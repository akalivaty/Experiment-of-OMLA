//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 0 0 1 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT64), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G137), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT11), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(G137), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT11), .ZN(new_n193));
  OAI211_X1 g007(.A(new_n188), .B(new_n193), .C1(new_n189), .C2(G137), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(new_n192), .A3(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G131), .ZN(new_n196));
  INV_X1    g010(.A(G131), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n191), .A2(new_n197), .A3(new_n192), .A4(new_n194), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  OR2_X1    g017(.A1(KEYINPUT0), .A2(G128), .ZN(new_n204));
  NAND2_X1  g018(.A1(KEYINPUT0), .A2(G128), .ZN(new_n205));
  AOI22_X1  g019(.A1(new_n201), .A2(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  AND3_X1   g020(.A1(new_n201), .A2(new_n203), .A3(new_n205), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n199), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G119), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G116), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT65), .B(G116), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n213), .B1(new_n214), .B2(G119), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n216));
  INV_X1    g030(.A(G113), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT2), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT2), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G113), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n215), .A2(new_n216), .A3(new_n221), .ZN(new_n222));
  AND2_X1   g036(.A1(KEYINPUT65), .A2(G116), .ZN(new_n223));
  NOR2_X1   g037(.A1(KEYINPUT65), .A2(G116), .ZN(new_n224));
  OAI21_X1  g038(.A(G119), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(new_n212), .A3(new_n221), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT66), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n212), .ZN(new_n228));
  INV_X1    g042(.A(new_n221), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n222), .A2(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G128), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(new_n201), .A3(new_n203), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n231), .A2(new_n200), .A3(G143), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n202), .B(G146), .C1(new_n231), .C2(KEYINPUT1), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n192), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n189), .A2(G137), .ZN(new_n238));
  OAI21_X1  g052(.A(G131), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n198), .A2(new_n236), .A3(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n210), .A2(new_n230), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n228), .A2(new_n229), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n216), .B1(new_n215), .B2(new_n221), .ZN(new_n243));
  AND4_X1   g057(.A1(new_n216), .A2(new_n225), .A3(new_n212), .A4(new_n221), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n208), .B1(new_n196), .B2(new_n198), .ZN(new_n246));
  INV_X1    g060(.A(new_n240), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n241), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT28), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n246), .A2(new_n247), .ZN(new_n251));
  AOI21_X1  g065(.A(KEYINPUT28), .B1(new_n251), .B2(new_n230), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  XOR2_X1   g067(.A(KEYINPUT26), .B(G101), .Z(new_n254));
  NOR2_X1   g068(.A1(G237), .A2(G953), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G210), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n254), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n257), .B(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n250), .A2(new_n253), .A3(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT29), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n187), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n264));
  OR2_X1    g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n264), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT30), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n267), .B1(new_n210), .B2(new_n240), .ZN(new_n268));
  NOR3_X1   g082(.A1(new_n246), .A2(new_n247), .A3(KEYINPUT30), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n245), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n241), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n262), .B(new_n261), .C1(new_n272), .C2(new_n260), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n265), .A2(new_n266), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G472), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(G472), .A2(G902), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n260), .B1(new_n250), .B2(new_n253), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n210), .A2(new_n267), .A3(new_n240), .ZN(new_n279));
  OAI21_X1  g093(.A(KEYINPUT30), .B1(new_n246), .B2(new_n247), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n230), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NOR3_X1   g095(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n282));
  NOR3_X1   g096(.A1(new_n281), .A2(new_n282), .A3(new_n259), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT31), .ZN(new_n284));
  OAI22_X1  g098(.A1(new_n278), .A2(KEYINPUT68), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT28), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n286), .B1(new_n241), .B2(new_n248), .ZN(new_n287));
  OAI211_X1 g101(.A(KEYINPUT68), .B(new_n259), .C1(new_n287), .C2(new_n252), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n270), .A2(new_n284), .A3(new_n241), .A4(new_n260), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NOR3_X1   g104(.A1(new_n285), .A2(KEYINPUT69), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT69), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n270), .A2(new_n241), .A3(new_n260), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n259), .B1(new_n287), .B2(new_n252), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT68), .ZN(new_n295));
  AOI22_X1  g109(.A1(KEYINPUT31), .A2(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n288), .A2(new_n289), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n292), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n277), .B1(new_n291), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT32), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT70), .ZN(new_n302));
  OAI211_X1 g116(.A(KEYINPUT32), .B(new_n277), .C1(new_n291), .C2(new_n298), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n299), .A2(KEYINPUT70), .A3(new_n300), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n276), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT25), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n231), .A2(G119), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n308), .B(KEYINPUT23), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n211), .A2(G128), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G110), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(KEYINPUT73), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n309), .A2(new_n312), .A3(new_n310), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT73), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n308), .A2(new_n310), .ZN(new_n317));
  XOR2_X1   g131(.A(KEYINPUT24), .B(G110), .Z(new_n318));
  OAI211_X1 g132(.A(new_n313), .B(new_n316), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT72), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT16), .ZN(new_n321));
  INV_X1    g135(.A(G140), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n322), .A3(G125), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(G125), .ZN(new_n324));
  INV_X1    g138(.A(G125), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G140), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n320), .B(new_n323), .C1(new_n327), .C2(new_n321), .ZN(new_n328));
  XNOR2_X1  g142(.A(G125), .B(G140), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(KEYINPUT72), .A3(KEYINPUT16), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n200), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n329), .A2(new_n200), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n319), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n317), .A2(new_n318), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n328), .A2(new_n200), .A3(new_n330), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  OAI221_X1 g151(.A(new_n335), .B1(new_n311), .B2(new_n312), .C1(new_n337), .C2(new_n331), .ZN(new_n338));
  INV_X1    g152(.A(G953), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(G221), .A3(G234), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n340), .B(KEYINPUT22), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n341), .B(G137), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n334), .A2(new_n338), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n342), .B1(new_n334), .B2(new_n338), .ZN(new_n344));
  NOR3_X1   g158(.A1(new_n343), .A2(new_n344), .A3(G902), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT74), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n307), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G217), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n348), .B1(G234), .B2(new_n187), .ZN(new_n349));
  INV_X1    g163(.A(new_n344), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n334), .A2(new_n338), .A3(new_n342), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n187), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(KEYINPUT74), .A3(KEYINPUT25), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n347), .A2(new_n349), .A3(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n349), .A2(G902), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT75), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n356), .B1(new_n350), .B2(new_n351), .ZN(new_n357));
  NOR3_X1   g171(.A1(new_n343), .A2(new_n344), .A3(KEYINPUT75), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n355), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n354), .A2(new_n359), .ZN(new_n360));
  XOR2_X1   g174(.A(KEYINPUT9), .B(G234), .Z(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(G221), .B1(new_n362), .B2(G902), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G469), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n365), .A2(new_n187), .ZN(new_n366));
  INV_X1    g180(.A(G107), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G104), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT3), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n369), .A2(KEYINPUT76), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT76), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n371), .A2(KEYINPUT3), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n368), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G101), .ZN(new_n374));
  OAI211_X1 g188(.A(G104), .B(new_n367), .C1(new_n369), .C2(KEYINPUT76), .ZN(new_n375));
  INV_X1    g189(.A(G104), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G107), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n373), .A2(new_n374), .A3(new_n375), .A4(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(KEYINPUT78), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT78), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(new_n376), .A3(G107), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n379), .A2(new_n381), .A3(new_n368), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G101), .ZN(new_n383));
  AND2_X1   g197(.A1(new_n378), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n384), .A2(new_n236), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n378), .A2(new_n383), .A3(new_n236), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n199), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT12), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n388), .B(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n391));
  INV_X1    g205(.A(new_n368), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n375), .B(new_n377), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT4), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(new_n394), .A3(G101), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT77), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n393), .A2(KEYINPUT77), .A3(new_n394), .A4(G101), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n394), .B1(new_n393), .B2(G101), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n397), .A2(new_n398), .B1(new_n378), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n209), .ZN(new_n401));
  INV_X1    g215(.A(new_n199), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT10), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n386), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n378), .A2(new_n383), .A3(KEYINPUT10), .A4(new_n236), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n401), .A2(new_n402), .A3(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n407), .A2(KEYINPUT79), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT79), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n404), .A2(new_n405), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n410), .B1(new_n209), .B2(new_n400), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n409), .B1(new_n411), .B2(new_n402), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n390), .B1(new_n408), .B2(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(G110), .B(G140), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n339), .A2(G227), .ZN(new_n415));
  XOR2_X1   g229(.A(new_n414), .B(new_n415), .Z(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n407), .A2(KEYINPUT79), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n411), .A2(new_n409), .A3(new_n402), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n411), .A2(new_n402), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  AOI22_X1  g236(.A1(new_n413), .A2(new_n417), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n366), .B1(new_n423), .B2(G469), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n420), .A2(new_n390), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n418), .A2(new_n419), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n416), .B1(new_n426), .B2(new_n422), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n365), .B(new_n187), .C1(new_n425), .C2(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n364), .B1(new_n424), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(G214), .B1(G237), .B2(G902), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n397), .A2(new_n398), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n399), .A2(new_n378), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(new_n245), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n222), .A2(new_n227), .ZN(new_n435));
  XNOR2_X1  g249(.A(KEYINPUT80), .B(KEYINPUT5), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n217), .B1(new_n436), .B2(new_n213), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n437), .B1(new_n228), .B2(new_n436), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n384), .A2(new_n435), .A3(KEYINPUT81), .A4(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT81), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n438), .B1(new_n243), .B2(new_n244), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n378), .A2(new_n383), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n434), .A2(new_n439), .A3(new_n443), .ZN(new_n444));
  XOR2_X1   g258(.A(G110), .B(G122), .Z(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n445), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n434), .A2(new_n443), .A3(new_n447), .A4(new_n439), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n446), .A2(KEYINPUT6), .A3(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT6), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n444), .A2(new_n450), .A3(new_n445), .ZN(new_n451));
  INV_X1    g265(.A(new_n236), .ZN(new_n452));
  AOI21_X1  g266(.A(KEYINPUT82), .B1(new_n452), .B2(new_n325), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(new_n325), .B2(new_n209), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n208), .A2(KEYINPUT82), .A3(G125), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n339), .A2(G224), .ZN(new_n457));
  XOR2_X1   g271(.A(new_n457), .B(KEYINPUT83), .Z(new_n458));
  XNOR2_X1  g272(.A(new_n456), .B(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n449), .A2(new_n451), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT85), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT5), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n461), .B1(new_n228), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n215), .A2(KEYINPUT85), .A3(KEYINPUT5), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n464), .A3(new_n437), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n435), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT86), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT86), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n465), .A2(new_n468), .A3(new_n435), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n467), .A2(new_n384), .A3(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(KEYINPUT84), .B(KEYINPUT8), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n445), .B(new_n471), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n470), .B(new_n472), .C1(new_n384), .C2(new_n441), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n457), .A2(KEYINPUT7), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n454), .A2(new_n474), .A3(new_n455), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n456), .A2(KEYINPUT7), .A3(new_n457), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n473), .A2(new_n475), .A3(new_n476), .A4(new_n448), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n460), .A2(new_n187), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(G210), .B1(G237), .B2(G902), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n460), .A2(new_n187), .A3(new_n477), .A4(new_n479), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n431), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n339), .A2(G952), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n484), .B1(G234), .B2(G237), .ZN(new_n485));
  XOR2_X1   g299(.A(KEYINPUT21), .B(G898), .Z(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(G234), .A2(G237), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n488), .A2(G902), .A3(G953), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n485), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT88), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n493), .B1(new_n231), .B2(G143), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n202), .A2(KEYINPUT88), .A3(G128), .ZN(new_n495));
  AOI22_X1  g309(.A1(new_n494), .A2(new_n495), .B1(KEYINPUT89), .B2(KEYINPUT13), .ZN(new_n496));
  NOR2_X1   g310(.A1(KEYINPUT89), .A2(KEYINPUT13), .ZN(new_n497));
  OR2_X1    g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT90), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n499), .B1(new_n202), .B2(G128), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n231), .A2(KEYINPUT90), .A3(G143), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n502), .B1(new_n496), .B2(new_n497), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n189), .B1(new_n498), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n494), .A2(new_n495), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n505), .A2(new_n189), .A3(new_n500), .A4(new_n501), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(G122), .B1(new_n223), .B2(new_n224), .ZN(new_n508));
  INV_X1    g322(.A(G122), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(G116), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n508), .A2(new_n367), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n367), .B1(new_n508), .B2(new_n510), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n504), .A2(new_n507), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(KEYINPUT91), .B1(new_n508), .B2(KEYINPUT14), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT91), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT14), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n214), .A2(new_n518), .A3(new_n519), .A4(G122), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n508), .A2(KEYINPUT14), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n517), .A2(new_n510), .A3(new_n520), .A4(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n512), .B1(new_n522), .B2(G107), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT92), .ZN(new_n524));
  INV_X1    g338(.A(new_n505), .ZN(new_n525));
  OAI21_X1  g339(.A(G134), .B1(new_n525), .B2(new_n502), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n506), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n523), .A2(new_n524), .A3(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n524), .B1(new_n523), .B2(new_n527), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n516), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NOR3_X1   g345(.A1(new_n362), .A2(new_n348), .A3(G953), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n523), .A2(new_n527), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT92), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n528), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(new_n516), .A3(new_n532), .ZN(new_n538));
  AOI21_X1  g352(.A(G902), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(G478), .ZN(new_n540));
  OR2_X1    g354(.A1(new_n540), .A2(KEYINPUT15), .ZN(new_n541));
  OR2_X1    g355(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n539), .A2(new_n541), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(G475), .ZN(new_n545));
  AOI21_X1  g359(.A(G143), .B1(new_n255), .B2(G214), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n255), .A2(G143), .A3(G214), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n197), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n548), .ZN(new_n550));
  NOR3_X1   g364(.A1(new_n550), .A2(new_n546), .A3(G131), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT17), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n549), .A2(KEYINPUT17), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n554), .A2(new_n336), .A3(new_n332), .A4(new_n555), .ZN(new_n556));
  OAI211_X1 g370(.A(KEYINPUT18), .B(G131), .C1(new_n550), .C2(new_n546), .ZN(new_n557));
  NAND2_X1  g371(.A1(KEYINPUT18), .A2(G131), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n547), .A2(new_n548), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n327), .A2(G146), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n333), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n557), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n556), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(G113), .B(G122), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(new_n376), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n556), .A2(new_n565), .A3(new_n562), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n545), .B1(new_n569), .B2(new_n187), .ZN(new_n570));
  INV_X1    g384(.A(new_n562), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n327), .A2(KEYINPUT19), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT19), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n329), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n575), .A2(G146), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n576), .A2(new_n331), .ZN(new_n577));
  INV_X1    g391(.A(new_n552), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n571), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(KEYINPUT87), .B1(new_n579), .B2(new_n565), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT87), .ZN(new_n581));
  NOR3_X1   g395(.A1(new_n552), .A2(new_n576), .A3(new_n331), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n581), .B(new_n566), .C1(new_n582), .C2(new_n571), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n580), .A2(new_n568), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(new_n545), .A3(new_n187), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT20), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT20), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n584), .A2(new_n587), .A3(new_n545), .A4(new_n187), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n570), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n544), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n429), .A2(new_n483), .A3(new_n492), .A4(new_n591), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n306), .A2(new_n360), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(new_n374), .ZN(G3));
  INV_X1    g408(.A(new_n277), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT69), .B1(new_n285), .B2(new_n290), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n296), .A2(new_n297), .A3(new_n292), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n187), .B1(new_n291), .B2(new_n298), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n598), .B1(new_n599), .B2(G472), .ZN(new_n600));
  INV_X1    g414(.A(new_n360), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n600), .A2(new_n601), .A3(new_n363), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n426), .A2(new_n422), .ZN(new_n603));
  AOI22_X1  g417(.A1(new_n603), .A2(new_n417), .B1(new_n420), .B2(new_n390), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n604), .A2(G469), .A3(G902), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n413), .A2(new_n417), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n420), .A2(new_n422), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n606), .A2(G469), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n366), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n602), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n532), .B1(new_n537), .B2(new_n516), .ZN(new_n613));
  AOI211_X1 g427(.A(new_n533), .B(new_n515), .C1(new_n536), .C2(new_n528), .ZN(new_n614));
  OAI21_X1  g428(.A(KEYINPUT33), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n534), .A2(new_n616), .A3(new_n538), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n615), .A2(new_n617), .A3(G478), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n539), .A2(new_n540), .ZN(new_n619));
  NAND2_X1  g433(.A1(G478), .A2(G902), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n621), .A2(new_n589), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n492), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT93), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n481), .A2(new_n482), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n625), .B1(new_n626), .B2(new_n430), .ZN(new_n627));
  AOI211_X1 g441(.A(KEYINPUT93), .B(new_n431), .C1(new_n481), .C2(new_n482), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n612), .A2(new_n624), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT94), .B(KEYINPUT34), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(G104), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n630), .B(new_n632), .ZN(G6));
  NAND2_X1  g447(.A1(new_n626), .A2(new_n430), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(KEYINPUT93), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n483), .A2(new_n625), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n544), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n588), .A2(KEYINPUT95), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n570), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n586), .A2(KEYINPUT95), .A3(new_n588), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n637), .A2(new_n638), .A3(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n643), .A2(new_n492), .A3(new_n612), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT35), .B(G107), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G9));
  INV_X1    g460(.A(KEYINPUT96), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n334), .A2(new_n338), .ZN(new_n648));
  INV_X1    g462(.A(new_n342), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(KEYINPUT36), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n648), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n355), .ZN(new_n652));
  AND3_X1   g466(.A1(new_n354), .A2(new_n647), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n647), .B1(new_n354), .B2(new_n652), .ZN(new_n654));
  OR2_X1    g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n656), .A2(KEYINPUT97), .A3(new_n600), .ZN(new_n657));
  INV_X1    g471(.A(new_n592), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT97), .ZN(new_n659));
  INV_X1    g473(.A(new_n600), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n659), .B1(new_n655), .B2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n657), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT37), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(new_n312), .ZN(G12));
  NAND2_X1  g478(.A1(new_n304), .A2(new_n305), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n655), .B1(new_n665), .B2(new_n275), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n363), .B1(new_n605), .B2(new_n610), .ZN(new_n667));
  INV_X1    g481(.A(new_n642), .ZN(new_n668));
  INV_X1    g482(.A(G900), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n485), .B1(new_n490), .B2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n668), .A2(new_n544), .A3(new_n671), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n637), .A2(new_n667), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n666), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G128), .ZN(G30));
  XOR2_X1   g489(.A(new_n670), .B(KEYINPUT39), .Z(new_n676));
  NAND2_X1  g490(.A1(new_n429), .A2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT98), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT40), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n430), .B1(new_n679), .B2(new_n680), .ZN(new_n682));
  XOR2_X1   g496(.A(new_n626), .B(KEYINPUT38), .Z(new_n683));
  NOR4_X1   g497(.A1(new_n681), .A2(new_n682), .A3(new_n656), .A4(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n272), .A2(new_n259), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n187), .B1(new_n249), .B2(new_n260), .ZN(new_n686));
  OAI21_X1  g500(.A(G472), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n688), .B1(new_n304), .B2(new_n305), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n689), .A2(new_n589), .A3(new_n638), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n684), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(KEYINPUT99), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT99), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n684), .A2(new_n693), .A3(new_n690), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT100), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(new_n202), .ZN(G45));
  INV_X1    g511(.A(new_n621), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n698), .A2(new_n590), .A3(new_n671), .ZN(new_n699));
  NOR4_X1   g513(.A1(new_n667), .A2(new_n627), .A3(new_n628), .A4(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n666), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(KEYINPUT101), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT101), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n666), .A2(new_n703), .A3(new_n700), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G146), .ZN(G48));
  NOR2_X1   g520(.A1(new_n306), .A2(new_n360), .ZN(new_n707));
  OAI21_X1  g521(.A(G469), .B1(new_n604), .B2(G902), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(new_n363), .A3(new_n428), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n709), .A2(new_n491), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n629), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n707), .A2(new_n622), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(KEYINPUT102), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT41), .B(G113), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G15));
  NAND3_X1  g529(.A1(new_n707), .A2(new_n643), .A3(new_n710), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G116), .ZN(G18));
  NAND3_X1  g531(.A1(new_n666), .A2(new_n591), .A3(new_n711), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G119), .ZN(G21));
  NOR2_X1   g533(.A1(new_n638), .A2(new_n589), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n635), .A2(new_n636), .A3(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT105), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n629), .A2(KEYINPUT105), .A3(new_n720), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(G902), .B1(new_n596), .B2(new_n597), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT103), .B(G472), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g542(.A(KEYINPUT104), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT104), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n599), .A2(new_n730), .A3(new_n727), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n294), .B1(new_n283), .B2(new_n284), .ZN(new_n732));
  INV_X1    g546(.A(new_n289), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n277), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n729), .A2(new_n731), .A3(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n360), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n725), .A2(new_n710), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  NOR4_X1   g552(.A1(new_n627), .A2(new_n628), .A3(new_n699), .A4(new_n709), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n655), .A2(new_n735), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G125), .ZN(G27));
  INV_X1    g556(.A(KEYINPUT42), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n481), .A2(new_n430), .A3(new_n482), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n667), .A2(new_n699), .A3(new_n744), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n598), .A2(KEYINPUT32), .B1(new_n274), .B2(G472), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n360), .B1(new_n746), .B2(new_n301), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n743), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n744), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n429), .A2(new_n749), .A3(new_n622), .A4(new_n671), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n750), .A2(KEYINPUT42), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n748), .B1(new_n707), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G131), .ZN(G33));
  INV_X1    g567(.A(new_n672), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n707), .A2(new_n429), .A3(new_n754), .A4(new_n749), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G134), .ZN(G36));
  NAND2_X1  g570(.A1(new_n423), .A2(KEYINPUT45), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n758));
  AOI211_X1 g572(.A(new_n417), .B(new_n421), .C1(new_n419), .C2(new_n418), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n416), .B1(new_n426), .B2(new_n390), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n757), .A2(G469), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(KEYINPUT106), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT106), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n757), .A2(new_n764), .A3(new_n761), .A4(G469), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n366), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n428), .B1(new_n766), .B2(KEYINPUT46), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT46), .ZN(new_n768));
  AOI211_X1 g582(.A(new_n768), .B(new_n366), .C1(new_n763), .C2(new_n765), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n363), .B(new_n676), .C1(new_n767), .C2(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n590), .A2(new_n621), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT107), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(KEYINPUT43), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n771), .B1(new_n773), .B2(KEYINPUT43), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n775), .B1(new_n776), .B2(new_n774), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(new_n660), .A3(new_n656), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n770), .B1(KEYINPUT44), .B2(new_n779), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n780), .B(new_n749), .C1(KEYINPUT44), .C2(new_n779), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G137), .ZN(G39));
  OAI21_X1  g596(.A(new_n363), .B1(new_n767), .B2(new_n769), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT108), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI211_X1 g599(.A(KEYINPUT108), .B(new_n363), .C1(new_n767), .C2(new_n769), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  XOR2_X1   g604(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n785), .A2(new_n792), .A3(new_n786), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n665), .A2(new_n275), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n794), .A2(new_n699), .A3(new_n744), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n790), .A2(new_n360), .A3(new_n793), .A4(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G140), .ZN(G42));
  AND2_X1   g611(.A1(new_n708), .A2(new_n428), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n771), .B1(new_n799), .B2(KEYINPUT49), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n800), .B1(KEYINPUT49), .B2(new_n799), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n360), .A2(new_n431), .A3(new_n364), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n801), .A2(new_n689), .A3(new_n683), .A4(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT116), .ZN(new_n804));
  INV_X1    g618(.A(new_n709), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n749), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT115), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n689), .A2(new_n601), .A3(new_n485), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n809), .A2(new_n589), .A3(new_n621), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n736), .A2(new_n777), .A3(new_n485), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n790), .A2(new_n793), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n798), .A2(new_n364), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n811), .B1(new_n815), .B2(new_n749), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n683), .A2(new_n431), .A3(new_n805), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(KEYINPUT113), .ZN(new_n818));
  OR2_X1    g632(.A1(KEYINPUT114), .A2(KEYINPUT50), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n818), .A2(new_n819), .A3(new_n812), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(KEYINPUT114), .A2(KEYINPUT50), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n819), .B(new_n822), .C1(new_n818), .C2(new_n812), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n777), .A2(new_n485), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n807), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n740), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n816), .A2(new_n821), .A3(new_n823), .A4(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT51), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n804), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n793), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n788), .B1(new_n785), .B2(new_n786), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n814), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n812), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n832), .A2(new_n749), .A3(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n834), .A2(new_n823), .A3(new_n826), .A4(new_n810), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n836), .A2(KEYINPUT116), .A3(KEYINPUT51), .A4(new_n821), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n829), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n828), .B1(new_n835), .B2(new_n820), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n354), .A2(new_n652), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n689), .A2(new_n840), .A3(new_n670), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n841), .A2(new_n725), .A3(new_n429), .ZN(new_n842));
  AOI22_X1  g656(.A1(new_n666), .A2(new_n673), .B1(new_n740), .B2(new_n739), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n666), .A2(new_n703), .A3(new_n700), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n703), .B1(new_n666), .B2(new_n700), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n842), .B(new_n843), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n705), .A2(KEYINPUT52), .A3(new_n843), .A4(new_n842), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NOR4_X1   g664(.A1(new_n602), .A2(new_n634), .A3(new_n611), .A4(new_n623), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT110), .B1(new_n593), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n794), .A2(new_n658), .A3(new_n601), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n612), .A2(new_n483), .A3(new_n624), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT110), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n544), .A2(new_n589), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(KEYINPUT111), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n612), .A2(new_n483), .A3(new_n492), .A4(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n852), .A2(new_n856), .A3(new_n662), .A4(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n750), .A2(new_n735), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n542), .A2(new_n543), .A3(new_n671), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n642), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n749), .A2(new_n863), .A3(KEYINPUT112), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(new_n429), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n306), .A2(new_n865), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n744), .A2(new_n642), .A3(new_n862), .ZN(new_n867));
  OR2_X1    g681(.A1(new_n867), .A2(KEYINPUT112), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n861), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n752), .B(new_n755), .C1(new_n869), .C2(new_n655), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n737), .A2(new_n712), .A3(new_n716), .A4(new_n718), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n860), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n850), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT53), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT54), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n850), .A2(new_n872), .A3(KEYINPUT53), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n850), .A2(new_n872), .A3(KEYINPUT53), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT53), .B1(new_n850), .B2(new_n872), .ZN(new_n880));
  OAI21_X1  g694(.A(KEYINPUT54), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n812), .A2(new_n637), .A3(new_n709), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n882), .B1(new_n622), .B2(new_n809), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n839), .A2(new_n878), .A3(new_n881), .A4(new_n883), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n484), .B(KEYINPUT117), .Z(new_n885));
  NAND2_X1  g699(.A1(new_n825), .A2(new_n747), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n886), .B(KEYINPUT48), .Z(new_n887));
  NOR4_X1   g701(.A1(new_n838), .A2(new_n884), .A3(new_n885), .A4(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(G952), .A2(G953), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(KEYINPUT118), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n803), .B1(new_n888), .B2(new_n890), .ZN(G75));
  AOI21_X1  g705(.A(new_n187), .B1(new_n875), .B2(new_n877), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(G210), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT56), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n449), .A2(new_n451), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(new_n459), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT55), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n893), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n897), .B1(new_n893), .B2(new_n894), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n339), .A2(G952), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(G51));
  XNOR2_X1  g715(.A(new_n366), .B(KEYINPUT57), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT119), .B1(new_n881), .B2(new_n878), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT119), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n875), .A2(new_n877), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n904), .B1(new_n905), .B2(KEYINPUT54), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n902), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(KEYINPUT120), .ZN(new_n908));
  INV_X1    g722(.A(new_n604), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT120), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n910), .B(new_n902), .C1(new_n903), .C2(new_n906), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n908), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n892), .A2(new_n765), .A3(new_n763), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n900), .B1(new_n912), .B2(new_n913), .ZN(G54));
  NAND3_X1  g728(.A1(new_n892), .A2(KEYINPUT58), .A3(G475), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(new_n584), .Z(new_n916));
  NOR2_X1   g730(.A1(new_n916), .A2(new_n900), .ZN(G60));
  NAND2_X1  g731(.A1(new_n615), .A2(new_n617), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n620), .B(KEYINPUT59), .Z(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n918), .B(new_n920), .C1(new_n903), .C2(new_n906), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n919), .B1(new_n881), .B2(new_n878), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n922), .A2(new_n918), .ZN(new_n923));
  INV_X1    g737(.A(new_n900), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n921), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT121), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n921), .A2(new_n923), .A3(KEYINPUT121), .A4(new_n924), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(G63));
  NAND2_X1  g743(.A1(G217), .A2(G902), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT60), .Z(new_n931));
  NAND3_X1  g745(.A1(new_n905), .A2(new_n651), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n924), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n357), .A2(new_n358), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT122), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n935), .B1(new_n905), .B2(new_n931), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n937));
  OAI22_X1  g751(.A1(new_n933), .A2(new_n936), .B1(KEYINPUT123), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(KEYINPUT123), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT124), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n938), .B(new_n940), .ZN(G66));
  INV_X1    g755(.A(G224), .ZN(new_n942));
  OAI21_X1  g756(.A(G953), .B1(new_n487), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n860), .A2(new_n871), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n943), .B1(new_n944), .B2(G953), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n895), .B1(G898), .B2(new_n339), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(G69));
  NOR2_X1   g761(.A1(new_n268), .A2(new_n269), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT125), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(new_n575), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n705), .A2(new_n843), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n692), .A2(new_n694), .A3(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT62), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(new_n955));
  OR2_X1    g769(.A1(new_n858), .A2(new_n622), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n707), .A2(new_n679), .A3(new_n956), .A4(new_n749), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n796), .A2(new_n781), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n950), .B1(new_n959), .B2(new_n339), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n339), .B1(G227), .B2(G900), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n950), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n752), .A2(new_n755), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(KEYINPUT126), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n796), .A2(new_n781), .A3(new_n952), .A4(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n725), .A2(new_n747), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n968), .A2(new_n770), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n965), .A2(KEYINPUT126), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n967), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n964), .B1(new_n971), .B2(new_n339), .ZN(new_n972));
  NAND2_X1  g786(.A1(G900), .A2(G953), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n961), .A2(new_n963), .A3(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n974), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n962), .B1(new_n960), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n975), .A2(new_n977), .ZN(G72));
  NAND2_X1  g792(.A1(G472), .A2(G902), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT63), .Z(new_n980));
  INV_X1    g794(.A(new_n944), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n980), .B1(new_n959), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n900), .B1(new_n982), .B2(new_n685), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n272), .A2(new_n260), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n905), .B(new_n980), .C1(new_n984), .C2(new_n283), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n971), .A2(new_n944), .ZN(new_n986));
  INV_X1    g800(.A(new_n980), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n259), .B(new_n272), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n983), .A2(new_n985), .A3(new_n988), .ZN(G57));
endmodule


