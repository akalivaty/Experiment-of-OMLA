//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 1 0 1 1 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n814, new_n815, new_n817, new_n818, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924;
  INV_X1    g000(.A(KEYINPUT95), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G43gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G99gat), .ZN(new_n204));
  XOR2_X1   g003(.A(KEYINPUT72), .B(G71gat), .Z(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G227gat), .A2(G233gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n207), .B(KEYINPUT64), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT70), .B(KEYINPUT1), .ZN(new_n209));
  XNOR2_X1  g008(.A(KEYINPUT68), .B(G120gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G113gat), .ZN(new_n211));
  INV_X1    g010(.A(G113gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G120gat), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n209), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G127gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G134gat), .ZN(new_n216));
  INV_X1    g015(.A(G134gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G127gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT69), .ZN(new_n219));
  AND3_X1   g018(.A1(new_n216), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n219), .B1(new_n216), .B2(new_n218), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT1), .ZN(new_n223));
  INV_X1    g022(.A(G120gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G113gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n213), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G127gat), .B(G134gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n223), .A2(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n215), .A2(KEYINPUT67), .A3(G134gat), .ZN(new_n230));
  AOI22_X1  g029(.A1(new_n214), .A2(new_n222), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OR2_X1    g030(.A1(G183gat), .A2(G190gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(G183gat), .A2(G190gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n232), .A2(KEYINPUT24), .A3(new_n233), .ZN(new_n234));
  OR2_X1    g033(.A1(new_n233), .A2(KEYINPUT24), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(G169gat), .A2(G176gat), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G169gat), .A2(G176gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT23), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT25), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n243), .B1(new_n238), .B2(KEYINPUT23), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n237), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(G169gat), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT65), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n248), .A2(G176gat), .ZN(new_n249));
  INV_X1    g048(.A(G176gat), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n250), .A2(KEYINPUT65), .ZN(new_n251));
  OAI211_X1 g050(.A(KEYINPUT23), .B(new_n247), .C1(new_n249), .C2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT66), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n252), .A2(new_n253), .A3(new_n242), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n253), .B1(new_n252), .B2(new_n242), .ZN(new_n255));
  NOR3_X1   g054(.A1(new_n254), .A2(new_n255), .A3(new_n236), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n246), .B1(new_n256), .B2(KEYINPUT25), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT27), .B(G183gat), .ZN(new_n258));
  INV_X1    g057(.A(G190gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OR2_X1    g059(.A1(new_n260), .A2(KEYINPUT28), .ZN(new_n261));
  OR2_X1    g060(.A1(new_n239), .A2(KEYINPUT26), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n239), .A2(KEYINPUT26), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n262), .A2(new_n240), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n260), .A2(KEYINPUT28), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n261), .A2(new_n233), .A3(new_n264), .A4(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n231), .B1(new_n257), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT23), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n250), .A2(KEYINPUT65), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n248), .A2(G176gat), .ZN(new_n270));
  AOI211_X1 g069(.A(new_n268), .B(G169gat), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n242), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT66), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n252), .A2(new_n253), .A3(new_n242), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n273), .A2(new_n237), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n245), .B1(new_n275), .B2(new_n243), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n226), .A2(new_n223), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n227), .A2(new_n228), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n277), .A2(new_n278), .A3(new_n230), .ZN(new_n279));
  INV_X1    g078(.A(new_n221), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n227), .A2(new_n219), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n209), .ZN(new_n283));
  OR2_X1    g082(.A1(KEYINPUT68), .A2(G120gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(KEYINPUT68), .A2(G120gat), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n212), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n213), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n283), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n279), .B1(new_n282), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n266), .ZN(new_n290));
  NOR3_X1   g089(.A1(new_n276), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n208), .B1(new_n267), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n206), .B1(new_n292), .B2(KEYINPUT32), .ZN(new_n293));
  INV_X1    g092(.A(new_n208), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n257), .A2(new_n231), .A3(new_n266), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n289), .B1(new_n276), .B2(new_n290), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(KEYINPUT71), .B1(new_n297), .B2(KEYINPUT33), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT71), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT33), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n292), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n293), .A2(new_n298), .A3(new_n301), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n292), .B(KEYINPUT32), .C1(new_n300), .C2(new_n206), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT34), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n295), .A2(new_n296), .A3(new_n305), .A4(new_n294), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT73), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n306), .B(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n295), .A2(new_n296), .A3(new_n294), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT34), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n304), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n302), .A2(new_n303), .A3(new_n310), .A4(new_n308), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n312), .A2(KEYINPUT36), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT74), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT74), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n312), .A2(new_n316), .A3(KEYINPUT36), .A4(new_n313), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT76), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n312), .A2(new_n319), .A3(new_n313), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n304), .A2(KEYINPUT76), .A3(new_n311), .ZN(new_n321));
  XOR2_X1   g120(.A(KEYINPUT75), .B(KEYINPUT36), .Z(new_n322));
  NAND3_X1  g121(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(KEYINPUT80), .A2(KEYINPUT30), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT77), .B(G211gat), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT22), .B1(new_n326), .B2(G218gat), .ZN(new_n327));
  XOR2_X1   g126(.A(G197gat), .B(G204gat), .Z(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  XOR2_X1   g128(.A(G211gat), .B(G218gat), .Z(new_n330));
  XNOR2_X1  g129(.A(new_n329), .B(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(G226gat), .A2(G233gat), .ZN(new_n333));
  XOR2_X1   g132(.A(new_n333), .B(KEYINPUT78), .Z(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT29), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n337), .B1(new_n257), .B2(new_n266), .ZN(new_n338));
  NOR3_X1   g137(.A1(new_n276), .A2(new_n290), .A3(new_n335), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n332), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n336), .B(new_n335), .C1(new_n276), .C2(new_n290), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n257), .A2(new_n266), .A3(new_n334), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n341), .A2(new_n342), .A3(new_n331), .ZN(new_n343));
  XNOR2_X1  g142(.A(G8gat), .B(G36gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(G64gat), .B(G92gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n344), .B(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n340), .A2(new_n343), .A3(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT80), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT30), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n325), .B1(new_n348), .B2(new_n352), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n340), .A2(new_n343), .A3(new_n347), .A4(new_n351), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n347), .B1(new_n340), .B2(new_n343), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT79), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI211_X1 g156(.A(KEYINPUT79), .B(new_n347), .C1(new_n340), .C2(new_n343), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n353), .B(new_n354), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(G141gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n361), .A2(G148gat), .ZN(new_n362));
  INV_X1    g161(.A(G148gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n363), .A2(G141gat), .ZN(new_n364));
  OAI21_X1  g163(.A(KEYINPUT81), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT2), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n363), .A2(G141gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n361), .A2(G148gat), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT81), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n365), .A2(new_n366), .A3(new_n370), .ZN(new_n371));
  AND2_X1   g170(.A1(G155gat), .A2(G162gat), .ZN(new_n372));
  NOR2_X1   g171(.A1(G155gat), .A2(G162gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(G162gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT83), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT83), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(G162gat), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n377), .A2(new_n379), .A3(G155gat), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n374), .B1(new_n380), .B2(KEYINPUT2), .ZN(new_n381));
  AND2_X1   g180(.A1(KEYINPUT82), .A2(G141gat), .ZN(new_n382));
  NOR2_X1   g181(.A1(KEYINPUT82), .A2(G141gat), .ZN(new_n383));
  OAI21_X1  g182(.A(G148gat), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n367), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n375), .A2(new_n386), .ZN(new_n387));
  NOR3_X1   g186(.A1(new_n387), .A2(new_n289), .A3(KEYINPUT4), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT4), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n371), .A2(new_n374), .B1(new_n381), .B2(new_n385), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n389), .B1(new_n231), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(G225gat), .A2(G233gat), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n394), .A2(new_n389), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT84), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT3), .ZN(new_n398));
  AND3_X1   g197(.A1(new_n375), .A2(new_n398), .A3(new_n386), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n398), .B1(new_n375), .B2(new_n386), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n397), .B1(new_n401), .B2(new_n289), .ZN(new_n402));
  INV_X1    g201(.A(new_n374), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n369), .B1(new_n367), .B2(new_n368), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n403), .B1(new_n406), .B2(new_n366), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n380), .A2(KEYINPUT2), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n385), .A2(new_n408), .A3(new_n403), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT3), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n390), .A2(new_n398), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n410), .A2(new_n411), .A3(new_n397), .A4(new_n289), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n393), .B(new_n396), .C1(new_n402), .C2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n394), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n387), .A2(new_n289), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n231), .A2(new_n390), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT5), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n410), .A2(new_n289), .A3(new_n411), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT84), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n392), .B1(new_n422), .B2(new_n412), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n415), .A2(KEYINPUT5), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n414), .A2(new_n420), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  XOR2_X1   g224(.A(G57gat), .B(G85gat), .Z(new_n426));
  XNOR2_X1  g225(.A(G1gat), .B(G29gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  XOR2_X1   g227(.A(KEYINPUT85), .B(KEYINPUT0), .Z(new_n429));
  XNOR2_X1  g228(.A(new_n429), .B(KEYINPUT86), .ZN(new_n430));
  XOR2_X1   g229(.A(new_n428), .B(new_n430), .Z(new_n431));
  AOI21_X1  g230(.A(KEYINPUT6), .B1(new_n425), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n431), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n419), .B1(new_n423), .B2(new_n396), .ZN(new_n434));
  INV_X1    g233(.A(new_n424), .ZN(new_n435));
  AOI211_X1 g234(.A(new_n435), .B(new_n392), .C1(new_n422), .C2(new_n412), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n433), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  OAI211_X1 g236(.A(KEYINPUT6), .B(new_n433), .C1(new_n434), .C2(new_n436), .ZN(new_n438));
  AOI22_X1  g237(.A1(new_n432), .A2(new_n437), .B1(new_n438), .B2(KEYINPUT87), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT6), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n423), .A2(new_n424), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n416), .A2(new_n389), .ZN(new_n442));
  INV_X1    g241(.A(new_n391), .ZN(new_n443));
  AOI221_X4 g242(.A(new_n395), .B1(new_n442), .B2(new_n443), .C1(new_n422), .C2(new_n412), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n431), .B(new_n441), .C1(new_n444), .C2(new_n419), .ZN(new_n445));
  AND4_X1   g244(.A1(KEYINPUT87), .A2(new_n437), .A3(new_n440), .A4(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n360), .B1(new_n439), .B2(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(G78gat), .B(G106gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n448), .B(KEYINPUT31), .ZN(new_n449));
  XNOR2_X1  g248(.A(KEYINPUT88), .B(G50gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n449), .B(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n451), .B(KEYINPUT89), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n398), .B1(new_n331), .B2(KEYINPUT29), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n453), .A2(new_n387), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n332), .B1(new_n336), .B2(new_n411), .ZN(new_n455));
  NAND2_X1  g254(.A1(G228gat), .A2(G233gat), .ZN(new_n456));
  XOR2_X1   g255(.A(new_n456), .B(G22gat), .Z(new_n457));
  OR3_X1    g256(.A1(new_n454), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n457), .B1(new_n454), .B2(new_n455), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n452), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n451), .A2(KEYINPUT89), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n458), .A2(new_n459), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n447), .A2(new_n464), .ZN(new_n465));
  XOR2_X1   g264(.A(new_n431), .B(KEYINPUT90), .Z(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n467), .B1(new_n434), .B2(new_n436), .ZN(new_n468));
  OR3_X1    g267(.A1(new_n416), .A2(new_n417), .A3(new_n415), .ZN(new_n469));
  OAI211_X1 g268(.A(KEYINPUT39), .B(new_n469), .C1(new_n423), .C2(new_n394), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n393), .B1(new_n402), .B2(new_n413), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT39), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n471), .A2(new_n472), .A3(new_n415), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n470), .A2(new_n473), .A3(new_n466), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT40), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n468), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n353), .A2(new_n354), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n355), .B(new_n356), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n474), .A2(KEYINPUT91), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT91), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n470), .A2(new_n473), .A3(new_n481), .A4(new_n466), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n480), .A2(new_n475), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT92), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n480), .A2(KEYINPUT92), .A3(new_n475), .A4(new_n482), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n479), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n438), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n488), .B1(new_n432), .B2(new_n468), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n340), .A2(new_n343), .ZN(new_n490));
  OR2_X1    g289(.A1(new_n490), .A2(KEYINPUT37), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(KEYINPUT37), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n346), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT38), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n341), .A2(new_n342), .A3(KEYINPUT93), .A4(new_n331), .ZN(new_n495));
  OAI211_X1 g294(.A(KEYINPUT37), .B(new_n495), .C1(new_n490), .C2(KEYINPUT93), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT38), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n496), .A2(new_n491), .A3(new_n497), .A4(new_n346), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n489), .A2(new_n348), .A3(new_n494), .A4(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n487), .A2(new_n463), .A3(new_n499), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n324), .A2(new_n465), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n320), .A2(new_n321), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT35), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n477), .A2(new_n503), .A3(new_n478), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n504), .A2(new_n489), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n502), .A2(new_n505), .A3(new_n463), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n312), .A2(new_n463), .A3(new_n313), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT35), .B1(new_n447), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT94), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AND3_X1   g309(.A1(new_n312), .A2(new_n463), .A3(new_n313), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n437), .A2(new_n445), .A3(new_n440), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n438), .A2(KEYINPUT87), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n432), .A2(KEYINPUT87), .A3(new_n437), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n359), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n517), .A2(KEYINPUT94), .A3(KEYINPUT35), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n506), .B1(new_n510), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n202), .B1(new_n501), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n502), .A2(new_n505), .A3(new_n463), .ZN(new_n521));
  AOI21_X1  g320(.A(KEYINPUT94), .B1(new_n517), .B2(KEYINPUT35), .ZN(new_n522));
  AOI211_X1 g321(.A(new_n509), .B(new_n503), .C1(new_n511), .C2(new_n516), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n324), .A2(new_n465), .A3(new_n500), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(KEYINPUT95), .A3(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G113gat), .B(G141gat), .ZN(new_n527));
  INV_X1    g326(.A(G197gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(KEYINPUT11), .B(G169gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(KEYINPUT12), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NOR2_X1   g332(.A1(G29gat), .A2(G36gat), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT14), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G43gat), .B(G50gat), .ZN(new_n537));
  INV_X1    g336(.A(G29gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(KEYINPUT96), .B(G36gat), .ZN(new_n539));
  OAI221_X1 g338(.A(new_n536), .B1(KEYINPUT15), .B2(new_n537), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n537), .A2(KEYINPUT15), .ZN(new_n541));
  XOR2_X1   g340(.A(new_n540), .B(new_n541), .Z(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(KEYINPUT17), .ZN(new_n543));
  INV_X1    g342(.A(G8gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(G15gat), .B(G22gat), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n545), .A2(G1gat), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n544), .B1(new_n546), .B2(KEYINPUT97), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT16), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n545), .B1(new_n548), .B2(G1gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n547), .B(new_n550), .Z(new_n551));
  NAND2_X1  g350(.A1(new_n543), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(G229gat), .A2(G233gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n547), .B(new_n550), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n542), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n552), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT18), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n552), .A2(KEYINPUT18), .A3(new_n553), .A4(new_n555), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n542), .B(new_n554), .ZN(new_n561));
  XOR2_X1   g360(.A(KEYINPUT98), .B(KEYINPUT13), .Z(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(new_n553), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT99), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n533), .B1(new_n560), .B2(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n564), .B(KEYINPUT99), .Z(new_n567));
  NAND4_X1  g366(.A1(new_n567), .A2(new_n532), .A3(new_n559), .A4(new_n558), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G85gat), .A2(G92gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT7), .ZN(new_n571));
  NAND2_X1  g370(.A1(G99gat), .A2(G106gat), .ZN(new_n572));
  INV_X1    g371(.A(G85gat), .ZN(new_n573));
  INV_X1    g372(.A(G92gat), .ZN(new_n574));
  AOI22_X1  g373(.A1(KEYINPUT8), .A2(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AND2_X1   g374(.A1(new_n575), .A2(KEYINPUT104), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n575), .A2(KEYINPUT104), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n571), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(G99gat), .B(G106gat), .Z(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(G71gat), .A2(G78gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT9), .ZN(new_n583));
  INV_X1    g382(.A(G71gat), .ZN(new_n584));
  INV_X1    g383(.A(G78gat), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(KEYINPUT101), .B(G57gat), .ZN(new_n587));
  INV_X1    g386(.A(G64gat), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n588), .A2(G57gat), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n586), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT102), .ZN(new_n592));
  XOR2_X1   g391(.A(new_n582), .B(KEYINPUT100), .Z(new_n593));
  NOR2_X1   g392(.A1(new_n588), .A2(G57gat), .ZN(new_n594));
  OAI21_X1  g393(.A(KEYINPUT9), .B1(new_n590), .B2(new_n594), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n593), .B(new_n595), .C1(new_n584), .C2(new_n585), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n581), .A2(KEYINPUT10), .A3(new_n592), .A4(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n592), .A2(new_n596), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n581), .B(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n597), .B1(new_n600), .B2(KEYINPUT10), .ZN(new_n601));
  NAND2_X1  g400(.A1(G230gat), .A2(G233gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n603), .B1(new_n599), .B2(new_n602), .ZN(new_n604));
  XNOR2_X1  g403(.A(G120gat), .B(G148gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(G176gat), .B(G204gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  OR2_X1    g406(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n604), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n520), .A2(new_n526), .A3(new_n569), .A4(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT21), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n551), .B1(new_n598), .B2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(G183gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n613), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n615), .B(new_n616), .Z(new_n617));
  AND2_X1   g416(.A1(G231gat), .A2(G233gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G127gat), .B(G155gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(G211gat), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n619), .A2(new_n622), .ZN(new_n627));
  NOR3_X1   g426(.A1(new_n624), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n617), .B(new_n618), .Z(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n621), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n625), .B1(new_n630), .B2(new_n623), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT103), .B(G134gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(new_n376), .ZN(new_n634));
  AOI21_X1  g433(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n543), .A2(new_n580), .ZN(new_n637));
  NAND3_X1  g436(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n542), .A2(new_n581), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G190gat), .B(G218gat), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n636), .B1(new_n642), .B2(KEYINPUT105), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n640), .B(new_n641), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n632), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n612), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n439), .A2(new_n446), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n648), .B(KEYINPUT106), .Z(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(G1gat), .ZN(G1324gat));
  NOR3_X1   g451(.A1(new_n612), .A2(new_n646), .A3(new_n360), .ZN(new_n653));
  NAND2_X1  g452(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n548), .A2(new_n544), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT42), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n658), .B(new_n659), .C1(new_n544), .C2(new_n653), .ZN(G1325gat));
  AOI21_X1  g459(.A(G15gat), .B1(new_n647), .B2(new_n502), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n324), .A2(KEYINPUT107), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT107), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n318), .A2(new_n663), .A3(new_n323), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  AND2_X1   g465(.A1(new_n666), .A2(G15gat), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n661), .B1(new_n647), .B2(new_n667), .ZN(G1326gat));
  NAND2_X1  g467(.A1(new_n647), .A2(new_n464), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT43), .B(G22gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1327gat));
  NOR3_X1   g470(.A1(new_n612), .A2(new_n645), .A3(new_n632), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n672), .A2(new_n538), .A3(new_n650), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT45), .ZN(new_n674));
  INV_X1    g473(.A(new_n645), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n520), .A2(new_n675), .A3(new_n526), .ZN(new_n676));
  AND3_X1   g475(.A1(new_n676), .A2(KEYINPUT109), .A3(KEYINPUT44), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n500), .A2(new_n465), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n679), .B1(new_n662), .B2(new_n664), .ZN(new_n680));
  OAI211_X1 g479(.A(new_n678), .B(new_n675), .C1(new_n680), .C2(new_n519), .ZN(new_n681));
  AOI22_X1  g480(.A1(new_n676), .A2(KEYINPUT44), .B1(new_n681), .B2(KEYINPUT109), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n626), .B1(new_n624), .B2(new_n627), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n630), .A2(new_n623), .A3(new_n625), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n610), .B(KEYINPUT108), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n686), .A2(new_n569), .A3(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  AND3_X1   g488(.A1(new_n683), .A2(new_n650), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n674), .B1(new_n690), .B2(new_n538), .ZN(G1328gat));
  NAND3_X1  g490(.A1(new_n672), .A2(new_n539), .A3(new_n359), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(KEYINPUT46), .ZN(new_n693));
  OR2_X1    g492(.A1(new_n692), .A2(KEYINPUT46), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n683), .A2(new_n359), .A3(new_n689), .ZN(new_n695));
  OAI211_X1 g494(.A(new_n693), .B(new_n694), .C1(new_n695), .C2(new_n539), .ZN(G1329gat));
  NAND4_X1  g495(.A1(new_n683), .A2(G43gat), .A3(new_n666), .A4(new_n689), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n672), .A2(new_n502), .ZN(new_n698));
  INV_X1    g497(.A(G43gat), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g500(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1330gat));
  INV_X1    g502(.A(G50gat), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n672), .A2(new_n704), .A3(new_n464), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n464), .B(new_n689), .C1(new_n677), .C2(new_n682), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n705), .B1(G50gat), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(KEYINPUT48), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT112), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n706), .A2(new_n709), .A3(G50gat), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n709), .B1(new_n706), .B2(G50gat), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n710), .A2(new_n711), .A3(new_n705), .ZN(new_n712));
  XOR2_X1   g511(.A(KEYINPUT111), .B(KEYINPUT48), .Z(new_n713));
  OAI21_X1  g512(.A(new_n708), .B1(new_n712), .B2(new_n713), .ZN(G1331gat));
  OR2_X1    g513(.A1(new_n680), .A2(new_n519), .ZN(new_n715));
  INV_X1    g514(.A(new_n687), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n686), .A2(new_n675), .A3(new_n569), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT113), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT113), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n715), .A2(new_n720), .A3(new_n717), .A4(new_n716), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n719), .A2(new_n650), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(new_n587), .ZN(G1332gat));
  AOI21_X1  g522(.A(KEYINPUT114), .B1(new_n719), .B2(new_n721), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n719), .A2(KEYINPUT114), .A3(new_n721), .ZN(new_n726));
  AND3_X1   g525(.A1(new_n725), .A2(new_n359), .A3(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n728));
  AND2_X1   g527(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n727), .B2(new_n728), .ZN(G1333gat));
  NAND4_X1  g530(.A1(new_n725), .A2(G71gat), .A3(new_n666), .A4(new_n726), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n719), .A2(new_n502), .A3(new_n721), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n584), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT50), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT50), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n732), .A2(new_n737), .A3(new_n734), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(G1334gat));
  NAND3_X1  g538(.A1(new_n725), .A2(new_n464), .A3(new_n726), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g540(.A1(new_n632), .A2(new_n569), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n715), .A2(new_n675), .A3(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT51), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT115), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n649), .A2(G85gat), .A3(new_n611), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT116), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n610), .B(new_n742), .C1(new_n677), .C2(new_n682), .ZN(new_n750));
  OAI21_X1  g549(.A(G85gat), .B1(new_n750), .B2(new_n649), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(G1336gat));
  OAI21_X1  g551(.A(G92gat), .B1(new_n750), .B2(new_n360), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n687), .A2(G92gat), .A3(new_n360), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT52), .B1(new_n745), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT117), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n715), .A2(new_n757), .A3(new_n675), .A4(new_n742), .ZN(new_n758));
  AOI21_X1  g557(.A(KEYINPUT51), .B1(new_n758), .B2(KEYINPUT118), .ZN(new_n759));
  AOI21_X1  g558(.A(KEYINPUT117), .B1(KEYINPUT118), .B2(KEYINPUT51), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n759), .B1(new_n743), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n754), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n763), .A2(new_n753), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n756), .B1(new_n764), .B2(new_n765), .ZN(G1337gat));
  INV_X1    g565(.A(new_n502), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n611), .A2(new_n767), .A3(G99gat), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n746), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(G99gat), .B1(new_n750), .B2(new_n665), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(G1338gat));
  NOR3_X1   g570(.A1(new_n687), .A2(G106gat), .A3(new_n463), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n762), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(G106gat), .B1(new_n750), .B2(new_n463), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT53), .ZN(new_n776));
  XNOR2_X1  g575(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n777), .B1(new_n745), .B2(new_n772), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT120), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n774), .A2(new_n778), .A3(KEYINPUT120), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n776), .A2(new_n781), .A3(new_n782), .ZN(G1339gat));
  INV_X1    g582(.A(new_n603), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT54), .B1(new_n601), .B2(new_n602), .ZN(new_n785));
  OR2_X1    g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n607), .B1(new_n603), .B2(KEYINPUT54), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n786), .A2(KEYINPUT55), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n608), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n553), .B1(new_n552), .B2(new_n555), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n561), .A2(new_n563), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n531), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n568), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT55), .B1(new_n786), .B2(new_n788), .ZN(new_n795));
  OR4_X1    g594(.A1(new_n645), .A2(new_n790), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n789), .A2(new_n569), .A3(new_n608), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n797), .A2(new_n795), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n794), .B1(new_n608), .B2(new_n609), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n645), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n686), .ZN(new_n802));
  INV_X1    g601(.A(new_n569), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n632), .A2(new_n645), .A3(new_n803), .A4(new_n611), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n649), .A2(new_n359), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n807), .A2(new_n511), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n808), .A2(new_n212), .A3(new_n569), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n767), .A2(new_n464), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(G113gat), .B1(new_n811), .B2(new_n803), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n809), .A2(new_n812), .ZN(G1340gat));
  NAND3_X1  g612(.A1(new_n808), .A2(new_n210), .A3(new_n610), .ZN(new_n814));
  OAI21_X1  g613(.A(G120gat), .B1(new_n811), .B2(new_n687), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(G1341gat));
  AOI21_X1  g615(.A(G127gat), .B1(new_n808), .B2(new_n632), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n811), .A2(new_n215), .A3(new_n686), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n817), .A2(new_n818), .ZN(G1342gat));
  NAND4_X1  g618(.A1(new_n805), .A2(new_n217), .A3(new_n511), .A4(new_n806), .ZN(new_n820));
  OAI21_X1  g619(.A(KEYINPUT56), .B1(new_n820), .B2(new_n645), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT121), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n807), .A2(new_n675), .A3(new_n810), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(G134gat), .ZN(new_n825));
  OR3_X1    g624(.A1(new_n820), .A2(KEYINPUT56), .A3(new_n645), .ZN(new_n826));
  OAI211_X1 g625(.A(KEYINPUT121), .B(KEYINPUT56), .C1(new_n820), .C2(new_n645), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n823), .A2(new_n825), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT122), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n828), .B(new_n829), .ZN(G1343gat));
  NOR2_X1   g629(.A1(new_n382), .A2(new_n383), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n665), .A2(new_n806), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n789), .A2(new_n569), .A3(new_n608), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n786), .A2(KEYINPUT124), .A3(new_n788), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT124), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n784), .A2(new_n785), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n836), .B1(new_n837), .B2(new_n787), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT55), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n835), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n799), .B1(new_n834), .B2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT125), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n645), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AOI211_X1 g642(.A(KEYINPUT125), .B(new_n799), .C1(new_n834), .C2(new_n840), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n796), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n686), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n463), .B1(new_n846), .B2(new_n804), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT57), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n463), .B1(new_n802), .B2(new_n804), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  XNOR2_X1  g649(.A(KEYINPUT123), .B(KEYINPUT57), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n833), .B1(new_n848), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n832), .B1(new_n854), .B2(new_n569), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n665), .A2(new_n464), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(KEYINPUT126), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n856), .A2(KEYINPUT126), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n807), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n859), .A2(G141gat), .A3(new_n803), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT58), .B1(new_n855), .B2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(new_n833), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863));
  AOI211_X1 g662(.A(new_n863), .B(new_n463), .C1(new_n846), .C2(new_n804), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n849), .A2(new_n851), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n862), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n831), .B1(new_n866), .B2(new_n803), .ZN(new_n867));
  INV_X1    g666(.A(new_n860), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT58), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n861), .A2(new_n870), .ZN(G1344gat));
  OAI22_X1  g670(.A1(new_n847), .A2(KEYINPUT57), .B1(new_n850), .B2(new_n852), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n610), .A3(new_n862), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n854), .A2(new_n875), .A3(new_n610), .ZN(new_n876));
  INV_X1    g675(.A(new_n859), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n875), .B1(new_n877), .B2(new_n610), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n874), .B(new_n876), .C1(G148gat), .C2(new_n878), .ZN(G1345gat));
  AOI21_X1  g678(.A(G155gat), .B1(new_n877), .B2(new_n632), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n632), .A2(G155gat), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n880), .B1(new_n854), .B2(new_n881), .ZN(G1346gat));
  NOR2_X1   g681(.A1(new_n866), .A2(new_n645), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n377), .A2(new_n379), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n675), .A2(new_n884), .ZN(new_n885));
  OAI22_X1  g684(.A1(new_n883), .A2(new_n884), .B1(new_n859), .B2(new_n885), .ZN(G1347gat));
  NOR2_X1   g685(.A1(new_n650), .A2(new_n360), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n805), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n888), .A2(new_n507), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(new_n247), .A3(new_n569), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n805), .A2(new_n810), .A3(new_n887), .ZN(new_n891));
  OAI21_X1  g690(.A(G169gat), .B1(new_n891), .B2(new_n803), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(G1348gat));
  AOI21_X1  g692(.A(G176gat), .B1(new_n889), .B2(new_n610), .ZN(new_n894));
  INV_X1    g693(.A(new_n891), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n687), .A2(new_n249), .A3(new_n251), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(G1349gat));
  NAND3_X1  g696(.A1(new_n889), .A2(new_n632), .A3(new_n258), .ZN(new_n898));
  OAI21_X1  g697(.A(G183gat), .B1(new_n891), .B2(new_n686), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g700(.A(new_n259), .B1(new_n895), .B2(new_n675), .ZN(new_n902));
  OR3_X1    g701(.A1(new_n902), .A2(KEYINPUT127), .A3(KEYINPUT61), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n889), .A2(new_n259), .A3(new_n675), .ZN(new_n904));
  NAND2_X1  g703(.A1(KEYINPUT127), .A2(KEYINPUT61), .ZN(new_n905));
  OR2_X1    g704(.A1(KEYINPUT127), .A2(KEYINPUT61), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n902), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n903), .A2(new_n904), .A3(new_n907), .ZN(G1351gat));
  NAND3_X1  g707(.A1(new_n872), .A2(new_n665), .A3(new_n887), .ZN(new_n909));
  OAI21_X1  g708(.A(G197gat), .B1(new_n909), .B2(new_n803), .ZN(new_n910));
  OR2_X1    g709(.A1(new_n888), .A2(new_n856), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n569), .A2(new_n528), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(G1352gat));
  NOR3_X1   g712(.A1(new_n911), .A2(G204gat), .A3(new_n611), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT62), .ZN(new_n915));
  OAI21_X1  g714(.A(G204gat), .B1(new_n909), .B2(new_n687), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(G1353gat));
  OR3_X1    g716(.A1(new_n911), .A2(new_n686), .A3(new_n326), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n872), .A2(new_n632), .A3(new_n665), .A4(new_n887), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n919), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n920));
  AOI21_X1  g719(.A(KEYINPUT63), .B1(new_n919), .B2(G211gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(G1354gat));
  OAI21_X1  g721(.A(G218gat), .B1(new_n909), .B2(new_n645), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n645), .A2(G218gat), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n923), .B1(new_n911), .B2(new_n924), .ZN(G1355gat));
endmodule


