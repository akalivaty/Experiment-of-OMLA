//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 0 0 1 1 1 0 1 0 0 1 0 1 0 1 0 0 1 1 0 1 1 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(KEYINPUT64), .B1(new_n212), .B2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR3_X1   g0014(.A1(new_n212), .A2(KEYINPUT64), .A3(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n217), .B(G250), .C1(G257), .C2(G264), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT0), .ZN(new_n219));
  INV_X1    g0019(.A(new_n201), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(G50), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n223), .A2(new_n210), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n227));
  AND2_X1   g0027(.A1(new_n227), .A2(KEYINPUT65), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(KEYINPUT65), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n226), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  OR2_X1    g0030(.A1(new_n230), .A2(KEYINPUT66), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n230), .A2(KEYINPUT66), .ZN(new_n233));
  AOI22_X1  g0033(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n234));
  NAND2_X1  g0034(.A1(G50), .A2(G226), .ZN(new_n235));
  NAND2_X1  g0035(.A1(G116), .A2(G270), .ZN(new_n236));
  NAND4_X1  g0036(.A1(new_n233), .A2(new_n234), .A3(new_n235), .A4(new_n236), .ZN(new_n237));
  OAI21_X1  g0037(.A(new_n212), .B1(new_n232), .B2(new_n237), .ZN(new_n238));
  OAI211_X1 g0038(.A(new_n219), .B(new_n225), .C1(KEYINPUT1), .C2(new_n238), .ZN(new_n239));
  AOI21_X1  g0039(.A(new_n239), .B1(KEYINPUT1), .B2(new_n238), .ZN(G361));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G232), .ZN(new_n242));
  XOR2_X1   g0042(.A(KEYINPUT2), .B(G226), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G264), .B(G270), .Z(new_n245));
  XNOR2_X1  g0045(.A(G250), .B(G257), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G358));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XOR2_X1   g0049(.A(G107), .B(G116), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G50), .B(G68), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G58), .B(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  OAI21_X1  g0055(.A(KEYINPUT68), .B1(new_n210), .B2(G1), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT68), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(new_n209), .A3(G20), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(new_n202), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n223), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n261), .A2(new_n266), .B1(new_n202), .B2(new_n263), .ZN(new_n267));
  INV_X1    g0067(.A(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(G20), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT67), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G58), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT8), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT8), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G58), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n210), .A2(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT67), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n271), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G20), .A2(G33), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n265), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n267), .A2(KEYINPUT9), .A3(new_n283), .ZN(new_n284));
  XOR2_X1   g0084(.A(new_n284), .B(KEYINPUT72), .Z(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT3), .B(G33), .ZN(new_n286));
  INV_X1    g0086(.A(G1698), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n286), .A2(G222), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n286), .A2(G223), .A3(G1698), .ZN(new_n289));
  INV_X1    g0089(.A(G77), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n288), .B(new_n289), .C1(new_n290), .C2(new_n286), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n223), .B1(G33), .B2(G41), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G41), .ZN(new_n294));
  INV_X1    g0094(.A(G45), .ZN(new_n295));
  AOI21_X1  g0095(.A(G1), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(G33), .A2(G41), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n297), .A2(G1), .A3(G13), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n296), .A2(new_n298), .A3(G274), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n292), .A2(new_n296), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n300), .B1(G226), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n293), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G190), .ZN(new_n304));
  OR3_X1    g0104(.A1(new_n303), .A2(KEYINPUT73), .A3(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(KEYINPUT73), .B1(new_n303), .B2(new_n304), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT9), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n267), .A2(new_n283), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n308), .A2(new_n309), .B1(new_n303), .B2(G200), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n285), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT10), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT10), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n285), .A2(new_n313), .A3(new_n307), .A4(new_n310), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n271), .A2(G77), .A3(new_n278), .ZN(new_n316));
  INV_X1    g0116(.A(G68), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n280), .A2(G50), .B1(G20), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(KEYINPUT11), .B1(new_n319), .B2(new_n265), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n266), .A2(G68), .A3(new_n259), .ZN(new_n321));
  OAI21_X1  g0121(.A(KEYINPUT74), .B1(new_n262), .B2(G68), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT12), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n322), .A2(new_n323), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n321), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT11), .ZN(new_n327));
  INV_X1    g0127(.A(new_n265), .ZN(new_n328));
  AOI211_X1 g0128(.A(new_n327), .B(new_n328), .C1(new_n316), .C2(new_n318), .ZN(new_n329));
  NOR3_X1   g0129(.A1(new_n320), .A2(new_n326), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT14), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n268), .A2(KEYINPUT3), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT3), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G33), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n333), .A2(new_n335), .A3(G232), .A4(G1698), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n333), .A2(new_n335), .A3(G226), .A4(new_n287), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G33), .A2(G97), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n292), .ZN(new_n340));
  INV_X1    g0140(.A(G274), .ZN(new_n341));
  INV_X1    g0141(.A(new_n223), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n341), .B1(new_n342), .B2(new_n297), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n301), .A2(G238), .B1(new_n343), .B2(new_n296), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT13), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n340), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n345), .B1(new_n340), .B2(new_n344), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n332), .B(G169), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n340), .A2(new_n344), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT13), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n340), .A2(new_n344), .A3(new_n345), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n350), .A2(G179), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n350), .A2(new_n351), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n332), .B1(new_n354), .B2(G169), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n331), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(G200), .B1(new_n346), .B2(new_n347), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n350), .A2(G190), .A3(new_n351), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n358), .A2(new_n359), .A3(new_n330), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n303), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n309), .B1(new_n363), .B2(G169), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT69), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n365), .ZN(new_n367));
  INV_X1    g0167(.A(G179), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n366), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n273), .A2(new_n275), .A3(KEYINPUT70), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(KEYINPUT70), .B1(new_n273), .B2(new_n275), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n280), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  XOR2_X1   g0174(.A(KEYINPUT15), .B(G87), .Z(new_n375));
  AOI22_X1  g0175(.A1(new_n375), .A2(new_n269), .B1(G20), .B2(G77), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n265), .ZN(new_n378));
  INV_X1    g0178(.A(new_n266), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n259), .A2(G77), .ZN(new_n380));
  OAI22_X1  g0180(.A1(new_n379), .A2(new_n380), .B1(G77), .B2(new_n262), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n333), .A2(new_n335), .A3(G232), .A4(new_n287), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n333), .A2(new_n335), .A3(G238), .A4(G1698), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n384), .B(new_n385), .C1(new_n206), .C2(new_n286), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n292), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n298), .A2(G244), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n299), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(G169), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n390), .B1(new_n386), .B2(new_n292), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n368), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n383), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n392), .A2(G200), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n395), .A2(G190), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n398), .A2(new_n399), .A3(new_n378), .A4(new_n382), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  XNOR2_X1  g0201(.A(new_n401), .B(KEYINPUT71), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n315), .A2(new_n362), .A3(new_n370), .A4(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT80), .ZN(new_n404));
  INV_X1    g0204(.A(G223), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n405), .A2(G1698), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n406), .A2(new_n333), .A3(new_n335), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT77), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n286), .A2(G226), .A3(G1698), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G33), .A2(G87), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n406), .A2(new_n333), .A3(new_n335), .A4(KEYINPUT77), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n409), .A2(new_n410), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n292), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT78), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT78), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n413), .A2(new_n416), .A3(new_n292), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n301), .A2(G232), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n299), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n419), .A2(G190), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n415), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n300), .B1(G232), .B2(new_n301), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n414), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(G200), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n333), .A2(new_n335), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT7), .B1(new_n427), .B2(new_n210), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT7), .ZN(new_n429));
  AOI211_X1 g0229(.A(new_n429), .B(G20), .C1(new_n333), .C2(new_n335), .ZN(new_n430));
  OAI21_X1  g0230(.A(G68), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT75), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(new_n272), .B2(new_n317), .ZN(new_n433));
  NAND3_X1  g0233(.A1(KEYINPUT75), .A2(G58), .A3(G68), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n433), .A2(new_n220), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(G20), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT76), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n280), .A2(G159), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT76), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n435), .A2(new_n439), .A3(G20), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n431), .A2(new_n437), .A3(new_n438), .A4(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT16), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n429), .B1(new_n286), .B2(G20), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n427), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n446), .A2(G68), .B1(G159), .B2(new_n280), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n447), .A2(KEYINPUT16), .A3(new_n437), .A4(new_n440), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n443), .A2(new_n448), .A3(new_n265), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n259), .A2(new_n276), .ZN(new_n450));
  OAI22_X1  g0250(.A1(new_n379), .A2(new_n450), .B1(new_n262), .B2(new_n276), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  AND4_X1   g0252(.A1(KEYINPUT17), .A2(new_n426), .A3(new_n449), .A4(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n328), .B1(new_n441), .B2(new_n442), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n451), .B1(new_n454), .B2(new_n448), .ZN(new_n455));
  AOI21_X1  g0255(.A(KEYINPUT17), .B1(new_n455), .B2(new_n426), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n404), .B1(new_n453), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n426), .A2(new_n449), .A3(new_n452), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT17), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n455), .A2(KEYINPUT17), .A3(new_n426), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n460), .A2(KEYINPUT80), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n457), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n449), .A2(new_n452), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n415), .A2(new_n368), .A3(new_n417), .A4(new_n422), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n423), .A2(new_n393), .ZN(new_n466));
  AND2_X1   g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n464), .A2(new_n467), .A3(KEYINPUT18), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT79), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT79), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n464), .A2(new_n467), .A3(new_n470), .A4(KEYINPUT18), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT18), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n465), .A2(new_n466), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n472), .B1(new_n455), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n469), .A2(new_n471), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n463), .A2(new_n475), .ZN(new_n476));
  OR3_X1    g0276(.A1(new_n403), .A2(new_n476), .A3(KEYINPUT81), .ZN(new_n477));
  OAI21_X1  g0277(.A(KEYINPUT81), .B1(new_n403), .B2(new_n476), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n333), .A2(new_n335), .A3(G244), .A4(G1698), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n333), .A2(new_n335), .A3(G238), .A4(new_n287), .ZN(new_n481));
  INV_X1    g0281(.A(G116), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n480), .B(new_n481), .C1(new_n268), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n292), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n209), .A2(G45), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n298), .A2(G250), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n298), .A2(G274), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n486), .B1(new_n487), .B2(new_n485), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n484), .A2(G190), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT84), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n488), .B1(new_n483), .B2(new_n292), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT84), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n492), .A2(new_n493), .A3(G190), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n492), .A2(new_n424), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n375), .A2(new_n262), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT19), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n210), .B1(new_n338), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(G87), .B2(new_n207), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n333), .A2(new_n335), .A3(new_n210), .A4(G68), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n498), .B1(new_n277), .B2(new_n205), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n497), .B1(new_n503), .B2(new_n265), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n209), .A2(G33), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n262), .A2(new_n505), .A3(new_n223), .A4(new_n264), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G87), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n496), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n484), .A2(new_n489), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n393), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n507), .A2(new_n375), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n368), .A2(new_n492), .B1(new_n504), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n495), .A2(new_n510), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n280), .A2(G77), .ZN(new_n516));
  XNOR2_X1  g0316(.A(G97), .B(G107), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT6), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n518), .A2(new_n205), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n517), .A2(new_n518), .B1(new_n206), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n516), .B1(new_n520), .B2(new_n210), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n206), .B1(new_n444), .B2(new_n445), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n265), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n262), .A2(G97), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n524), .B1(new_n507), .B2(G97), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n333), .A2(new_n335), .A3(G244), .A4(new_n287), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT4), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n286), .A2(KEYINPUT4), .A3(G244), .A4(new_n287), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G283), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n286), .A2(G250), .A3(G1698), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n529), .A2(new_n530), .A3(new_n531), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n292), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n295), .A2(G1), .ZN(new_n535));
  XNOR2_X1  g0335(.A(KEYINPUT5), .B(G41), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n343), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AND2_X1   g0337(.A1(KEYINPUT5), .A2(G41), .ZN(new_n538));
  NOR2_X1   g0338(.A1(KEYINPUT5), .A2(G41), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n535), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n540), .A2(G257), .A3(new_n298), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT82), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT82), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n537), .A2(new_n541), .A3(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n534), .A2(new_n543), .A3(new_n368), .A4(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n526), .A2(new_n546), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n537), .A2(new_n541), .A3(new_n544), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n544), .B1(new_n537), .B2(new_n541), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(G169), .B1(new_n550), .B2(new_n534), .ZN(new_n551));
  OAI21_X1  g0351(.A(KEYINPUT83), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n526), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n534), .A2(new_n543), .A3(new_n545), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(G200), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n553), .B(new_n555), .C1(new_n304), .C2(new_n554), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n554), .A2(new_n393), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT83), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n557), .A2(new_n558), .A3(new_n526), .A4(new_n546), .ZN(new_n559));
  AND4_X1   g0359(.A1(new_n515), .A2(new_n552), .A3(new_n556), .A4(new_n559), .ZN(new_n560));
  OR2_X1    g0360(.A1(G250), .A2(G1698), .ZN(new_n561));
  INV_X1    g0361(.A(G257), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(G1698), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g0364(.A(KEYINPUT86), .B(G294), .ZN(new_n565));
  OAI22_X1  g0365(.A1(new_n564), .A2(new_n427), .B1(new_n565), .B2(new_n268), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT87), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n333), .A2(new_n561), .A3(new_n335), .A4(new_n563), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n569), .B(KEYINPUT87), .C1(new_n268), .C2(new_n565), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n568), .A2(new_n292), .A3(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n540), .A2(G264), .A3(new_n298), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n571), .A2(new_n304), .A3(new_n537), .A4(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n537), .ZN(new_n574));
  INV_X1    g0374(.A(new_n572), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n298), .B1(new_n566), .B2(new_n567), .ZN(new_n576));
  AOI211_X1 g0376(.A(new_n574), .B(new_n575), .C1(new_n576), .C2(new_n570), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n573), .B1(new_n577), .B2(G200), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT25), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(new_n262), .B2(G107), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  NOR3_X1   g0381(.A1(new_n262), .A2(new_n579), .A3(G107), .ZN(new_n582));
  OAI22_X1  g0382(.A1(new_n581), .A2(new_n582), .B1(new_n206), .B2(new_n506), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n333), .A2(new_n335), .A3(new_n210), .A4(G87), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT22), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT22), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n286), .A2(new_n586), .A3(new_n210), .A4(G87), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NOR3_X1   g0388(.A1(new_n268), .A2(new_n482), .A3(G20), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT23), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(new_n210), .B2(G107), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n589), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(KEYINPUT24), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT24), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n588), .A2(new_n596), .A3(new_n593), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n583), .B1(new_n598), .B2(new_n265), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n578), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n571), .A2(new_n537), .A3(new_n572), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n393), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n571), .A2(new_n368), .A3(new_n537), .A4(new_n572), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n328), .B1(new_n595), .B2(new_n597), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n602), .B(new_n603), .C1(new_n604), .C2(new_n583), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(KEYINPUT85), .A2(KEYINPUT21), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n540), .A2(G270), .A3(new_n298), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n287), .A2(G264), .ZN(new_n609));
  NOR2_X1   g0409(.A1(G257), .A2(G1698), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n611), .A2(new_n427), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n292), .B1(new_n286), .B2(G303), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n537), .B(new_n608), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(G169), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n263), .A2(new_n482), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n616), .B1(new_n506), .B2(new_n482), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n264), .A2(new_n223), .B1(G20), .B2(new_n482), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n531), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n619));
  AOI21_X1  g0419(.A(KEYINPUT20), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n618), .A2(KEYINPUT20), .A3(new_n619), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n617), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n607), .B1(new_n615), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n614), .A2(G200), .ZN(new_n625));
  INV_X1    g0425(.A(G303), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n298), .B1(new_n427), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n627), .B1(new_n427), .B2(new_n611), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n628), .A2(G190), .A3(new_n537), .A4(new_n608), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n625), .A2(new_n629), .A3(new_n623), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n614), .A2(new_n368), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n507), .A2(G116), .ZN(new_n632));
  INV_X1    g0432(.A(new_n622), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n632), .B(new_n616), .C1(new_n633), .C2(new_n620), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n607), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n634), .A2(G169), .A3(new_n614), .A4(new_n636), .ZN(new_n637));
  AND4_X1   g0437(.A1(new_n624), .A2(new_n630), .A3(new_n635), .A4(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n606), .A2(new_n639), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n479), .A2(new_n560), .A3(new_n640), .ZN(G372));
  INV_X1    g0441(.A(KEYINPUT26), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n552), .A2(new_n559), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n642), .B1(new_n643), .B2(new_n515), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT88), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n645), .B1(new_n511), .B2(new_n393), .ZN(new_n646));
  NOR3_X1   g0446(.A1(new_n492), .A2(KEYINPUT88), .A3(G169), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n514), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n495), .A2(new_n510), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n526), .A2(new_n546), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n649), .A2(new_n648), .A3(new_n650), .A4(new_n557), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n648), .B1(new_n651), .B2(KEYINPUT26), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n644), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n624), .A2(new_n635), .A3(new_n637), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n605), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n511), .A2(new_n645), .A3(new_n393), .ZN(new_n657));
  OAI21_X1  g0457(.A(KEYINPUT88), .B1(new_n492), .B2(G169), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n514), .A2(new_n659), .B1(new_n495), .B2(new_n510), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n656), .A2(new_n600), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n552), .A2(new_n556), .A3(new_n559), .ZN(new_n662));
  OAI21_X1  g0462(.A(KEYINPUT89), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n660), .A2(new_n600), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n552), .A2(new_n556), .A3(new_n559), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT89), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n664), .A2(new_n665), .A3(new_n666), .A4(new_n656), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n653), .A2(new_n663), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n479), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n370), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n356), .B1(new_n361), .B2(new_n397), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n463), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n468), .A2(new_n474), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n670), .B1(new_n674), .B2(new_n315), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n669), .A2(new_n675), .ZN(G369));
  NAND3_X1  g0476(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT90), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(G213), .ZN(new_n680));
  OR3_X1    g0480(.A1(new_n678), .A2(KEYINPUT91), .A3(KEYINPUT27), .ZN(new_n681));
  OAI21_X1  g0481(.A(KEYINPUT91), .B1(new_n678), .B2(KEYINPUT27), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n680), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G343), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(new_n623), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n654), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n639), .B2(new_n685), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n687), .A2(G330), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n599), .A2(new_n684), .ZN(new_n689));
  OAI22_X1  g0489(.A1(new_n606), .A2(new_n689), .B1(new_n605), .B2(new_n684), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n654), .A2(new_n684), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n693), .A2(new_n605), .A3(new_n600), .ZN(new_n694));
  INV_X1    g0494(.A(new_n684), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n605), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n691), .A2(new_n698), .ZN(G399));
  NOR2_X1   g0499(.A1(new_n216), .A2(G41), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n702));
  AND3_X1   g0502(.A1(new_n701), .A2(G1), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n703), .B1(new_n222), .B2(new_n700), .ZN(new_n704));
  XOR2_X1   g0504(.A(new_n704), .B(KEYINPUT28), .Z(new_n705));
  INV_X1    g0505(.A(new_n648), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n706), .B1(new_n651), .B2(KEYINPUT26), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n643), .A2(new_n642), .A3(new_n515), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n707), .B(new_n708), .C1(new_n661), .C2(new_n662), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n709), .A2(KEYINPUT29), .A3(new_n684), .ZN(new_n710));
  XOR2_X1   g0510(.A(new_n710), .B(KEYINPUT95), .Z(new_n711));
  NAND2_X1  g0511(.A1(new_n668), .A2(new_n684), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT94), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n712), .B(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n711), .B1(new_n714), .B2(KEYINPUT29), .ZN(new_n715));
  INV_X1    g0515(.A(G330), .ZN(new_n716));
  AND4_X1   g0516(.A1(new_n605), .A2(new_n600), .A3(new_n638), .A4(new_n684), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n560), .A2(new_n717), .A3(KEYINPUT93), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT93), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n552), .A2(new_n515), .A3(new_n556), .A4(new_n559), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n600), .A2(new_n605), .A3(new_n638), .A4(new_n684), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n719), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n614), .A2(new_n368), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n492), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n725), .A2(new_n554), .A3(new_n601), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(KEYINPUT92), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT30), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n631), .A2(new_n492), .A3(new_n572), .A4(new_n571), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n728), .B1(new_n729), .B2(new_n554), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n571), .A2(new_n492), .A3(new_n572), .ZN(new_n731));
  AND3_X1   g0531(.A1(new_n534), .A2(new_n543), .A3(new_n545), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n731), .A2(new_n732), .A3(KEYINPUT30), .A4(new_n631), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT92), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n725), .A2(new_n601), .A3(new_n554), .A4(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n727), .A2(new_n730), .A3(new_n733), .A4(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(KEYINPUT31), .B1(new_n736), .B2(new_n695), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n730), .A2(new_n733), .A3(new_n726), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n738), .A2(KEYINPUT31), .A3(new_n695), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n716), .B1(new_n723), .B2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n715), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(KEYINPUT96), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT96), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n715), .A2(new_n745), .A3(new_n742), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n705), .B1(new_n747), .B2(G1), .ZN(G364));
  AND2_X1   g0548(.A1(new_n210), .A2(G13), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n209), .B1(new_n749), .B2(G45), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n700), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n688), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(G330), .B2(new_n687), .ZN(new_n754));
  INV_X1    g0554(.A(new_n752), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n223), .B1(G20), .B2(new_n393), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n304), .A2(G179), .A3(G200), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n210), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n205), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n210), .A2(new_n368), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n424), .A2(G190), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n760), .B1(G68), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT97), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n304), .A2(new_n424), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n761), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G190), .A2(G200), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n761), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI22_X1  g0572(.A1(G50), .A2(new_n769), .B1(new_n772), .B2(G77), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n761), .A2(G190), .A3(new_n424), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n210), .A2(G179), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n767), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n775), .A2(G58), .B1(new_n778), .B2(G87), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT32), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n776), .A2(new_n770), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n780), .B1(new_n782), .B2(G159), .ZN(new_n783));
  INV_X1    g0583(.A(G159), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n781), .A2(KEYINPUT32), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n776), .A2(new_n762), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n206), .ZN(new_n787));
  NOR4_X1   g0587(.A1(new_n783), .A2(new_n785), .A3(new_n787), .A4(new_n427), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n766), .A2(new_n773), .A3(new_n779), .A4(new_n788), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n775), .A2(G322), .B1(new_n782), .B2(G329), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n286), .B1(new_n769), .B2(G326), .ZN(new_n791));
  AND2_X1   g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI22_X1  g0592(.A1(G311), .A2(new_n772), .B1(new_n778), .B2(G303), .ZN(new_n793));
  XNOR2_X1  g0593(.A(KEYINPUT33), .B(G317), .ZN(new_n794));
  INV_X1    g0594(.A(new_n786), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n764), .A2(new_n794), .B1(new_n795), .B2(G283), .ZN(new_n796));
  INV_X1    g0596(.A(new_n759), .ZN(new_n797));
  INV_X1    g0597(.A(new_n565), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n792), .A2(new_n793), .A3(new_n796), .A4(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n757), .B1(new_n789), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n217), .A2(G355), .A3(new_n286), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n216), .A2(new_n286), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(G45), .B2(new_n221), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n254), .A2(G45), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n802), .B1(G116), .B2(new_n217), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(G13), .A2(G33), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(G20), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n756), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n755), .B(new_n801), .C1(new_n806), .C2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n809), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n687), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n754), .A2(new_n813), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT98), .Z(G396));
  INV_X1    g0615(.A(KEYINPUT102), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n328), .B1(new_n374), .B2(new_n376), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n817), .A2(new_n381), .B1(new_n395), .B2(G169), .ZN(new_n818));
  INV_X1    g0618(.A(new_n396), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n816), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n383), .A2(new_n394), .A3(KEYINPUT102), .A4(new_n396), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n683), .A2(new_n383), .A3(G343), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n820), .A2(new_n821), .A3(new_n822), .A4(new_n400), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n397), .A2(new_n684), .ZN(new_n824));
  AOI21_X1  g0624(.A(KEYINPUT103), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n823), .A2(new_n824), .A3(KEYINPUT103), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n668), .A2(new_n684), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n714), .B2(new_n828), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n752), .B1(new_n830), .B2(new_n742), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n742), .B2(new_n830), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n756), .A2(new_n807), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(KEYINPUT99), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n775), .A2(G294), .B1(new_n764), .B2(G283), .ZN(new_n835));
  AOI22_X1  g0635(.A1(G87), .A2(new_n795), .B1(new_n782), .B2(G311), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n427), .B1(new_n768), .B2(new_n626), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n206), .A2(new_n777), .B1(new_n771), .B2(new_n482), .ZN(new_n839));
  NOR4_X1   g0639(.A1(new_n837), .A2(new_n760), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(G137), .ZN(new_n841));
  INV_X1    g0641(.A(G150), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n768), .A2(new_n841), .B1(new_n763), .B2(new_n842), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT100), .ZN(new_n844));
  INV_X1    g0644(.A(G143), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n844), .B1(new_n845), .B2(new_n774), .C1(new_n784), .C2(new_n771), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT34), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n286), .B1(new_n777), .B2(new_n202), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n795), .A2(G68), .ZN(new_n849));
  INV_X1    g0649(.A(G132), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n849), .B1(new_n850), .B2(new_n781), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n848), .B(new_n851), .C1(G58), .C2(new_n797), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n840), .B1(new_n847), .B2(new_n852), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n752), .B1(G77), .B2(new_n834), .C1(new_n853), .C2(new_n757), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(KEYINPUT101), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n808), .B2(new_n828), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n832), .A2(new_n856), .ZN(G384));
  INV_X1    g0657(.A(new_n520), .ZN(new_n858));
  OR2_X1    g0658(.A1(new_n858), .A2(KEYINPUT35), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(KEYINPUT35), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n859), .A2(G116), .A3(new_n224), .A4(new_n860), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n861), .B(KEYINPUT36), .Z(new_n862));
  NAND4_X1  g0662(.A1(new_n222), .A2(G77), .A3(new_n433), .A4(new_n434), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n202), .A2(G68), .ZN(new_n864));
  AOI211_X1 g0664(.A(new_n209), .B(G13), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n479), .B(new_n711), .C1(new_n714), .C2(KEYINPUT29), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n675), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT39), .ZN(new_n869));
  XOR2_X1   g0669(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n464), .A2(new_n683), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n453), .A2(new_n456), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n872), .B1(new_n873), .B2(new_n673), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n464), .A2(new_n467), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n875), .A2(new_n872), .A3(new_n458), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(KEYINPUT37), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT37), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n875), .A2(new_n872), .A3(new_n878), .A4(new_n458), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT106), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n874), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n877), .A2(KEYINPUT106), .A3(new_n879), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n871), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n872), .B1(new_n463), .B2(new_n475), .ZN(new_n885));
  INV_X1    g0685(.A(new_n880), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT38), .ZN(new_n887));
  NOR3_X1   g0687(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n869), .B1(new_n884), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n357), .A2(new_n684), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n887), .B1(new_n885), .B2(new_n886), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT18), .B1(new_n464), .B2(new_n467), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(KEYINPUT79), .B2(new_n468), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n894), .A2(new_n471), .B1(new_n457), .B2(new_n462), .ZN(new_n895));
  OAI211_X1 g0695(.A(KEYINPUT38), .B(new_n880), .C1(new_n895), .C2(new_n872), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n892), .A2(new_n896), .A3(KEYINPUT39), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n889), .A2(new_n891), .A3(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n673), .A2(new_n683), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n684), .A2(new_n330), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n356), .A2(new_n360), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(G169), .B1(new_n346), .B2(new_n347), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(KEYINPUT14), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n360), .A2(new_n904), .A3(new_n352), .A4(new_n348), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT104), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n905), .A2(new_n906), .A3(new_n900), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n902), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n906), .B1(new_n905), .B2(new_n900), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n820), .A2(new_n821), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n684), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n910), .B1(new_n829), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n892), .A2(new_n896), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n899), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n898), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n868), .B(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT40), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n892), .A2(new_n896), .A3(new_n918), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n736), .A2(KEYINPUT31), .A3(new_n695), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n920), .A2(new_n737), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n723), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n828), .B1(new_n908), .B2(new_n909), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT107), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n924), .A2(new_n918), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n922), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n919), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT93), .B1(new_n560), .B2(new_n717), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n720), .A2(new_n721), .A3(new_n719), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n921), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n823), .A2(new_n824), .A3(KEYINPUT103), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n931), .A2(new_n825), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n902), .A2(new_n907), .ZN(new_n933));
  INV_X1    g0733(.A(new_n909), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n924), .B1(new_n930), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n880), .A2(new_n881), .ZN(new_n937));
  INV_X1    g0737(.A(new_n874), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n937), .A2(new_n883), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n870), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n936), .B1(new_n940), .B2(new_n896), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n927), .B1(new_n941), .B2(new_n918), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n942), .A2(new_n479), .A3(new_n930), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n923), .B1(new_n723), .B2(new_n921), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n884), .A2(new_n888), .B1(new_n944), .B2(new_n924), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n945), .A2(KEYINPUT40), .B1(new_n919), .B2(new_n926), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n479), .A2(new_n930), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n943), .A2(G330), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n917), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n209), .B2(new_n749), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n917), .A2(new_n949), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n866), .B1(new_n951), .B2(new_n952), .ZN(G367));
  NAND3_X1  g0753(.A1(new_n778), .A2(KEYINPUT46), .A3(G116), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT46), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n777), .B2(new_n482), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n954), .B(new_n956), .C1(new_n565), .C2(new_n763), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT111), .Z(new_n958));
  INV_X1    g0758(.A(G317), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n427), .B1(new_n781), .B2(new_n959), .C1(new_n205), .C2(new_n786), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT112), .Z(new_n961));
  INV_X1    g0761(.A(G283), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n771), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(G311), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n774), .A2(new_n626), .B1(new_n768), .B2(new_n964), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n963), .B(new_n965), .C1(G107), .C2(new_n797), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n961), .A2(new_n966), .ZN(new_n967));
  AOI22_X1  g0767(.A1(G50), .A2(new_n772), .B1(new_n782), .B2(G137), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n968), .B1(new_n272), .B2(new_n777), .C1(new_n784), .C2(new_n763), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n797), .A2(G68), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n970), .B1(new_n768), .B2(new_n845), .C1(new_n842), .C2(new_n774), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n795), .A2(G77), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n286), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT113), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n958), .A2(new_n967), .B1(new_n972), .B2(new_n975), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT47), .Z(new_n977));
  NOR2_X1   g0777(.A1(new_n977), .A2(new_n757), .ZN(new_n978));
  INV_X1    g0778(.A(new_n803), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n979), .A2(new_n247), .ZN(new_n980));
  INV_X1    g0780(.A(new_n810), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(new_n216), .B2(new_n375), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n755), .B(new_n978), .C1(new_n980), .C2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n695), .A2(new_n509), .ZN(new_n984));
  MUX2_X1   g0784(.A(new_n706), .B(new_n660), .S(new_n984), .Z(new_n985));
  OAI21_X1  g0785(.A(new_n983), .B1(new_n812), .B2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n746), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n745), .B1(new_n715), .B2(new_n742), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n665), .B1(new_n553), .B2(new_n684), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n695), .A2(new_n650), .A3(new_n557), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n698), .ZN(new_n992));
  XOR2_X1   g0792(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n993));
  XNOR2_X1  g0793(.A(new_n992), .B(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n991), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n995), .A2(KEYINPUT44), .A3(new_n697), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT44), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n991), .B2(new_n698), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n996), .A2(KEYINPUT109), .A3(new_n998), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n998), .A2(KEYINPUT109), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n994), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n691), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n690), .A2(new_n693), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT110), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n694), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(new_n1005), .B2(new_n1004), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(new_n688), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n987), .A2(new_n988), .B1(new_n1003), .B2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n700), .B(KEYINPUT41), .Z(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n751), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n995), .A2(new_n694), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT42), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n995), .A2(new_n605), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n684), .B1(new_n1015), .B2(new_n643), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n1014), .A2(new_n1016), .B1(KEYINPUT43), .B2(new_n985), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n985), .A2(KEYINPUT43), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n995), .A2(new_n691), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1019), .A2(new_n1022), .A3(new_n1020), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n986), .B1(new_n1012), .B2(new_n1026), .ZN(G387));
  INV_X1    g0827(.A(new_n1008), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n747), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n744), .A2(new_n746), .A3(new_n1008), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1029), .A2(new_n700), .A3(new_n1030), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n690), .A2(new_n812), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n217), .A2(new_n286), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n1033), .A2(new_n702), .B1(G107), .B2(new_n217), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n372), .A2(new_n373), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n202), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT50), .Z(new_n1037));
  AOI21_X1  g0837(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1037), .A2(new_n702), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n979), .B1(new_n244), .B2(G45), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1034), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n752), .B1(new_n1041), .B2(new_n981), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n317), .A2(new_n771), .B1(new_n777), .B2(new_n290), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n427), .B(new_n1043), .C1(G97), .C2(new_n795), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n769), .A2(G159), .B1(new_n782), .B2(G150), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n775), .A2(G50), .B1(new_n764), .B2(new_n276), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n797), .A2(new_n375), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n797), .A2(G283), .B1(new_n778), .B2(new_n798), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G322), .A2(new_n769), .B1(new_n764), .B2(G311), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n626), .B2(new_n771), .C1(new_n959), .C2(new_n774), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT48), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1049), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT114), .Z(new_n1054));
  NAND2_X1  g0854(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1054), .A2(KEYINPUT49), .A3(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n286), .B1(new_n782), .B2(G326), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1056), .B(new_n1057), .C1(new_n482), .C2(new_n786), .ZN(new_n1058));
  AOI21_X1  g0858(.A(KEYINPUT49), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1048), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1042), .B1(new_n1060), .B2(new_n756), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n1028), .A2(new_n751), .B1(new_n1032), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1031), .A2(new_n1062), .ZN(G393));
  INV_X1    g0863(.A(new_n1003), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n751), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n803), .A2(new_n251), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n810), .B1(new_n217), .B2(new_n205), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n752), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n774), .A2(new_n964), .B1(new_n768), .B2(new_n959), .ZN(new_n1069));
  XOR2_X1   g0869(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n1070));
  XOR2_X1   g0870(.A(new_n1069), .B(new_n1070), .Z(new_n1071));
  AOI211_X1 g0871(.A(new_n286), .B(new_n787), .C1(G116), .C2(new_n797), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(G294), .A2(new_n772), .B1(new_n778), .B2(G283), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G303), .A2(new_n764), .B1(new_n782), .B2(G322), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n774), .A2(new_n784), .B1(new_n768), .B2(new_n842), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT51), .Z(new_n1077));
  OAI22_X1  g0877(.A1(new_n202), .A2(new_n763), .B1(new_n777), .B2(new_n317), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(G143), .B2(new_n782), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1035), .A2(new_n772), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n759), .A2(new_n290), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n427), .B1(new_n795), .B2(G87), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1079), .A2(new_n1080), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n1071), .A2(new_n1075), .B1(new_n1077), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1068), .B1(new_n1085), .B2(new_n756), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n991), .B2(new_n812), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1064), .B(new_n1028), .C1(new_n987), .C2(new_n988), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n700), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1064), .B1(new_n747), .B2(new_n1028), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1065), .B(new_n1087), .C1(new_n1089), .C2(new_n1090), .ZN(G390));
  AND3_X1   g0891(.A1(new_n930), .A2(G330), .A3(new_n935), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n829), .A2(new_n912), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n910), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n889), .A2(new_n897), .B1(new_n1095), .B2(new_n890), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n884), .A2(new_n888), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n709), .A2(new_n828), .A3(new_n684), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n1098), .A2(new_n912), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1099), .A2(new_n910), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n890), .B(KEYINPUT116), .ZN(new_n1101));
  NOR3_X1   g0901(.A1(new_n1097), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1092), .B1(new_n1096), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(KEYINPUT39), .B1(new_n940), .B2(new_n896), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n897), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n1104), .A2(new_n1105), .B1(new_n891), .B2(new_n913), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1101), .B1(new_n940), .B2(new_n896), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n910), .B2(new_n1099), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n716), .B(new_n932), .C1(new_n723), .C2(new_n740), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n1094), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1106), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1103), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n479), .A2(G330), .A3(new_n930), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n867), .A2(new_n675), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1110), .A2(new_n1099), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n922), .A2(new_n716), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1094), .B1(new_n1117), .B2(new_n828), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT118), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1093), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n740), .B1(new_n928), .B2(new_n929), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1123), .A2(G330), .A3(new_n828), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n910), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1092), .B1(new_n1125), .B2(KEYINPUT117), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT117), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1124), .A2(new_n1127), .A3(new_n910), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n1121), .B(new_n1122), .C1(new_n1126), .C2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(KEYINPUT117), .B1(new_n1109), .B2(new_n1094), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n930), .A2(G330), .A3(new_n935), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1130), .A2(new_n1131), .A3(new_n1128), .ZN(new_n1132));
  AOI21_X1  g0932(.A(KEYINPUT118), .B1(new_n1132), .B2(new_n1093), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1120), .B1(new_n1129), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1112), .A2(new_n1115), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1103), .A2(new_n1111), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1094), .B1(new_n741), .B2(new_n828), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1131), .B1(new_n1137), .B2(new_n1127), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1128), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1093), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n1121), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1132), .A2(KEYINPUT118), .A3(new_n1093), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1119), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1136), .B1(new_n1143), .B2(new_n1114), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1135), .A2(new_n1144), .A3(new_n700), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n807), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n752), .B1(new_n276), .B2(new_n834), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n777), .A2(new_n842), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1148), .B(KEYINPUT53), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n775), .A2(G132), .B1(new_n782), .B2(G125), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(KEYINPUT54), .B(G143), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1149), .B(new_n1150), .C1(new_n771), .C2(new_n1151), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(G128), .A2(new_n769), .B1(new_n764), .B2(G137), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n427), .B1(new_n795), .B2(G50), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1153), .B(new_n1154), .C1(new_n784), .C2(new_n759), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n775), .A2(G116), .B1(new_n782), .B2(G294), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n1156), .B1(new_n205), .B2(new_n771), .C1(new_n206), .C2(new_n763), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n286), .B1(new_n778), .B2(G87), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n769), .A2(G283), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1082), .A2(new_n1158), .A3(new_n849), .A4(new_n1159), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n1152), .A2(new_n1155), .B1(new_n1157), .B2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1147), .B1(new_n1161), .B2(new_n756), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n1112), .A2(new_n751), .B1(new_n1146), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1145), .A2(new_n1163), .ZN(G378));
  XOR2_X1   g0964(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1165));
  NAND2_X1  g0965(.A1(new_n315), .A2(new_n370), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n683), .A2(new_n309), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT120), .Z(new_n1168));
  NOR2_X1   g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1165), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1171), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1165), .ZN(new_n1174));
  NOR3_X1   g0974(.A1(new_n1173), .A2(new_n1169), .A3(new_n1174), .ZN(new_n1175));
  OR2_X1    g0975(.A1(new_n1172), .A2(new_n1175), .ZN(new_n1176));
  NOR3_X1   g0976(.A1(new_n946), .A2(new_n716), .A3(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1172), .A2(new_n1175), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n942), .B2(G330), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n916), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT121), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1176), .B1(new_n946), .B2(new_n716), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n942), .A2(G330), .A3(new_n1178), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n916), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1180), .A2(new_n1181), .A3(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1115), .B1(new_n1143), .B2(new_n1136), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1182), .A2(new_n1184), .A3(new_n1183), .A4(KEYINPUT121), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT57), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1190), .B1(new_n1180), .B2(new_n1185), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n701), .B1(new_n1192), .B2(new_n1187), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1186), .A2(new_n751), .A3(new_n1188), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n752), .B1(G50), .B2(new_n834), .ZN(new_n1196));
  INV_X1    g0996(.A(G128), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n774), .A2(new_n1197), .B1(new_n763), .B2(new_n850), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(G125), .A2(new_n769), .B1(new_n772), .B2(G137), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n777), .B2(new_n1151), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1198), .B(new_n1200), .C1(G150), .C2(new_n797), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT59), .ZN(new_n1202));
  OR2_X1    g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n268), .B(new_n294), .C1(new_n786), .C2(new_n784), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(G124), .B2(new_n782), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1203), .A2(new_n1204), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n427), .A2(new_n294), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(G77), .B2(new_n778), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT119), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(G116), .A2(new_n769), .B1(new_n772), .B2(new_n375), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1211), .B1(new_n272), .B2(new_n786), .C1(new_n206), .C2(new_n774), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n970), .B1(new_n205), .B2(new_n763), .C1(new_n962), .C2(new_n781), .ZN(new_n1213));
  NOR3_X1   g1013(.A1(new_n1210), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n1214), .A2(KEYINPUT58), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(KEYINPUT58), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1208), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1207), .A2(new_n1215), .A3(new_n1216), .A4(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1196), .B1(new_n1218), .B2(new_n756), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1219), .B1(new_n1178), .B2(new_n808), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1195), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1194), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT122), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1221), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(KEYINPUT122), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1225), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(G375));
  NAND2_X1  g1029(.A1(new_n910), .A2(new_n807), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n752), .B1(G68), .B2(new_n834), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n774), .A2(new_n841), .B1(new_n771), .B2(new_n842), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n427), .B(new_n1232), .C1(G58), .C2(new_n795), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n768), .A2(new_n850), .B1(new_n763), .B2(new_n1151), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n777), .A2(new_n784), .B1(new_n781), .B2(new_n1197), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1233), .B(new_n1236), .C1(new_n202), .C2(new_n759), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(G116), .A2(new_n764), .B1(new_n782), .B2(G303), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1238), .B1(new_n205), .B2(new_n777), .C1(new_n962), .C2(new_n774), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(G294), .A2(new_n769), .B1(new_n772), .B2(G107), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1240), .A2(new_n427), .A3(new_n973), .A4(new_n1047), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1237), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n1242), .A2(KEYINPUT123), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n757), .B1(new_n1242), .B2(KEYINPUT123), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1231), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n1134), .A2(new_n751), .B1(new_n1230), .B2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1011), .B1(new_n1143), .B2(new_n1114), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1114), .B(new_n1120), .C1(new_n1129), .C2(new_n1133), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1246), .B1(new_n1247), .B2(new_n1249), .ZN(G381));
  INV_X1    g1050(.A(G378), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1065), .A2(new_n1087), .ZN(new_n1252));
  AND2_X1   g1052(.A1(new_n1088), .A2(new_n700), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1090), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1252), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1255), .A2(new_n832), .A3(new_n856), .ZN(new_n1256));
  INV_X1    g1056(.A(G396), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1031), .A2(new_n1257), .A3(new_n1062), .ZN(new_n1258));
  NOR4_X1   g1058(.A1(new_n1256), .A2(G387), .A3(G381), .A4(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1228), .A2(new_n1251), .A3(new_n1259), .ZN(G407));
  INV_X1    g1060(.A(G343), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(G213), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1228), .A2(new_n1251), .A3(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(G407), .A2(new_n1264), .A3(G213), .ZN(G409));
  NAND3_X1  g1065(.A1(new_n1194), .A2(G378), .A3(new_n1222), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1186), .A2(new_n1187), .A3(new_n1011), .A4(new_n1188), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1220), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1180), .A2(new_n1185), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1268), .B1(new_n1269), .B2(new_n751), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1267), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1251), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1266), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT124), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT60), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1275), .B1(new_n1134), .B2(new_n1115), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1274), .B1(new_n1276), .B2(new_n1249), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1114), .B1(new_n1278), .B2(new_n1120), .ZN(new_n1279));
  OAI211_X1 g1079(.A(KEYINPUT124), .B(new_n1248), .C1(new_n1279), .C2(new_n1275), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n701), .B1(new_n1249), .B2(KEYINPUT60), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1277), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1246), .B1(KEYINPUT125), .B2(G384), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1282), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1282), .A2(new_n1286), .A3(new_n1284), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1273), .A2(new_n1290), .A3(new_n1262), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(KEYINPUT62), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT61), .ZN(new_n1293));
  INV_X1    g1093(.A(G2897), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1262), .A2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1282), .A2(new_n1286), .A3(new_n1284), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1286), .B1(new_n1282), .B2(new_n1284), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1296), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1288), .A2(new_n1295), .A3(new_n1289), .ZN(new_n1300));
  AOI21_X1  g1100(.A(G378), .B1(new_n1267), .B2(new_n1270), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1301), .B1(new_n1226), .B2(G378), .ZN(new_n1302));
  OAI211_X1 g1102(.A(new_n1299), .B(new_n1300), .C1(new_n1302), .C2(new_n1263), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT62), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1273), .A2(new_n1290), .A3(new_n1304), .A4(new_n1262), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1292), .A2(new_n1293), .A3(new_n1303), .A4(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(new_n750), .ZN(new_n1308));
  AND2_X1   g1108(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1310), .A2(G390), .A3(new_n986), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1255), .A2(G387), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1257), .B1(new_n1031), .B2(new_n1062), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  AOI22_X1  g1114(.A1(new_n1311), .A2(new_n1312), .B1(new_n1258), .B2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  AND3_X1   g1116(.A1(new_n1031), .A2(new_n1257), .A3(new_n1062), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1317), .A2(new_n1313), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1318), .A2(new_n1311), .A3(new_n1312), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1316), .A2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1306), .A2(new_n1320), .ZN(new_n1321));
  NOR3_X1   g1121(.A1(new_n1297), .A2(new_n1298), .A3(new_n1296), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1295), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1323));
  OAI21_X1  g1123(.A(KEYINPUT126), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT126), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1299), .A2(new_n1300), .A3(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1273), .A2(new_n1262), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1324), .A2(new_n1326), .A3(new_n1327), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1273), .A2(new_n1290), .A3(KEYINPUT63), .A4(new_n1262), .ZN(new_n1329));
  AND3_X1   g1129(.A1(new_n1318), .A2(new_n1311), .A3(new_n1312), .ZN(new_n1330));
  NOR3_X1   g1130(.A1(new_n1330), .A2(new_n1315), .A3(KEYINPUT61), .ZN(new_n1331));
  AND2_X1   g1131(.A1(new_n1329), .A2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT63), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1291), .A2(new_n1333), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1328), .A2(new_n1332), .A3(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1321), .A2(new_n1335), .ZN(G405));
  OAI211_X1 g1136(.A(KEYINPUT127), .B(new_n1266), .C1(new_n1228), .C2(G378), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT127), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1225), .A2(new_n1227), .A3(new_n1338), .A4(new_n1251), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1337), .A2(new_n1339), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1320), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1316), .A2(new_n1290), .A3(new_n1319), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1340), .A2(new_n1343), .ZN(new_n1344));
  NAND4_X1  g1144(.A1(new_n1337), .A2(new_n1341), .A3(new_n1339), .A4(new_n1342), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1344), .A2(new_n1345), .ZN(G402));
endmodule


