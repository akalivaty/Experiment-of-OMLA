//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 1 0 0 0 0 0 0 1 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n836, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n205), .B(new_n206), .Z(new_n207));
  XNOR2_X1  g006(.A(G15gat), .B(G22gat), .ZN(new_n208));
  AND2_X1   g007(.A1(KEYINPUT88), .A2(G1gat), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT16), .B1(KEYINPUT88), .B2(G1gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n211), .B(KEYINPUT89), .C1(G1gat), .C2(new_n208), .ZN(new_n212));
  XOR2_X1   g011(.A(new_n212), .B(G8gat), .Z(new_n213));
  OAI21_X1  g012(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  NOR3_X1   g014(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(G29gat), .A2(G36gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT87), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(KEYINPUT87), .B1(G29gat), .B2(G36gat), .ZN(new_n220));
  OAI22_X1  g019(.A1(new_n215), .A2(new_n216), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT15), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI221_X1 g022(.A(KEYINPUT15), .B1(new_n219), .B2(new_n220), .C1(new_n215), .C2(new_n216), .ZN(new_n224));
  XNOR2_X1  g023(.A(G43gat), .B(G50gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  OR3_X1    g025(.A1(new_n221), .A2(new_n222), .A3(new_n225), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT17), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n228), .B1(new_n226), .B2(new_n227), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n213), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(G229gat), .A2(G233gat), .ZN(new_n233));
  OR2_X1    g032(.A1(new_n212), .A2(G8gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n212), .A2(G8gat), .ZN(new_n235));
  AOI22_X1  g034(.A1(new_n234), .A2(new_n235), .B1(new_n226), .B2(new_n227), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n232), .A2(new_n233), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT18), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT91), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n226), .A2(new_n227), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT17), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(new_n229), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n236), .B1(new_n243), .B2(new_n213), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT91), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n244), .A2(new_n245), .A3(KEYINPUT18), .A4(new_n233), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n240), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT90), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n238), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n244), .A2(KEYINPUT90), .A3(new_n233), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n249), .A2(new_n250), .A3(new_n239), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n213), .A2(new_n226), .A3(new_n227), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(new_n237), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n233), .B(KEYINPUT13), .Z(new_n254));
  AND2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  AND4_X1   g055(.A1(new_n207), .A2(new_n247), .A3(new_n251), .A4(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n255), .B1(new_n240), .B2(new_n246), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n207), .B1(new_n258), .B2(new_n251), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(G78gat), .B(G106gat), .Z(new_n261));
  XNOR2_X1  g060(.A(KEYINPUT31), .B(G50gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n261), .B(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n263), .A2(KEYINPUT81), .ZN(new_n264));
  AND2_X1   g063(.A1(G155gat), .A2(G162gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(G155gat), .A2(G162gat), .ZN(new_n266));
  OAI21_X1  g065(.A(KEYINPUT73), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G155gat), .ZN(new_n268));
  INV_X1    g067(.A(G162gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT73), .ZN(new_n271));
  NAND2_X1  g070(.A1(G155gat), .A2(G162gat), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G141gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(G148gat), .ZN(new_n276));
  INV_X1    g075(.A(G148gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(G141gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n272), .A2(KEYINPUT2), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n274), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT3), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT74), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n284), .B1(new_n277), .B2(G141gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n275), .A2(KEYINPUT74), .A3(G148gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(new_n278), .A3(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n272), .B1(new_n270), .B2(KEYINPUT2), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n282), .A2(new_n283), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT29), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AND2_X1   g091(.A1(G211gat), .A2(G218gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(G211gat), .A2(G218gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AND2_X1   g094(.A1(G197gat), .A2(G204gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(G197gat), .A2(G204gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n295), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(G211gat), .B(G218gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(G197gat), .B(G204gat), .ZN(new_n302));
  INV_X1    g101(.A(new_n299), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n300), .A2(new_n304), .A3(KEYINPUT69), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT69), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n306), .B(new_n295), .C1(new_n298), .C2(new_n299), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n308), .ZN(new_n309));
  AOI22_X1  g108(.A1(new_n274), .A2(new_n281), .B1(new_n287), .B2(new_n288), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT29), .B1(new_n300), .B2(new_n304), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n311), .B1(KEYINPUT3), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(G228gat), .A2(G233gat), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n264), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n263), .A2(KEYINPUT81), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(G22gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n308), .A2(KEYINPUT70), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT70), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n305), .A2(new_n320), .A3(new_n307), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n315), .B1(new_n322), .B2(new_n292), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n305), .A2(new_n291), .A3(new_n307), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT79), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT3), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n305), .A2(new_n307), .A3(KEYINPUT79), .A4(new_n291), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n310), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT80), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n323), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n324), .A2(new_n325), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n331), .A2(new_n283), .A3(new_n327), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(new_n311), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n333), .A2(KEYINPUT80), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n316), .B(new_n318), .C1(new_n330), .C2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n333), .A2(KEYINPUT80), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n328), .A2(new_n329), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n338), .A3(new_n323), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n318), .B1(new_n339), .B2(new_n316), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n308), .ZN(new_n342));
  INV_X1    g141(.A(G226gat), .ZN(new_n343));
  INV_X1    g142(.A(G233gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G183gat), .A2(G190gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT24), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT24), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n349), .A2(G183gat), .A3(G190gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g150(.A1(G183gat), .A2(G190gat), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(G169gat), .ZN(new_n355));
  INV_X1    g154(.A(G176gat), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(new_n356), .A3(KEYINPUT23), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT23), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n358), .B1(G169gat), .B2(G176gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(G169gat), .A2(G176gat), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n357), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n354), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT25), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT64), .ZN(new_n364));
  INV_X1    g163(.A(G190gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(G183gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(KEYINPUT64), .A2(G190gat), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n351), .A2(new_n369), .ZN(new_n370));
  AND4_X1   g169(.A1(KEYINPUT25), .A2(new_n357), .A3(new_n359), .A4(new_n360), .ZN(new_n371));
  AOI22_X1  g170(.A1(new_n362), .A2(new_n363), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(G169gat), .A2(G176gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT26), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT26), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n375), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n374), .B(new_n347), .C1(new_n376), .C2(new_n373), .ZN(new_n377));
  AND2_X1   g176(.A1(KEYINPUT64), .A2(G190gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(KEYINPUT64), .A2(G190gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT27), .B(G183gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT28), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n380), .A2(new_n381), .A3(KEYINPUT28), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n377), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(KEYINPUT71), .B1(new_n372), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n370), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n352), .B1(new_n348), .B2(new_n350), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n357), .A2(new_n359), .A3(new_n360), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n363), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n377), .ZN(new_n393));
  AND3_X1   g192(.A1(new_n380), .A2(new_n381), .A3(KEYINPUT28), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT28), .B1(new_n380), .B2(new_n381), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT71), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n392), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n346), .B1(new_n387), .B2(new_n398), .ZN(new_n399));
  AOI211_X1 g198(.A(KEYINPUT29), .B(new_n345), .C1(new_n392), .C2(new_n396), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n342), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n345), .A2(KEYINPUT29), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n387), .A2(new_n402), .A3(new_n398), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n392), .A2(new_n396), .A3(new_n345), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n403), .A2(new_n404), .A3(new_n322), .ZN(new_n405));
  XOR2_X1   g204(.A(G8gat), .B(G36gat), .Z(new_n406));
  XNOR2_X1  g205(.A(G64gat), .B(G92gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n401), .A2(new_n405), .A3(new_n408), .ZN(new_n409));
  XOR2_X1   g208(.A(new_n408), .B(KEYINPUT72), .Z(new_n410));
  AOI21_X1  g209(.A(new_n410), .B1(new_n401), .B2(new_n405), .ZN(new_n411));
  OAI21_X1  g210(.A(KEYINPUT30), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n401), .A2(new_n405), .A3(new_n408), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT30), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(G120gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(G113gat), .ZN(new_n418));
  INV_X1    g217(.A(G113gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(G120gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT1), .ZN(new_n422));
  XNOR2_X1  g221(.A(G127gat), .B(G134gat), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n421), .B(new_n422), .C1(new_n423), .C2(KEYINPUT65), .ZN(new_n424));
  INV_X1    g223(.A(G127gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(G134gat), .ZN(new_n426));
  INV_X1    g225(.A(G134gat), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(G127gat), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n422), .A2(KEYINPUT65), .ZN(new_n430));
  XNOR2_X1  g229(.A(G113gat), .B(G120gat), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n429), .B(new_n430), .C1(new_n431), .C2(KEYINPUT1), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n424), .A2(new_n432), .ZN(new_n433));
  AOI22_X1  g232(.A1(new_n267), .A2(new_n273), .B1(new_n279), .B2(new_n280), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n287), .A2(new_n288), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n282), .A2(new_n289), .A3(new_n424), .A4(new_n432), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n436), .A2(KEYINPUT75), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT75), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n311), .A2(new_n439), .A3(new_n433), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(G225gat), .A2(G233gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT3), .B1(new_n435), .B2(new_n434), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n444), .A2(new_n290), .A3(new_n433), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT4), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n437), .A2(new_n446), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n424), .A2(new_n432), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n448), .A2(KEYINPUT4), .A3(new_n310), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n445), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n442), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n443), .A2(new_n452), .A3(KEYINPUT39), .ZN(new_n453));
  XNOR2_X1  g252(.A(G57gat), .B(G85gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n454), .B(KEYINPUT78), .ZN(new_n455));
  XOR2_X1   g254(.A(KEYINPUT77), .B(KEYINPUT0), .Z(new_n456));
  XNOR2_X1  g255(.A(new_n455), .B(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(G1gat), .B(G29gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n457), .B(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT39), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n450), .A2(new_n461), .A3(new_n451), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n453), .A2(KEYINPUT40), .A3(new_n460), .A4(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n438), .A2(new_n451), .A3(new_n440), .ZN(new_n464));
  XOR2_X1   g263(.A(KEYINPUT76), .B(KEYINPUT5), .Z(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n445), .A2(new_n447), .A3(new_n442), .A4(new_n449), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OR2_X1    g268(.A1(new_n468), .A2(new_n465), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n469), .A2(new_n459), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n463), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n452), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n459), .B1(new_n473), .B2(new_n461), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT40), .B1(new_n474), .B2(new_n453), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n341), .B1(new_n416), .B2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(KEYINPUT82), .B(KEYINPUT37), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n401), .A2(new_n405), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT83), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n401), .A2(KEYINPUT83), .A3(new_n405), .A4(new_n478), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n410), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT38), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n403), .A2(new_n404), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n487), .A2(new_n319), .A3(new_n321), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n387), .A2(new_n398), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n400), .B1(new_n489), .B2(new_n345), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(new_n308), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n486), .B1(new_n492), .B2(KEYINPUT37), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n483), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n468), .A2(new_n465), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n495), .B1(new_n468), .B2(new_n467), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT6), .B1(new_n496), .B2(new_n459), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n469), .A2(new_n470), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n460), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n469), .A2(KEYINPUT6), .A3(new_n470), .A4(new_n459), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT84), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n496), .A2(KEYINPUT84), .A3(KEYINPUT6), .A4(new_n459), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n494), .A2(new_n500), .A3(new_n413), .A4(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n401), .A2(new_n405), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n408), .B1(new_n507), .B2(KEYINPUT37), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n485), .B1(new_n483), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n477), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT85), .ZN(new_n511));
  INV_X1    g310(.A(new_n340), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(new_n335), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n507), .A2(new_n484), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n414), .B1(new_n514), .B2(new_n413), .ZN(new_n515));
  INV_X1    g314(.A(new_n415), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n500), .A2(new_n501), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n513), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(G227gat), .A2(G233gat), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n433), .B1(new_n372), .B2(new_n386), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n392), .A2(new_n396), .A3(new_n448), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT32), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT66), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G15gat), .B(G43gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(G71gat), .B(G99gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n520), .ZN(new_n529));
  AND3_X1   g328(.A1(new_n392), .A2(new_n448), .A3(new_n396), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n448), .B1(new_n392), .B2(new_n396), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT33), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n528), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT66), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n532), .A2(new_n535), .A3(KEYINPUT32), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n525), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT67), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT67), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n525), .A2(new_n534), .A3(new_n539), .A4(new_n536), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n528), .A2(new_n533), .ZN(new_n542));
  NOR3_X1   g341(.A1(new_n523), .A2(new_n524), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n521), .A2(new_n522), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT34), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n547), .B1(new_n520), .B2(KEYINPUT68), .ZN(new_n548));
  OR3_X1    g347(.A1(new_n546), .A2(new_n529), .A3(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n548), .B1(new_n546), .B2(new_n529), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n545), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n551), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n541), .A2(new_n544), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n552), .A2(KEYINPUT36), .A3(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT36), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n553), .B1(new_n541), .B2(new_n544), .ZN(new_n557));
  AOI211_X1 g356(.A(new_n543), .B(new_n551), .C1(new_n538), .C2(new_n540), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n519), .B1(new_n555), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT85), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n477), .B(new_n561), .C1(new_n506), .C2(new_n509), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n511), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n501), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n564), .B1(new_n497), .B2(new_n499), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n416), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n566), .A2(new_n552), .A3(new_n554), .A4(new_n513), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT35), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n557), .A2(new_n558), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n505), .A2(new_n500), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n416), .A2(KEYINPUT35), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n569), .A2(new_n513), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n260), .B1(new_n563), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(G64gat), .ZN(new_n575));
  AND2_X1   g374(.A1(new_n575), .A2(G57gat), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n575), .A2(G57gat), .ZN(new_n577));
  AND2_X1   g376(.A1(G71gat), .A2(G78gat), .ZN(new_n578));
  OAI22_X1  g377(.A1(new_n576), .A2(new_n577), .B1(KEYINPUT9), .B2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G71gat), .B(G78gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT21), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G127gat), .B(G155gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n213), .B1(new_n583), .B2(new_n582), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT92), .ZN(new_n590));
  XOR2_X1   g389(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G183gat), .B(G211gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n588), .B(new_n594), .ZN(new_n595));
  AND2_X1   g394(.A1(G232gat), .A2(G233gat), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n596), .A2(KEYINPUT41), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT93), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(G134gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(G162gat), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT95), .B(G85gat), .ZN(new_n602));
  INV_X1    g401(.A(G92gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G85gat), .A2(G92gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT7), .ZN(new_n606));
  INV_X1    g405(.A(G99gat), .ZN(new_n607));
  INV_X1    g406(.A(G106gat), .ZN(new_n608));
  OAI21_X1  g407(.A(KEYINPUT8), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n604), .A2(new_n606), .A3(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(G99gat), .B(G106gat), .Z(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n611), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n613), .A2(new_n604), .A3(new_n606), .A4(new_n609), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n612), .A2(KEYINPUT96), .A3(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT96), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n610), .A2(new_n616), .A3(new_n611), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(KEYINPUT97), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT97), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n615), .A2(new_n620), .A3(new_n617), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n243), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  AOI22_X1  g421(.A1(new_n618), .A2(new_n241), .B1(KEYINPUT41), .B2(new_n596), .ZN(new_n623));
  XNOR2_X1  g422(.A(G190gat), .B(G218gat), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT94), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n624), .B1(new_n622), .B2(new_n623), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n601), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n622), .A2(new_n623), .ZN(new_n629));
  INV_X1    g428(.A(new_n624), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n631), .A2(KEYINPUT94), .A3(new_n625), .A4(new_n600), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(G120gat), .B(G148gat), .Z(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT100), .ZN(new_n635));
  XNOR2_X1  g434(.A(G176gat), .B(G204gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(G230gat), .A2(G233gat), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n615), .A2(new_n582), .A3(new_n617), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT10), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n581), .A2(new_n612), .A3(new_n614), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n581), .A2(KEYINPUT10), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n618), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n639), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n638), .B1(new_n640), .B2(new_n642), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n637), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n643), .A2(KEYINPUT98), .A3(new_n645), .ZN(new_n649));
  AOI21_X1  g448(.A(KEYINPUT98), .B1(new_n643), .B2(new_n645), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n649), .A2(new_n650), .A3(new_n639), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT99), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n637), .B1(new_n647), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n653), .B1(new_n652), .B2(new_n647), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n648), .B1(new_n651), .B2(new_n654), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n595), .A2(new_n633), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n574), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n657), .A2(new_n518), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n658), .B(G1gat), .Z(G1324gat));
  INV_X1    g458(.A(KEYINPUT42), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n657), .A2(new_n517), .ZN(new_n661));
  XOR2_X1   g460(.A(KEYINPUT16), .B(G8gat), .Z(new_n662));
  AOI21_X1  g461(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(G8gat), .B1(new_n657), .B2(new_n517), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT101), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n660), .A2(KEYINPUT101), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n666), .B1(new_n662), .B2(new_n667), .ZN(new_n668));
  AOI22_X1  g467(.A1(new_n663), .A2(new_n664), .B1(new_n661), .B2(new_n668), .ZN(G1325gat));
  NAND2_X1  g468(.A1(new_n555), .A2(new_n559), .ZN(new_n670));
  OAI21_X1  g469(.A(G15gat), .B1(new_n657), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n569), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n672), .A2(G15gat), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n671), .B1(new_n657), .B2(new_n673), .ZN(G1326gat));
  NOR2_X1   g473(.A1(new_n657), .A2(new_n513), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT43), .B(G22gat), .Z(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1327gat));
  INV_X1    g476(.A(new_n655), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n595), .A2(new_n633), .A3(new_n678), .ZN(new_n679));
  AOI211_X1 g478(.A(new_n260), .B(new_n679), .C1(new_n563), .C2(new_n573), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n681), .A2(G29gat), .A3(new_n518), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n682), .B(KEYINPUT45), .Z(new_n683));
  INV_X1    g482(.A(new_n633), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n684), .B1(new_n563), .B2(new_n573), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n685), .A2(KEYINPUT44), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687));
  AOI211_X1 g486(.A(new_n687), .B(new_n684), .C1(new_n563), .C2(new_n573), .ZN(new_n688));
  INV_X1    g487(.A(new_n260), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n655), .B(KEYINPUT102), .Z(new_n690));
  NAND3_X1  g489(.A1(new_n689), .A2(new_n690), .A3(new_n595), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n686), .A2(new_n688), .A3(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(G29gat), .B1(new_n693), .B2(new_n518), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n683), .A2(new_n694), .ZN(G1328gat));
  NOR3_X1   g494(.A1(new_n681), .A2(G36gat), .A3(new_n517), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT46), .ZN(new_n697));
  OAI21_X1  g496(.A(G36gat), .B1(new_n693), .B2(new_n517), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(G1329gat));
  INV_X1    g498(.A(new_n670), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n692), .A2(G43gat), .A3(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n681), .A2(new_n672), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n701), .B1(G43gat), .B2(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g503(.A(KEYINPUT48), .ZN(new_n705));
  INV_X1    g504(.A(G50gat), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n706), .B1(new_n692), .B2(new_n341), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n513), .A2(G50gat), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n680), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n705), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n563), .A2(new_n573), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n633), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(new_n687), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n685), .A2(KEYINPUT44), .ZN(new_n714));
  INV_X1    g513(.A(new_n691), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n713), .A2(new_n341), .A3(new_n714), .A4(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(G50gat), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT104), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT103), .ZN(new_n719));
  INV_X1    g518(.A(new_n679), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n574), .A2(new_n719), .A3(new_n720), .A4(new_n708), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(KEYINPUT48), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n719), .B1(new_n680), .B2(new_n708), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n717), .A2(new_n718), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n718), .B1(new_n717), .B2(new_n724), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n710), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT105), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n710), .B(KEYINPUT105), .C1(new_n725), .C2(new_n726), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(G1331gat));
  NOR4_X1   g530(.A1(new_n689), .A2(new_n690), .A3(new_n595), .A4(new_n633), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n711), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n565), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(G57gat), .ZN(G1332gat));
  AND2_X1   g534(.A1(new_n733), .A2(new_n416), .ZN(new_n736));
  NOR2_X1   g535(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n737));
  AND2_X1   g536(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n739), .B1(new_n736), .B2(new_n737), .ZN(G1333gat));
  NAND2_X1  g539(.A1(new_n733), .A2(new_n700), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n672), .A2(G71gat), .ZN(new_n742));
  AOI22_X1  g541(.A1(new_n741), .A2(G71gat), .B1(new_n733), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(KEYINPUT106), .B(KEYINPUT50), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(G1334gat));
  NAND2_X1  g544(.A1(new_n733), .A2(new_n341), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(G78gat), .ZN(G1335gat));
  INV_X1    g546(.A(new_n595), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n689), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n685), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n753), .A2(KEYINPUT107), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT107), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n750), .A2(new_n755), .A3(new_n751), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n752), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n757), .A2(new_n565), .A3(new_n602), .A4(new_n655), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n686), .A2(new_n688), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n689), .A2(new_n678), .A3(new_n748), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n761), .A2(new_n518), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n758), .B1(new_n602), .B2(new_n762), .ZN(G1336gat));
  NAND3_X1  g562(.A1(new_n759), .A2(new_n416), .A3(new_n760), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT52), .B1(new_n764), .B2(G92gat), .ZN(new_n765));
  INV_X1    g564(.A(new_n757), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n690), .A2(G92gat), .A3(new_n517), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n765), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  OR2_X1    g568(.A1(new_n752), .A2(KEYINPUT108), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n752), .A2(KEYINPUT108), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n770), .B(new_n771), .C1(new_n754), .C2(new_n756), .ZN(new_n772));
  AOI22_X1  g571(.A1(new_n772), .A2(new_n767), .B1(G92gat), .B2(new_n764), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n769), .B1(new_n773), .B2(new_n774), .ZN(G1337gat));
  NAND4_X1  g574(.A1(new_n757), .A2(new_n607), .A3(new_n569), .A4(new_n655), .ZN(new_n776));
  OAI21_X1  g575(.A(G99gat), .B1(new_n761), .B2(new_n670), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(G1338gat));
  NAND3_X1  g577(.A1(new_n759), .A2(new_n341), .A3(new_n760), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT53), .B1(new_n779), .B2(G106gat), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n690), .A2(G106gat), .A3(new_n513), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n780), .B1(new_n766), .B2(new_n782), .ZN(new_n783));
  AOI22_X1  g582(.A1(new_n772), .A2(new_n781), .B1(G106gat), .B2(new_n779), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n783), .B1(new_n784), .B2(new_n785), .ZN(G1339gat));
  NAND2_X1  g585(.A1(new_n656), .A2(new_n260), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n258), .A2(new_n207), .A3(new_n251), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n253), .A2(new_n254), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n244), .A2(new_n233), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n205), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n651), .A2(new_n654), .ZN(new_n795));
  XOR2_X1   g594(.A(KEYINPUT110), .B(KEYINPUT54), .Z(new_n796));
  NAND2_X1  g595(.A1(new_n646), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n637), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n638), .B1(new_n618), .B2(new_n644), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n643), .A2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT109), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n643), .A2(new_n799), .A3(KEYINPUT109), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n802), .A2(KEYINPUT54), .A3(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n650), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n643), .A2(KEYINPUT98), .A3(new_n645), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n805), .A2(new_n638), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n798), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n795), .B1(new_n808), .B2(KEYINPUT55), .ZN(new_n809));
  INV_X1    g608(.A(new_n637), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n810), .B1(new_n646), .B2(new_n796), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n802), .A2(KEYINPUT54), .A3(new_n803), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n811), .B1(new_n651), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814));
  AOI22_X1  g613(.A1(new_n813), .A2(new_n814), .B1(new_n628), .B2(new_n632), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n794), .A2(new_n809), .A3(new_n815), .ZN(new_n816));
  AND3_X1   g615(.A1(new_n789), .A2(new_n655), .A3(new_n792), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n247), .A2(new_n251), .A3(new_n256), .ZN(new_n818));
  INV_X1    g617(.A(new_n207), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AOI22_X1  g619(.A1(new_n820), .A2(new_n789), .B1(new_n814), .B2(new_n813), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n817), .B1(new_n821), .B2(new_n809), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n816), .B1(new_n822), .B2(new_n633), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n788), .B1(new_n823), .B2(new_n595), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n824), .A2(new_n672), .A3(new_n341), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n518), .A2(new_n416), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(G113gat), .B1(new_n827), .B2(new_n260), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n689), .A2(new_n419), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(KEYINPUT111), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n828), .B1(new_n827), .B2(new_n830), .ZN(G1340gat));
  NOR3_X1   g630(.A1(new_n827), .A2(new_n417), .A3(new_n690), .ZN(new_n832));
  INV_X1    g631(.A(new_n827), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n655), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n832), .B1(new_n417), .B2(new_n834), .ZN(G1341gat));
  NOR2_X1   g634(.A1(new_n827), .A2(new_n595), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(new_n425), .ZN(G1342gat));
  NAND3_X1  g636(.A1(new_n825), .A2(new_n633), .A3(new_n826), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(G134gat), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT112), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n839), .B(new_n840), .ZN(new_n841));
  OR3_X1    g640(.A1(new_n838), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT56), .B1(new_n838), .B2(G134gat), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT113), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n839), .B(KEYINPUT112), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT113), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n846), .A2(new_n847), .A3(new_n843), .A4(new_n842), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n845), .A2(new_n848), .ZN(G1343gat));
  NAND2_X1  g648(.A1(new_n670), .A2(new_n826), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT57), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n851), .B1(new_n824), .B2(new_n513), .ZN(new_n852));
  INV_X1    g651(.A(new_n815), .ZN(new_n853));
  OAI22_X1  g652(.A1(new_n813), .A2(new_n814), .B1(new_n651), .B2(new_n654), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n853), .A2(new_n793), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n813), .A2(new_n814), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n856), .B1(new_n257), .B2(new_n259), .ZN(new_n857));
  OAI22_X1  g656(.A1(new_n857), .A2(new_n854), .B1(new_n678), .B2(new_n793), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n855), .B1(new_n858), .B2(new_n684), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n787), .B1(new_n859), .B2(new_n748), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(KEYINPUT57), .A3(new_n341), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n850), .B1(new_n852), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n275), .B1(new_n862), .B2(new_n689), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT58), .B1(new_n863), .B2(KEYINPUT114), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT115), .ZN(new_n865));
  INV_X1    g664(.A(new_n850), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n824), .A2(new_n851), .A3(new_n513), .ZN(new_n867));
  AOI21_X1  g666(.A(KEYINPUT57), .B1(new_n860), .B2(new_n341), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n689), .B(new_n866), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(G141gat), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n860), .A2(new_n341), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n689), .A2(new_n275), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n871), .A2(new_n850), .A3(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n865), .B1(new_n870), .B2(new_n874), .ZN(new_n875));
  AOI211_X1 g674(.A(KEYINPUT115), .B(new_n873), .C1(new_n869), .C2(G141gat), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n864), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(KEYINPUT115), .B1(new_n863), .B2(new_n873), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n870), .A2(new_n874), .A3(new_n865), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT114), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n870), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n878), .A2(new_n879), .A3(KEYINPUT58), .A4(new_n881), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n877), .A2(new_n882), .ZN(G1344gat));
  NOR2_X1   g682(.A1(new_n850), .A2(new_n678), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n860), .A2(new_n277), .A3(new_n341), .A4(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n886));
  INV_X1    g685(.A(new_n884), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n809), .A2(new_n815), .A3(KEYINPUT116), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n794), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT116), .B1(new_n809), .B2(new_n815), .ZN(new_n890));
  OAI22_X1  g689(.A1(new_n822), .A2(new_n633), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT117), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n748), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI221_X1 g692(.A(KEYINPUT117), .B1(new_n889), .B2(new_n890), .C1(new_n822), .C2(new_n633), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n788), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n851), .B1(new_n895), .B2(new_n513), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n887), .B1(new_n896), .B2(new_n861), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT118), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n277), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n891), .A2(new_n892), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n894), .A3(new_n595), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n513), .B1(new_n901), .B2(new_n787), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n861), .B1(new_n902), .B2(KEYINPUT57), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n884), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(KEYINPUT118), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n886), .B1(new_n899), .B2(new_n905), .ZN(new_n906));
  AOI211_X1 g705(.A(KEYINPUT59), .B(new_n277), .C1(new_n862), .C2(new_n655), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n885), .B1(new_n906), .B2(new_n907), .ZN(G1345gat));
  NOR2_X1   g707(.A1(new_n871), .A2(new_n850), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n748), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(KEYINPUT119), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n911), .A2(G155gat), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(KEYINPUT119), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n595), .A2(new_n268), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT120), .ZN(new_n915));
  AOI22_X1  g714(.A1(new_n912), .A2(new_n913), .B1(new_n862), .B2(new_n915), .ZN(G1346gat));
  NAND2_X1  g715(.A1(new_n862), .A2(new_n633), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n684), .A2(G162gat), .ZN(new_n918));
  AOI22_X1  g717(.A1(new_n917), .A2(G162gat), .B1(new_n909), .B2(new_n918), .ZN(new_n919));
  XOR2_X1   g718(.A(new_n919), .B(KEYINPUT121), .Z(G1347gat));
  NOR2_X1   g719(.A1(new_n517), .A2(new_n565), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n825), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(G169gat), .B1(new_n922), .B2(new_n689), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n921), .B(KEYINPUT122), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n825), .A2(new_n924), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n925), .A2(new_n355), .A3(new_n260), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n923), .A2(new_n926), .ZN(G1348gat));
  NAND3_X1  g726(.A1(new_n922), .A2(new_n356), .A3(new_n655), .ZN(new_n928));
  OAI21_X1  g727(.A(G176gat), .B1(new_n925), .B2(new_n690), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(G1349gat));
  NAND3_X1  g729(.A1(new_n825), .A2(new_n748), .A3(new_n924), .ZN(new_n931));
  OR2_X1    g730(.A1(new_n931), .A2(KEYINPUT123), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n367), .B1(new_n931), .B2(KEYINPUT123), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n748), .A2(new_n381), .ZN(new_n934));
  AOI22_X1  g733(.A1(new_n932), .A2(new_n933), .B1(new_n922), .B2(new_n934), .ZN(new_n935));
  XOR2_X1   g734(.A(KEYINPUT124), .B(KEYINPUT60), .Z(new_n936));
  XNOR2_X1  g735(.A(new_n935), .B(new_n936), .ZN(G1350gat));
  NAND3_X1  g736(.A1(new_n922), .A2(new_n380), .A3(new_n633), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n825), .A2(new_n633), .A3(new_n924), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT61), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n939), .A2(new_n940), .A3(G190gat), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n940), .B1(new_n939), .B2(G190gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n938), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT125), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n943), .B(new_n944), .ZN(G1351gat));
  AND2_X1   g744(.A1(new_n924), .A2(new_n670), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n903), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(G197gat), .B1(new_n947), .B2(new_n260), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n670), .A2(new_n341), .A3(new_n921), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n860), .A2(new_n949), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n950), .A2(G197gat), .A3(new_n260), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT126), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n948), .A2(new_n952), .ZN(G1352gat));
  NOR3_X1   g752(.A1(new_n950), .A2(G204gat), .A3(new_n678), .ZN(new_n954));
  XOR2_X1   g753(.A(new_n954), .B(KEYINPUT127), .Z(new_n955));
  INV_X1    g754(.A(KEYINPUT62), .ZN(new_n956));
  OR2_X1    g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n955), .A2(new_n956), .ZN(new_n958));
  OAI21_X1  g757(.A(G204gat), .B1(new_n947), .B2(new_n690), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(G1353gat));
  OR3_X1    g759(.A1(new_n950), .A2(G211gat), .A3(new_n595), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n903), .A2(new_n748), .A3(new_n946), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n962), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n963));
  AOI21_X1  g762(.A(KEYINPUT63), .B1(new_n962), .B2(G211gat), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(G1354gat));
  OAI21_X1  g764(.A(G218gat), .B1(new_n947), .B2(new_n684), .ZN(new_n966));
  OR3_X1    g765(.A1(new_n950), .A2(G218gat), .A3(new_n684), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(G1355gat));
endmodule


