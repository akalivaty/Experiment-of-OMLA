//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 1 0 1 1 0 1 0 1 1 0 0 1 1 1 0 0 0 0 0 1 1 0 0 0 1 1 1 0 0 1 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1219,
    new_n1220, new_n1221, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1282, new_n1283, new_n1284, new_n1285;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  OAI21_X1  g0006(.A(G50), .B1(G58), .B2(G68), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT64), .ZN(new_n208));
  AND2_X1   g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  NAND3_X1  g0009(.A1(new_n208), .A2(G20), .A3(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G13), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT0), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n210), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n220));
  INV_X1    g0020(.A(G116), .ZN(new_n221));
  INV_X1    g0021(.A(G270), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G97), .A2(G257), .ZN(new_n225));
  INV_X1    g0025(.A(G68), .ZN(new_n226));
  INV_X1    g0026(.A(G238), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n224), .B(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  AOI211_X1 g0028(.A(new_n223), .B(new_n228), .C1(G58), .C2(G232), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n213), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT1), .Z(new_n231));
  AOI211_X1 g0031(.A(new_n219), .B(new_n231), .C1(new_n218), .C2(new_n217), .ZN(G361));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT2), .ZN(new_n235));
  INV_X1    g0035(.A(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G264), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(new_n222), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT65), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G107), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(new_n221), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G351));
  NAND2_X1  g0049(.A1(G33), .A2(G97), .ZN(new_n250));
  OR2_X1    g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G1698), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n253), .B1(G232), .B2(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G226), .A2(G1698), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n250), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  AND2_X1   g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G1), .A2(G13), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G41), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n209), .B(KEYINPUT67), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT67), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n265), .B1(new_n258), .B2(new_n259), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G45), .ZN(new_n268));
  AOI21_X1  g0068(.A(G1), .B1(new_n263), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT66), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G274), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n273), .B1(new_n269), .B2(KEYINPUT66), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n267), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n267), .A2(G238), .A3(new_n270), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT71), .ZN(new_n277));
  AND3_X1   g0077(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n277), .B1(new_n275), .B2(new_n276), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n261), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT13), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT72), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT13), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n283), .B(new_n261), .C1(new_n278), .C2(new_n279), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n281), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n280), .A2(KEYINPUT72), .A3(KEYINPUT13), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(G169), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT14), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n281), .A2(G179), .A3(new_n284), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT14), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n285), .A2(new_n290), .A3(G169), .A4(new_n286), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n288), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n211), .A2(G13), .A3(G20), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(G68), .ZN(new_n294));
  OR2_X1    g0094(.A1(new_n294), .A2(KEYINPUT73), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT12), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n296), .B1(new_n294), .B2(KEYINPUT73), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(new_n297), .ZN(new_n299));
  NAND3_X1  g0099(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n259), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n211), .A2(G20), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n298), .B(new_n299), .C1(new_n226), .C2(new_n304), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n305), .B(KEYINPUT74), .ZN(new_n306));
  NOR2_X1   g0106(.A1(G20), .A2(G33), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G50), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n212), .A2(G33), .ZN(new_n310));
  OAI22_X1  g0110(.A1(new_n308), .A2(new_n309), .B1(new_n310), .B2(new_n202), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n212), .A2(G68), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n301), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n313), .B(KEYINPUT11), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n306), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n292), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g0116(.A(KEYINPUT8), .B(G58), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n318), .A2(new_n307), .B1(G20), .B2(G77), .ZN(new_n319));
  XNOR2_X1  g0119(.A(KEYINPUT15), .B(G87), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n319), .B1(new_n310), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n293), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n321), .A2(new_n301), .B1(new_n202), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n302), .A2(G77), .A3(new_n303), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n275), .ZN(new_n326));
  AND2_X1   g0126(.A1(KEYINPUT3), .A2(G33), .ZN(new_n327));
  NOR2_X1   g0127(.A1(KEYINPUT3), .A2(G33), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n329), .A2(G1698), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G232), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n329), .A2(G107), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n253), .A2(G1698), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n333), .B(KEYINPUT69), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n331), .B(new_n332), .C1(new_n334), .C2(new_n227), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n326), .B1(new_n335), .B2(new_n260), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n269), .B1(new_n264), .B2(new_n266), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G244), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n325), .B1(new_n339), .B2(G179), .ZN(new_n340));
  AOI21_X1  g0140(.A(G169), .B1(new_n336), .B2(new_n338), .ZN(new_n341));
  OR2_X1    g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AND2_X1   g0142(.A1(new_n316), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n315), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n285), .A2(G200), .A3(new_n286), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n281), .A2(G190), .A3(new_n284), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n293), .A2(G50), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n304), .A2(new_n309), .ZN(new_n350));
  INV_X1    g0150(.A(G150), .ZN(new_n351));
  OAI22_X1  g0151(.A1(new_n317), .A2(new_n310), .B1(new_n351), .B2(new_n308), .ZN(new_n352));
  XNOR2_X1  g0152(.A(new_n352), .B(KEYINPUT70), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(new_n212), .B2(new_n201), .ZN(new_n354));
  AOI211_X1 g0154(.A(new_n349), .B(new_n350), .C1(new_n354), .C2(new_n301), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n330), .A2(G222), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT68), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n357), .B(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n329), .A2(G77), .ZN(new_n360));
  INV_X1    g0160(.A(G223), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n359), .B(new_n360), .C1(new_n361), .C2(new_n334), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n260), .ZN(new_n363));
  INV_X1    g0163(.A(new_n337), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n364), .A2(new_n236), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n363), .A2(new_n275), .A3(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n356), .B1(new_n367), .B2(G179), .ZN(new_n368));
  AOI211_X1 g0168(.A(new_n326), .B(new_n365), .C1(new_n362), .C2(new_n260), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n369), .A2(G169), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n363), .A2(G190), .A3(new_n275), .A4(new_n366), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n355), .A2(KEYINPUT9), .ZN(new_n373));
  INV_X1    g0173(.A(G200), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n372), .B(new_n373), .C1(new_n369), .C2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n355), .A2(KEYINPUT9), .ZN(new_n376));
  OAI21_X1  g0176(.A(KEYINPUT10), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n367), .A2(G200), .B1(KEYINPUT9), .B2(new_n355), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT10), .ZN(new_n379));
  INV_X1    g0179(.A(new_n376), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n378), .A2(new_n379), .A3(new_n380), .A4(new_n372), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n371), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n325), .B1(new_n339), .B2(G200), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n336), .A2(G190), .A3(new_n338), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI211_X1 g0185(.A(G223), .B(new_n254), .C1(new_n327), .C2(new_n328), .ZN(new_n386));
  OAI211_X1 g0186(.A(G226), .B(G1698), .C1(new_n327), .C2(new_n328), .ZN(new_n387));
  NAND2_X1  g0187(.A1(G33), .A2(G87), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT78), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n386), .A2(new_n387), .A3(KEYINPUT78), .A4(new_n388), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n391), .A2(new_n260), .A3(new_n392), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n266), .A2(new_n264), .B1(new_n270), .B2(new_n271), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n394), .A2(new_n274), .B1(new_n337), .B2(G232), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(G169), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n393), .A2(G179), .A3(new_n395), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AND2_X1   g0199(.A1(G58), .A2(G68), .ZN(new_n400));
  NOR2_X1   g0200(.A1(G58), .A2(G68), .ZN(new_n401));
  OAI21_X1  g0201(.A(G20), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(KEYINPUT75), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n307), .A2(G159), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT75), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n405), .B(G20), .C1(new_n400), .C2(new_n401), .ZN(new_n406));
  AND3_X1   g0206(.A1(new_n403), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(KEYINPUT7), .B1(new_n329), .B2(new_n212), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT7), .ZN(new_n409));
  NOR4_X1   g0209(.A1(new_n327), .A2(new_n328), .A3(new_n409), .A4(G20), .ZN(new_n410));
  OAI21_X1  g0210(.A(G68), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT76), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n407), .B(new_n411), .C1(new_n412), .C2(KEYINPUT16), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT16), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n403), .A2(new_n412), .A3(new_n404), .A4(new_n406), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n251), .A2(new_n212), .A3(new_n252), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n409), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n251), .A2(KEYINPUT7), .A3(new_n212), .A4(new_n252), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n226), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n403), .A2(new_n404), .A3(new_n406), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n414), .B(new_n415), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n413), .A2(new_n421), .A3(new_n301), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n318), .A2(new_n303), .ZN(new_n423));
  XNOR2_X1  g0223(.A(new_n423), .B(KEYINPUT77), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n322), .A2(new_n301), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n424), .A2(new_n425), .B1(new_n322), .B2(new_n317), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n399), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT18), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n397), .A2(new_n398), .B1(new_n422), .B2(new_n426), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT18), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n393), .A2(G190), .A3(new_n395), .ZN(new_n433));
  AND3_X1   g0233(.A1(new_n422), .A2(new_n426), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT17), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n396), .A2(G200), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n436), .A2(new_n422), .A3(new_n426), .A4(new_n433), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT17), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n430), .A2(new_n432), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n382), .A2(new_n385), .A3(new_n440), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n348), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n322), .A2(new_n221), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n211), .A2(G33), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n293), .A2(new_n444), .A3(new_n259), .A4(new_n300), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n443), .B1(new_n445), .B2(new_n221), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n221), .A2(G20), .ZN(new_n447));
  AOI21_X1  g0247(.A(G20), .B1(G33), .B2(G283), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n262), .A2(G97), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT83), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n450), .B1(new_n448), .B2(new_n449), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n301), .B(new_n447), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT20), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n448), .A2(new_n449), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT83), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n302), .B1(new_n458), .B2(new_n451), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n459), .A2(KEYINPUT20), .A3(new_n447), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n446), .B1(new_n456), .B2(new_n460), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n251), .A2(new_n252), .B1(G257), .B2(new_n254), .ZN(new_n462));
  NAND2_X1  g0262(.A1(G264), .A2(G1698), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G303), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n329), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n464), .A2(new_n260), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT80), .ZN(new_n468));
  XOR2_X1   g0268(.A(KEYINPUT5), .B(G41), .Z(new_n469));
  NAND4_X1  g0269(.A1(new_n265), .A2(new_n211), .A3(G45), .A4(G274), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n470), .ZN(new_n472));
  XNOR2_X1  g0272(.A(KEYINPUT5), .B(G41), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n472), .A2(KEYINPUT80), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n473), .A2(new_n211), .A3(G45), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n267), .A2(G270), .A3(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n467), .A2(new_n475), .A3(G179), .A4(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n461), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n456), .A2(new_n460), .ZN(new_n480));
  INV_X1    g0280(.A(new_n446), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(G169), .ZN(new_n483));
  INV_X1    g0283(.A(new_n260), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n484), .B1(new_n462), .B2(new_n463), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n485), .A2(new_n466), .B1(new_n471), .B2(new_n474), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n483), .B1(new_n486), .B2(new_n477), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n482), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT21), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n479), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n253), .A2(G257), .A3(G1698), .ZN(new_n491));
  NAND2_X1  g0291(.A1(G33), .A2(G294), .ZN(new_n492));
  OAI211_X1 g0292(.A(G250), .B(new_n254), .C1(new_n327), .C2(new_n328), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n260), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n267), .A2(G264), .A3(new_n476), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n495), .A2(new_n475), .A3(new_n496), .ZN(new_n497));
  OR2_X1    g0297(.A1(new_n497), .A2(G179), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n483), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n212), .B(G87), .C1(new_n327), .C2(new_n328), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT22), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT22), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n253), .A2(new_n502), .A3(new_n212), .A4(G87), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n212), .A2(G33), .A3(G116), .ZN(new_n505));
  XNOR2_X1  g0305(.A(new_n505), .B(KEYINPUT85), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n212), .A2(G107), .ZN(new_n508));
  XNOR2_X1  g0308(.A(new_n508), .B(KEYINPUT23), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n504), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(KEYINPUT24), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT24), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n504), .A2(new_n512), .A3(new_n507), .A4(new_n509), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n302), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT79), .ZN(new_n515));
  XNOR2_X1  g0315(.A(new_n445), .B(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(G107), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n293), .A2(G107), .ZN(new_n518));
  XNOR2_X1  g0318(.A(new_n518), .B(KEYINPUT25), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n498), .B(new_n499), .C1(new_n514), .C2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT84), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n467), .A2(new_n475), .A3(new_n477), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(G169), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n461), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n522), .B1(new_n525), .B2(KEYINPUT21), .ZN(new_n526));
  NOR4_X1   g0326(.A1(new_n461), .A2(new_n524), .A3(KEYINPUT84), .A4(new_n489), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n490), .B(new_n521), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n253), .A2(new_n212), .A3(G68), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT19), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n212), .B1(new_n250), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(G87), .B2(new_n205), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n531), .B1(new_n250), .B2(G20), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n530), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n535), .A2(new_n301), .B1(new_n322), .B2(new_n320), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n445), .A2(new_n515), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n445), .A2(new_n515), .ZN(new_n539));
  OAI21_X1  g0339(.A(G87), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT82), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n516), .A2(KEYINPUT82), .A3(G87), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n537), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(G244), .B(G1698), .C1(new_n327), .C2(new_n328), .ZN(new_n545));
  OAI211_X1 g0345(.A(G238), .B(new_n254), .C1(new_n327), .C2(new_n328), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n545), .B(new_n546), .C1(new_n262), .C2(new_n221), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n260), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n267), .B(G250), .C1(G1), .C2(new_n268), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n548), .A2(new_n549), .A3(new_n470), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n374), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n472), .B1(new_n547), .B2(new_n260), .ZN(new_n552));
  INV_X1    g0352(.A(G190), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n552), .A2(new_n553), .A3(new_n549), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  XOR2_X1   g0355(.A(new_n320), .B(KEYINPUT81), .Z(new_n556));
  NAND2_X1  g0356(.A1(new_n516), .A2(new_n556), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n483), .A2(new_n550), .B1(new_n557), .B2(new_n536), .ZN(new_n558));
  INV_X1    g0358(.A(G179), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n552), .A2(new_n559), .A3(new_n549), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n544), .A2(new_n555), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n511), .A2(new_n513), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n301), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n497), .A2(new_n374), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n495), .A2(new_n553), .A3(new_n475), .A4(new_n496), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n520), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n563), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n254), .A2(KEYINPUT4), .A3(G244), .ZN(new_n569));
  INV_X1    g0369(.A(G250), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n569), .B1(new_n570), .B2(new_n254), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n571), .A2(new_n253), .B1(G33), .B2(G283), .ZN(new_n572));
  OAI211_X1 g0372(.A(G244), .B(new_n254), .C1(new_n327), .C2(new_n328), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT4), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n484), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n267), .A2(G257), .A3(new_n476), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n577), .A2(new_n553), .A3(new_n475), .A4(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n475), .ZN(new_n580));
  INV_X1    g0380(.A(new_n578), .ZN(new_n581));
  NOR3_X1   g0381(.A1(new_n580), .A2(new_n576), .A3(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n579), .B1(new_n582), .B2(G200), .ZN(new_n583));
  OAI21_X1  g0383(.A(G107), .B1(new_n408), .B2(new_n410), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT6), .ZN(new_n585));
  INV_X1    g0385(.A(G97), .ZN(new_n586));
  INV_X1    g0386(.A(G107), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n585), .B1(new_n588), .B2(new_n204), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n587), .A2(KEYINPUT6), .A3(G97), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(G20), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n307), .A2(G77), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n584), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n301), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n293), .A2(G97), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n516), .A2(G97), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n595), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n583), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n582), .A2(new_n559), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n577), .A2(new_n475), .A3(new_n578), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n483), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n595), .A2(new_n597), .A3(new_n598), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n601), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n561), .A2(new_n568), .A3(new_n600), .A4(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n523), .A2(new_n553), .ZN(new_n607));
  AOI211_X1 g0407(.A(new_n607), .B(new_n482), .C1(G200), .C2(new_n523), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n442), .A2(new_n529), .A3(new_n609), .ZN(G372));
  NAND2_X1  g0410(.A1(new_n550), .A2(new_n483), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n557), .A2(new_n536), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n611), .A2(new_n612), .A3(new_n560), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n529), .B2(new_n606), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n601), .A2(new_n603), .A3(new_n604), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n616), .A2(new_n561), .A3(KEYINPUT26), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(KEYINPUT86), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT86), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n616), .A2(new_n561), .A3(new_n619), .A4(KEYINPUT26), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT26), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n552), .A2(new_n553), .A3(new_n549), .ZN(new_n622));
  AOI21_X1  g0422(.A(G200), .B1(new_n552), .B2(new_n549), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n540), .A2(new_n541), .ZN(new_n625));
  AOI21_X1  g0425(.A(KEYINPUT82), .B1(new_n516), .B2(G87), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n536), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n613), .B1(new_n624), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n621), .B1(new_n628), .B2(new_n605), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n618), .A2(new_n620), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n615), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n442), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n371), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n377), .A2(new_n381), .ZN(new_n634));
  INV_X1    g0434(.A(new_n347), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n437), .A2(new_n439), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NOR3_X1   g0437(.A1(new_n343), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n430), .A2(new_n432), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n634), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n632), .A2(new_n633), .A3(new_n641), .ZN(G369));
  OR2_X1    g0442(.A1(new_n526), .A2(new_n527), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n490), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n214), .A2(G20), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n211), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(G213), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(G343), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n461), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n644), .A2(new_n653), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n643), .B(new_n490), .C1(new_n461), .C2(new_n652), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n608), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(G330), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n651), .B1(new_n514), .B2(new_n520), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n568), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(new_n521), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n521), .A2(new_n651), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n657), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT87), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n644), .A2(new_n660), .A3(new_n521), .A4(new_n652), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n661), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT88), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n666), .A2(KEYINPUT88), .A3(new_n661), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n665), .B1(new_n670), .B2(new_n672), .ZN(G399));
  OR3_X1    g0473(.A1(new_n215), .A2(KEYINPUT89), .A3(G41), .ZN(new_n674));
  OAI21_X1  g0474(.A(KEYINPUT89), .B1(new_n215), .B2(G41), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n205), .A2(G87), .A3(G116), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G1), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n208), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n678), .B1(new_n679), .B2(new_n676), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT28), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT29), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n631), .A2(new_n682), .A3(new_n652), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n617), .A2(new_n629), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n684), .B(new_n613), .C1(new_n529), .C2(new_n606), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n682), .B1(new_n685), .B2(new_n652), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(G330), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n602), .A2(new_n478), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n495), .A2(new_n496), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(new_n550), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT30), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n691), .A2(KEYINPUT30), .A3(new_n693), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n582), .A2(G179), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n698), .A2(new_n523), .A3(new_n497), .A4(new_n550), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n696), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n651), .ZN(new_n701));
  NOR4_X1   g0501(.A1(new_n528), .A2(new_n606), .A3(new_n608), .A4(new_n651), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT31), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n696), .A2(new_n699), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT90), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n696), .A2(KEYINPUT90), .A3(new_n699), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(new_n697), .A3(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n709), .A2(KEYINPUT31), .A3(new_n651), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n690), .B1(new_n704), .B2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n689), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n681), .B1(new_n714), .B2(G1), .ZN(G364));
  NOR2_X1   g0515(.A1(new_n656), .A2(G330), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT91), .ZN(new_n717));
  INV_X1    g0517(.A(new_n676), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n211), .B1(new_n645), .B2(G45), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n717), .A2(new_n657), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n245), .A2(G45), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n215), .A2(new_n253), .ZN(new_n725));
  OAI211_X1 g0525(.A(new_n724), .B(new_n725), .C1(G45), .C2(new_n679), .ZN(new_n726));
  INV_X1    g0526(.A(G355), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n216), .A2(new_n253), .ZN(new_n728));
  OAI221_X1 g0528(.A(new_n726), .B1(G116), .B2(new_n216), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n259), .B1(G20), .B2(new_n483), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT93), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(G13), .A2(G33), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n733), .B(KEYINPUT92), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(G20), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(G179), .A2(G200), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n212), .B1(new_n737), .B2(G190), .ZN(new_n738));
  INV_X1    g0538(.A(G294), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n559), .A2(G200), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n212), .A2(G190), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(G311), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n212), .A2(new_n553), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n374), .A2(G179), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI221_X1 g0547(.A(new_n329), .B1(new_n743), .B2(new_n744), .C1(new_n465), .C2(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n553), .ZN(new_n750));
  AOI211_X1 g0550(.A(new_n740), .B(new_n748), .C1(G326), .C2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n745), .A2(new_n741), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G322), .ZN(new_n754));
  OR2_X1    g0554(.A1(new_n742), .A2(KEYINPUT94), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n742), .A2(KEYINPUT94), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n755), .A2(new_n746), .A3(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G283), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n749), .A2(G190), .ZN(new_n760));
  AND2_X1   g0560(.A1(new_n760), .A2(KEYINPUT95), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(KEYINPUT95), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  XNOR2_X1  g0564(.A(KEYINPUT33), .B(G317), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n755), .A2(new_n756), .A3(new_n737), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n764), .A2(new_n765), .B1(new_n767), .B2(G329), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n751), .A2(new_n754), .A3(new_n759), .A4(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(G159), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT32), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n757), .A2(new_n587), .ZN(new_n773));
  INV_X1    g0573(.A(G87), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n253), .B1(new_n743), .B2(new_n202), .C1(new_n774), .C2(new_n747), .ZN(new_n775));
  INV_X1    g0575(.A(new_n750), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n776), .A2(new_n309), .B1(new_n738), .B2(new_n586), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n773), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n772), .B(new_n778), .C1(new_n226), .C2(new_n763), .ZN(new_n779));
  INV_X1    g0579(.A(G58), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n752), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n769), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n729), .A2(new_n736), .B1(new_n732), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n735), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n721), .B(new_n783), .C1(new_n656), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n723), .A2(new_n785), .ZN(G396));
  NAND2_X1  g0586(.A1(new_n631), .A2(new_n652), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n340), .A2(new_n341), .A3(new_n651), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n325), .A2(new_n651), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n385), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n788), .B1(new_n790), .B2(new_n342), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n787), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n630), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n791), .B(new_n652), .C1(new_n794), .C2(new_n614), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(new_n711), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(new_n722), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n757), .A2(new_n226), .ZN(new_n799));
  INV_X1    g0599(.A(G132), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n253), .B1(new_n780), .B2(new_n738), .C1(new_n766), .C2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n743), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n802), .A2(G159), .B1(G137), .B2(new_n750), .ZN(new_n803));
  INV_X1    g0603(.A(G143), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n803), .B1(new_n804), .B2(new_n752), .C1(new_n763), .C2(new_n351), .ZN(new_n805));
  XNOR2_X1  g0605(.A(KEYINPUT98), .B(KEYINPUT34), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n799), .B(new_n801), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n807), .B1(new_n309), .B2(new_n747), .C1(new_n806), .C2(new_n805), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n776), .A2(new_n465), .B1(new_n738), .B2(new_n586), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n766), .A2(new_n744), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n757), .A2(new_n774), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n329), .B1(new_n752), .B2(new_n739), .C1(new_n587), .C2(new_n747), .ZN(new_n812));
  NOR4_X1   g0612(.A1(new_n809), .A2(new_n810), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  OR2_X1    g0613(.A1(new_n764), .A2(KEYINPUT97), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n764), .A2(KEYINPUT97), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(G283), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n813), .B1(new_n221), .B2(new_n743), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n731), .B1(new_n808), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n731), .A2(new_n734), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(KEYINPUT96), .Z(new_n821));
  AOI21_X1  g0621(.A(new_n819), .B1(new_n202), .B2(new_n821), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n721), .B(new_n822), .C1(new_n791), .C2(new_n734), .ZN(new_n823));
  XOR2_X1   g0623(.A(new_n823), .B(KEYINPUT99), .Z(new_n824));
  NAND2_X1  g0624(.A1(new_n798), .A2(new_n824), .ZN(G384));
  NOR2_X1   g0625(.A1(new_n701), .A2(new_n703), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n792), .B1(new_n704), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n315), .A2(new_n651), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n316), .A2(new_n347), .A3(new_n829), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n315), .B(new_n651), .C1(new_n292), .C2(new_n635), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n828), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT38), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT37), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n431), .B2(KEYINPUT101), .ZN(new_n836));
  AND3_X1   g0636(.A1(new_n399), .A2(KEYINPUT101), .A3(new_n427), .ZN(new_n837));
  INV_X1    g0637(.A(new_n649), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n427), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n438), .ZN(new_n840));
  NOR3_X1   g0640(.A1(new_n836), .A2(new_n837), .A3(new_n840), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n839), .A2(new_n438), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n835), .B1(new_n842), .B2(new_n428), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n839), .B1(new_n639), .B2(new_n636), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n834), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT101), .ZN(new_n847));
  AOI21_X1  g0647(.A(KEYINPUT37), .B1(new_n428), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n431), .A2(KEYINPUT101), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n848), .A2(new_n842), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(KEYINPUT16), .B1(new_n407), .B2(new_n411), .ZN(new_n851));
  OAI21_X1  g0651(.A(KEYINPUT100), .B1(new_n851), .B2(new_n302), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n407), .A2(new_n411), .A3(KEYINPUT16), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n414), .B1(new_n419), .B2(new_n420), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT100), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n854), .A2(new_n855), .A3(new_n301), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n852), .A2(new_n853), .A3(new_n856), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n857), .A2(new_n426), .B1(new_n397), .B2(new_n398), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n649), .B1(new_n857), .B2(new_n426), .ZN(new_n859));
  INV_X1    g0659(.A(new_n438), .ZN(new_n860));
  NOR3_X1   g0660(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n850), .B1(new_n861), .B2(new_n835), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n639), .A2(new_n636), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n859), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n862), .A2(new_n864), .A3(KEYINPUT38), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n846), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(KEYINPUT40), .ZN(new_n867));
  OR3_X1    g0667(.A1(new_n833), .A2(KEYINPUT103), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n857), .A2(new_n426), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n869), .A2(new_n838), .B1(new_n434), .B2(new_n436), .ZN(new_n870));
  INV_X1    g0670(.A(new_n858), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n835), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n859), .ZN(new_n873));
  OAI22_X1  g0673(.A1(new_n872), .A2(new_n841), .B1(new_n440), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n834), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n865), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n828), .A2(new_n876), .A3(new_n832), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT40), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT103), .B1(new_n833), .B2(new_n867), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n868), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n704), .A2(new_n827), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n442), .A2(new_n882), .ZN(new_n883));
  XOR2_X1   g0683(.A(new_n881), .B(new_n883), .Z(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(G330), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n688), .A2(new_n348), .A3(new_n441), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n641), .A2(new_n886), .A3(new_n633), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n885), .B(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n316), .A2(new_n651), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT39), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n846), .A2(new_n890), .A3(new_n865), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n890), .B1(new_n875), .B2(new_n865), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n889), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n640), .A2(new_n649), .ZN(new_n894));
  INV_X1    g0694(.A(new_n788), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n795), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n896), .A2(new_n876), .A3(new_n832), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n893), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT102), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n893), .A2(KEYINPUT102), .A3(new_n894), .A4(new_n897), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n888), .B(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n903), .B1(new_n211), .B2(new_n645), .ZN(new_n904));
  OAI211_X1 g0704(.A(G20), .B(new_n209), .C1(new_n591), .C2(KEYINPUT35), .ZN(new_n905));
  AOI211_X1 g0705(.A(new_n221), .B(new_n905), .C1(KEYINPUT35), .C2(new_n591), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n906), .B(KEYINPUT36), .Z(new_n907));
  NOR3_X1   g0707(.A1(new_n679), .A2(new_n202), .A3(new_n400), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n226), .A2(G50), .ZN(new_n909));
  OAI211_X1 g0709(.A(G1), .B(new_n214), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n904), .A2(new_n907), .A3(new_n910), .ZN(G367));
  NAND2_X1  g0711(.A1(new_n627), .A2(new_n651), .ZN(new_n912));
  XOR2_X1   g0712(.A(new_n912), .B(KEYINPUT104), .Z(new_n913));
  MUX2_X1   g0713(.A(new_n613), .B(new_n628), .S(new_n913), .Z(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n735), .ZN(new_n915));
  INV_X1    g0715(.A(new_n725), .ZN(new_n916));
  OAI221_X1 g0716(.A(new_n736), .B1(new_n216), .B2(new_n320), .C1(new_n240), .C2(new_n916), .ZN(new_n917));
  OAI221_X1 g0717(.A(new_n253), .B1(new_n752), .B2(new_n351), .C1(new_n780), .C2(new_n747), .ZN(new_n918));
  INV_X1    g0718(.A(new_n738), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(G68), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n776), .B2(new_n804), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n758), .A2(G77), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(G137), .B2(new_n767), .ZN(new_n925));
  OAI221_X1 g0725(.A(new_n925), .B1(new_n309), .B2(new_n743), .C1(new_n770), .C2(new_n816), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT46), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n747), .A2(new_n927), .A3(new_n221), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n743), .A2(new_n817), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n927), .B1(new_n747), .B2(new_n221), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT108), .ZN(new_n931));
  OAI221_X1 g0731(.A(new_n329), .B1(new_n465), .B2(new_n752), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  AOI211_X1 g0732(.A(new_n929), .B(new_n932), .C1(new_n931), .C2(new_n930), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n776), .A2(new_n744), .B1(new_n738), .B2(new_n587), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n757), .A2(new_n586), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n934), .B(new_n935), .C1(G317), .C2(new_n767), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n933), .B(new_n936), .C1(new_n739), .C2(new_n816), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n926), .B1(new_n928), .B2(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT47), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n732), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n915), .A2(new_n721), .A3(new_n917), .A4(new_n940), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n600), .B(new_n605), .C1(new_n599), .C2(new_n652), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n616), .A2(new_n651), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n669), .A2(new_n671), .A3(new_n945), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n946), .A2(KEYINPUT107), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(KEYINPUT107), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT44), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n947), .A2(new_n948), .A3(KEYINPUT44), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n945), .B1(new_n669), .B2(new_n671), .ZN(new_n953));
  XOR2_X1   g0753(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n954));
  XNOR2_X1  g0754(.A(new_n953), .B(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n951), .A2(new_n952), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n664), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n644), .A2(new_n652), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n662), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n666), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n657), .B(new_n960), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n713), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n951), .A2(new_n665), .A3(new_n952), .A4(new_n955), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n957), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n714), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n676), .B(KEYINPUT41), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n720), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n666), .A2(new_n945), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT42), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n605), .B1(new_n942), .B2(new_n521), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n652), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n974), .A2(KEYINPUT105), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(KEYINPUT105), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT43), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n977), .B1(new_n978), .B2(new_n914), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n664), .A2(new_n944), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n914), .B(KEYINPUT43), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(new_n975), .B2(new_n976), .ZN(new_n983));
  OR3_X1    g0783(.A1(new_n979), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n981), .B1(new_n979), .B2(new_n983), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n941), .B1(new_n969), .B2(new_n986), .ZN(G387));
  INV_X1    g0787(.A(KEYINPUT111), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n722), .B1(new_n662), .B2(new_n735), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n237), .A2(new_n268), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n677), .B(new_n268), .C1(new_n226), .C2(new_n202), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT50), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n317), .B2(G50), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n318), .A2(KEYINPUT50), .A3(new_n309), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n991), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NOR3_X1   g0795(.A1(new_n990), .A2(new_n916), .A3(new_n995), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n728), .A2(new_n677), .B1(G107), .B2(new_n216), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT109), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n736), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n989), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n556), .A2(new_n919), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n309), .B2(new_n752), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT110), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n253), .B1(new_n743), .B2(new_n226), .C1(new_n202), .C2(new_n747), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n757), .A2(new_n586), .B1(new_n770), .B2(new_n776), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n1004), .B(new_n1005), .C1(G150), .C2(new_n767), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1003), .B(new_n1006), .C1(new_n317), .C2(new_n763), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n802), .A2(G303), .B1(G322), .B2(new_n750), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n816), .B2(new_n744), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(G317), .B2(new_n753), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT48), .Z(new_n1011));
  NAND2_X1  g0811(.A1(new_n919), .A2(G283), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n747), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(G294), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1011), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT49), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n253), .B1(new_n767), .B2(G326), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n757), .A2(new_n221), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1007), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1000), .B1(new_n1022), .B2(new_n732), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n961), .A2(new_n719), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n676), .B1(new_n713), .B2(new_n961), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n962), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n988), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1025), .A2(new_n1027), .A3(new_n988), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(G393));
  NAND3_X1  g0831(.A1(new_n957), .A2(KEYINPUT112), .A3(new_n964), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n964), .A2(KEYINPUT112), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n718), .B(new_n965), .C1(new_n1034), .C2(new_n963), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n945), .A2(new_n735), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n816), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(G303), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n753), .A2(G311), .B1(G317), .B2(new_n750), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT52), .Z(new_n1040));
  NAND2_X1  g0840(.A1(new_n767), .A2(G322), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n329), .B1(new_n738), .B2(new_n221), .C1(new_n739), .C2(new_n743), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n1042), .B(new_n773), .C1(G283), .C2(new_n1013), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1038), .A2(new_n1040), .A3(new_n1041), .A4(new_n1043), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n253), .B1(new_n743), .B2(new_n317), .C1(new_n226), .C2(new_n747), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1045), .B(new_n811), .C1(G77), .C2(new_n919), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n804), .B2(new_n766), .C1(new_n816), .C2(new_n309), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n753), .A2(G159), .B1(G150), .B2(new_n750), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT51), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1044), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n722), .B1(new_n1050), .B2(new_n732), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n736), .B1(new_n586), .B2(new_n216), .C1(new_n248), .C2(new_n916), .ZN(new_n1052));
  AND3_X1   g0852(.A1(new_n1036), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(new_n1034), .B2(new_n720), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1035), .A2(new_n1054), .ZN(G390));
  NAND2_X1  g0855(.A1(new_n1013), .A2(G150), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT53), .ZN(new_n1057));
  INV_X1    g0857(.A(G125), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n309), .A2(new_n757), .B1(new_n766), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(G128), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n776), .A2(new_n1060), .B1(new_n738), .B2(new_n770), .ZN(new_n1061));
  XOR2_X1   g0861(.A(KEYINPUT54), .B(G143), .Z(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n253), .B1(new_n1063), .B2(new_n743), .ZN(new_n1064));
  NOR4_X1   g0864(.A1(new_n1057), .A2(new_n1059), .A3(new_n1061), .A4(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(G137), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1065), .B1(new_n800), .B2(new_n752), .C1(new_n1066), .C2(new_n816), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n776), .A2(new_n817), .B1(new_n738), .B2(new_n202), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n766), .A2(new_n739), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n329), .B1(new_n743), .B2(new_n586), .C1(new_n774), .C2(new_n747), .ZN(new_n1070));
  NOR4_X1   g0870(.A1(new_n1068), .A2(new_n799), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1071), .B1(new_n221), .B2(new_n752), .C1(new_n816), .C2(new_n587), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n731), .B1(new_n1067), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n317), .B2(new_n821), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n874), .A2(new_n834), .ZN(new_n1075));
  AOI21_X1  g0875(.A(KEYINPUT38), .B1(new_n862), .B2(new_n864), .ZN(new_n1076));
  OAI21_X1  g0876(.A(KEYINPUT39), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n846), .A2(new_n890), .A3(new_n865), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n721), .B(new_n1074), .C1(new_n1079), .C2(new_n734), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n790), .A2(new_n342), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n685), .A2(new_n652), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n895), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT113), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1082), .A2(KEYINPUT113), .A3(new_n895), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1085), .A2(new_n832), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n889), .B1(new_n865), .B2(new_n846), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n795), .A2(new_n895), .B1(new_n830), .B2(new_n831), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1077), .B(new_n1078), .C1(new_n1090), .C2(new_n889), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n711), .A2(new_n791), .A3(new_n832), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  AND3_X1   g0893(.A1(new_n1089), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n828), .A2(G330), .A3(new_n832), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1080), .B1(new_n1098), .B2(new_n719), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n609), .A2(new_n529), .A3(new_n652), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n1100), .A2(KEYINPUT31), .B1(new_n651), .B2(new_n700), .ZN(new_n1101));
  OAI211_X1 g0901(.A(G330), .B(new_n791), .C1(new_n1101), .C2(new_n826), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n830), .A2(new_n831), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1092), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  AND3_X1   g0907(.A1(new_n709), .A2(KEYINPUT31), .A3(new_n651), .ZN(new_n1108));
  OAI211_X1 g0908(.A(G330), .B(new_n791), .C1(new_n1101), .C2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n1103), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(KEYINPUT114), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT114), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1109), .A2(new_n1103), .A3(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1111), .A2(new_n1095), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1107), .B1(new_n1114), .B2(new_n896), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n348), .A2(new_n441), .A3(new_n882), .A4(G330), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n641), .A2(new_n886), .A3(new_n1116), .A4(new_n633), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1098), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n676), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n1111), .A2(new_n1095), .A3(new_n1113), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n896), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1106), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1117), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n1098), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1099), .B1(new_n1120), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(G378));
  NAND4_X1  g0928(.A1(new_n868), .A2(G330), .A3(new_n879), .A4(new_n880), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n355), .A2(new_n649), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT116), .ZN(new_n1134));
  OR2_X1    g0934(.A1(new_n382), .A2(new_n1134), .ZN(new_n1135));
  AOI211_X1 g0935(.A(KEYINPUT116), .B(new_n371), .C1(new_n377), .C2(new_n381), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1133), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n382), .A2(new_n1134), .ZN(new_n1139));
  NOR3_X1   g0939(.A1(new_n1139), .A2(new_n1136), .A3(new_n1132), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1131), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1135), .A2(new_n1137), .A3(new_n1133), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1132), .B1(new_n1139), .B2(new_n1136), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1142), .A2(new_n1143), .A3(new_n1130), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n900), .A2(new_n901), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1145), .B1(new_n900), .B2(new_n901), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1129), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1145), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1079), .A2(new_n889), .B1(new_n876), .B2(new_n1090), .ZN(new_n1150));
  AOI21_X1  g0950(.A(KEYINPUT102), .B1(new_n1150), .B2(new_n894), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n901), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1149), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1129), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n900), .A2(new_n901), .A3(new_n1145), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1124), .B1(new_n1098), .B2(new_n1115), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1148), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT57), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1148), .A2(new_n1156), .A3(new_n1157), .A4(KEYINPUT57), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1160), .A2(new_n718), .A3(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1148), .A2(new_n1156), .A3(new_n720), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n757), .A2(new_n780), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n920), .B1(new_n221), .B2(new_n776), .C1(new_n766), .C2(new_n817), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n1164), .B(new_n1165), .C1(G97), .C2(new_n764), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n263), .B(new_n329), .C1(new_n747), .C2(new_n202), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT115), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n556), .A2(new_n802), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1166), .B(new_n1169), .C1(new_n1168), .C2(new_n1167), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(G107), .B2(new_n753), .ZN(new_n1171));
  XOR2_X1   g0971(.A(new_n1171), .B(KEYINPUT58), .Z(new_n1172));
  OAI21_X1  g0972(.A(new_n309), .B1(new_n327), .B2(G41), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n776), .A2(new_n1058), .B1(new_n351), .B2(new_n738), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n1063), .A2(new_n747), .B1(new_n743), .B2(new_n1066), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1174), .B(new_n1175), .C1(new_n764), .C2(G132), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n1060), .B2(new_n752), .ZN(new_n1177));
  OR2_X1    g0977(.A1(new_n1177), .A2(KEYINPUT59), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(KEYINPUT59), .ZN(new_n1179));
  AOI21_X1  g0979(.A(G33), .B1(new_n758), .B2(G159), .ZN(new_n1180));
  AOI21_X1  g0980(.A(G41), .B1(new_n767), .B2(G124), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .A4(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1172), .A2(new_n1173), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n722), .B1(new_n1183), .B2(new_n732), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1184), .B1(G50), .B2(new_n820), .C1(new_n1145), .C2(new_n734), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1163), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1162), .A2(new_n1186), .ZN(G375));
  OAI211_X1 g0987(.A(new_n1117), .B(new_n1106), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1125), .A2(new_n968), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n722), .B1(new_n821), .B2(new_n226), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n1190), .B(KEYINPUT117), .Z(new_n1191));
  NOR2_X1   g0991(.A1(new_n832), .A2(new_n734), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1037), .A2(G116), .B1(G107), .B2(new_n802), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n739), .B2(new_n776), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT118), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n766), .A2(new_n465), .B1(new_n586), .B2(new_n747), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT119), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n253), .B(new_n1197), .C1(G283), .C2(new_n753), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1195), .A2(new_n923), .A3(new_n1001), .A4(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n752), .A2(new_n1066), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n766), .A2(new_n1060), .B1(new_n770), .B2(new_n747), .ZN(new_n1201));
  XOR2_X1   g1001(.A(new_n1201), .B(KEYINPUT120), .Z(new_n1202));
  OAI22_X1  g1002(.A1(new_n776), .A2(new_n800), .B1(new_n738), .B2(new_n309), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n253), .B1(new_n743), .B2(new_n351), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(new_n1164), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1202), .B(new_n1205), .C1(new_n816), .C2(new_n1063), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1199), .B1(new_n1200), .B2(new_n1206), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1191), .B(new_n1192), .C1(new_n732), .C2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n1123), .B2(new_n720), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1189), .A2(new_n1209), .ZN(G381));
  AND2_X1   g1010(.A1(new_n1186), .A2(new_n1127), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n1162), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1029), .A2(new_n785), .A3(new_n723), .A4(new_n1030), .ZN(new_n1213));
  OR3_X1    g1013(.A1(new_n1213), .A2(G381), .A3(G384), .ZN(new_n1214));
  NOR3_X1   g1014(.A1(new_n1214), .A2(G387), .A3(G390), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT121), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1212), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n1216), .B2(new_n1215), .ZN(G407));
  NAND2_X1  g1018(.A1(new_n650), .A2(G213), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1219), .B(KEYINPUT122), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  OAI211_X1 g1021(.A(G407), .B(G213), .C1(new_n1212), .C2(new_n1221), .ZN(G409));
  INV_X1    g1022(.A(KEYINPUT124), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT60), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1188), .A2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1115), .A2(KEYINPUT60), .A3(new_n1117), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1225), .A2(new_n1125), .A3(new_n718), .A4(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1227), .A2(G384), .A3(new_n1209), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(G384), .B1(new_n1227), .B2(new_n1209), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1223), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1227), .A2(new_n1209), .ZN(new_n1232));
  INV_X1    g1032(.A(G384), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1234), .A2(KEYINPUT124), .A3(new_n1228), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1231), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(G375), .A2(G378), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1148), .A2(new_n1156), .A3(new_n1157), .A4(new_n968), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1186), .A2(new_n1127), .A3(new_n1238), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1236), .A2(new_n1237), .A3(new_n1221), .A4(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT61), .B1(new_n1240), .B2(KEYINPUT62), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1220), .A2(G2897), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(new_n1236), .B2(new_n1243), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1237), .A2(new_n1221), .A3(new_n1239), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1237), .A2(KEYINPUT123), .A3(new_n1239), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT123), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1127), .B1(new_n1162), .B2(new_n1186), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1239), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1249), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1248), .A2(new_n1252), .A3(new_n1221), .A4(new_n1236), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1241), .B(new_n1247), .C1(new_n1253), .C2(KEYINPUT62), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1030), .ZN(new_n1255));
  OAI21_X1  g1055(.A(G396), .B1(new_n1255), .B2(new_n1028), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1213), .A2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1257), .A2(new_n1035), .A3(new_n1054), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1257), .B1(new_n1035), .B2(new_n1054), .ZN(new_n1260));
  OAI21_X1  g1060(.A(G387), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(G390), .A2(new_n1213), .A3(new_n1256), .ZN(new_n1262));
  INV_X1    g1062(.A(G387), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1262), .A2(new_n1263), .A3(new_n1258), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1261), .A2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1254), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT63), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1253), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT125), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1253), .A2(KEYINPUT125), .A3(new_n1267), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT61), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1261), .A2(new_n1264), .A3(new_n1273), .ZN(new_n1274));
  OR2_X1    g1074(.A1(new_n1274), .A2(KEYINPUT126), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1248), .A2(new_n1252), .A3(new_n1221), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1245), .ZN(new_n1277));
  OR2_X1    g1077(.A1(new_n1240), .A2(new_n1267), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1274), .A2(KEYINPUT126), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1275), .A2(new_n1277), .A3(new_n1278), .A4(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1266), .B1(new_n1272), .B2(new_n1280), .ZN(G405));
  XNOR2_X1  g1081(.A(new_n1265), .B(KEYINPUT127), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1250), .B1(new_n1162), .B2(new_n1211), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1236), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1284), .B1(new_n1242), .B2(new_n1283), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1282), .B(new_n1285), .ZN(G402));
endmodule


