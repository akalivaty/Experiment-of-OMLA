//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 0 0 1 0 0 1 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 1 1 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n548, new_n549,
    new_n550, new_n551, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n563, new_n565, new_n566,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n613, new_n615, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1134, new_n1135;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT65), .Z(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT66), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G125), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT67), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n459), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(new_n466), .A3(KEYINPUT67), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n458), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  XNOR2_X1  g044(.A(new_n469), .B(KEYINPUT68), .ZN(new_n470));
  OAI21_X1  g045(.A(G2105), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT69), .B(G2104), .ZN(new_n472));
  OAI211_X1 g047(.A(G137), .B(new_n465), .C1(new_n472), .C2(new_n462), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(G101), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n471), .A2(new_n477), .ZN(G160));
  OR2_X1    g053(.A1(new_n472), .A2(new_n462), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(new_n465), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(new_n476), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(G124), .ZN(new_n483));
  OR3_X1    g058(.A1(new_n482), .A2(KEYINPUT70), .A3(new_n483), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(new_n476), .B2(G112), .ZN(new_n485));
  INV_X1    g060(.A(G100), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(new_n476), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n480), .A2(G2105), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(new_n488), .B2(G136), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT70), .B1(new_n482), .B2(new_n483), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n484), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT71), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  OAI211_X1 g068(.A(G126), .B(new_n465), .C1(new_n472), .C2(new_n462), .ZN(new_n494));
  NAND2_X1  g069(.A1(G114), .A2(G2104), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  AND2_X1   g072(.A1(KEYINPUT4), .A2(G138), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n465), .B(new_n498), .C1(new_n472), .C2(new_n462), .ZN(new_n499));
  NAND2_X1  g074(.A1(G102), .A2(G2104), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(new_n476), .ZN(new_n502));
  AND3_X1   g077(.A1(new_n465), .A2(new_n466), .A3(KEYINPUT67), .ZN(new_n503));
  AOI21_X1  g078(.A(KEYINPUT67), .B1(new_n465), .B2(new_n466), .ZN(new_n504));
  OAI211_X1 g079(.A(G138), .B(new_n476), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n497), .A2(new_n502), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT72), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n476), .B1(new_n494), .B2(new_n495), .ZN(new_n510));
  AOI21_X1  g085(.A(G2105), .B1(new_n499), .B2(new_n500), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT72), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(new_n513), .A3(new_n507), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n509), .A2(new_n514), .ZN(G164));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n517), .B2(KEYINPUT73), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT73), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n519), .A2(KEYINPUT5), .A3(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  XOR2_X1   g097(.A(KEYINPUT6), .B(G651), .Z(new_n523));
  OAI21_X1  g098(.A(KEYINPUT74), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT74), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT6), .B(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n521), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G88), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n530));
  INV_X1    g105(.A(G651), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n526), .A2(G50), .A3(G543), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n529), .A2(new_n532), .A3(new_n533), .ZN(G303));
  INV_X1    g109(.A(G303), .ZN(G166));
  NAND2_X1  g110(.A1(new_n528), .A2(G89), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT75), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n523), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n526), .A2(KEYINPUT75), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n538), .A2(G543), .A3(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G51), .ZN(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT7), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n545));
  NAND4_X1  g120(.A1(new_n536), .A2(new_n542), .A3(new_n544), .A4(new_n545), .ZN(G286));
  INV_X1    g121(.A(G286), .ZN(G168));
  NAND2_X1  g122(.A1(new_n528), .A2(G90), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(new_n531), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n541), .A2(G52), .ZN(new_n551));
  AND3_X1   g126(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(G171));
  NAND2_X1  g127(.A1(new_n524), .A2(new_n527), .ZN(new_n553));
  INV_X1    g128(.A(G81), .ZN(new_n554));
  INV_X1    g129(.A(G43), .ZN(new_n555));
  OAI22_X1  g130(.A1(new_n553), .A2(new_n554), .B1(new_n555), .B2(new_n540), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT76), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n558), .A2(new_n531), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  AND3_X1   g137(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G36), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n563), .A2(new_n566), .ZN(G188));
  NAND4_X1  g142(.A1(new_n538), .A2(G53), .A3(G543), .A4(new_n539), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT77), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AND2_X1   g146(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n569), .A2(new_n570), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n571), .B1(new_n568), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT78), .ZN(new_n575));
  OR3_X1    g150(.A1(new_n572), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n572), .B2(new_n574), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  XOR2_X1   g154(.A(KEYINPUT79), .B(G65), .Z(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n522), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n528), .A2(G91), .B1(G651), .B2(new_n581), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G299));
  INV_X1    g159(.A(G171), .ZN(G301));
  NAND2_X1  g160(.A1(new_n528), .A2(G87), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n541), .A2(G49), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G288));
  AND3_X1   g164(.A1(new_n526), .A2(G48), .A3(G543), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n521), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G86), .ZN(new_n593));
  OAI221_X1 g168(.A(new_n591), .B1(new_n531), .B2(new_n592), .C1(new_n553), .C2(new_n593), .ZN(G305));
  AOI22_X1  g169(.A1(new_n528), .A2(G85), .B1(G47), .B2(new_n541), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n531), .B2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  INV_X1    g173(.A(G54), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n521), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n600));
  OAI22_X1  g175(.A1(new_n540), .A2(new_n599), .B1(new_n531), .B2(new_n600), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT80), .ZN(new_n602));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  OAI21_X1  g178(.A(KEYINPUT10), .B1(new_n553), .B2(new_n603), .ZN(new_n604));
  OR3_X1    g179(.A1(new_n553), .A2(KEYINPUT10), .A3(new_n603), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n602), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n598), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n598), .B1(new_n607), .B2(G868), .ZN(G321));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(new_n583), .B2(G868), .ZN(G297));
  OAI21_X1  g186(.A(new_n610), .B1(new_n583), .B2(G868), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n607), .B1(new_n613), .B2(G860), .ZN(G148));
  NOR2_X1   g189(.A1(new_n606), .A2(G559), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G868), .B2(new_n561), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI21_X1  g194(.A(G2105), .B1(new_n464), .B2(new_n467), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(new_n472), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT12), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2100), .ZN(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n625), .A2(KEYINPUT81), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(KEYINPUT81), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n626), .B(new_n627), .C1(G111), .C2(new_n476), .ZN(new_n628));
  INV_X1    g203(.A(new_n488), .ZN(new_n629));
  INV_X1    g204(.A(G135), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n631), .B1(G123), .B2(new_n481), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2096), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n624), .A2(new_n633), .ZN(G156));
  XOR2_X1   g209(.A(KEYINPUT15), .B(G2435), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2438), .ZN(new_n636));
  XOR2_X1   g211(.A(G2427), .B(G2430), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT83), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n636), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(KEYINPUT14), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2451), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(G2454), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n640), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n646), .B(new_n647), .Z(new_n648));
  AND2_X1   g223(.A1(new_n648), .A2(G14), .ZN(G401));
  XNOR2_X1  g224(.A(G2084), .B(G2090), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT84), .Z(new_n651));
  XOR2_X1   g226(.A(G2067), .B(G2678), .Z(new_n652));
  NOR2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2072), .B(G2078), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT18), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n654), .B(KEYINPUT17), .Z(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n651), .B2(new_n652), .ZN(new_n658));
  INV_X1    g233(.A(new_n652), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n659), .A2(new_n654), .ZN(new_n660));
  AOI211_X1 g235(.A(new_n653), .B(new_n658), .C1(new_n651), .C2(new_n660), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT85), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2096), .B(G2100), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(G227));
  XOR2_X1   g240(.A(G1956), .B(G2474), .Z(new_n666));
  XOR2_X1   g241(.A(G1961), .B(G1966), .Z(new_n667));
  NOR2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1971), .B(G1976), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n666), .A2(new_n667), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT20), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n672), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n669), .A2(new_n671), .A3(new_n673), .ZN(new_n677));
  OAI211_X1 g252(.A(new_n676), .B(new_n677), .C1(new_n675), .C2(new_n674), .ZN(new_n678));
  XOR2_X1   g253(.A(G1981), .B(G1986), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G1991), .B(G1996), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT86), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n682), .B(new_n684), .Z(G229));
  MUX2_X1   g260(.A(G6), .B(G305), .S(G16), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT89), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT32), .B(G1981), .Z(new_n688));
  XOR2_X1   g263(.A(new_n687), .B(new_n688), .Z(new_n689));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G22), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(G166), .B2(new_n690), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(G1971), .Z(new_n693));
  NOR2_X1   g268(.A1(G16), .A2(G23), .ZN(new_n694));
  INV_X1    g269(.A(G288), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n694), .B1(new_n695), .B2(G16), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT33), .B(G1976), .Z(new_n697));
  XOR2_X1   g272(.A(new_n696), .B(new_n697), .Z(new_n698));
  NAND3_X1  g273(.A1(new_n689), .A2(new_n693), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(KEYINPUT34), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT90), .ZN(new_n701));
  INV_X1    g276(.A(G25), .ZN(new_n702));
  OAI21_X1  g277(.A(KEYINPUT87), .B1(new_n702), .B2(G29), .ZN(new_n703));
  OR3_X1    g278(.A1(new_n702), .A2(KEYINPUT87), .A3(G29), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n481), .A2(G119), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n488), .A2(G131), .ZN(new_n706));
  NOR2_X1   g281(.A1(G95), .A2(G2105), .ZN(new_n707));
  OAI21_X1  g282(.A(G2104), .B1(new_n476), .B2(G107), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n705), .B(new_n706), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT88), .ZN(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n703), .B(new_n704), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT35), .B(G1991), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n712), .B(new_n713), .Z(new_n714));
  OAI211_X1 g289(.A(new_n701), .B(new_n714), .C1(KEYINPUT34), .C2(new_n699), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT91), .B(KEYINPUT36), .Z(new_n716));
  MUX2_X1   g291(.A(G24), .B(G290), .S(G16), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(G1986), .ZN(new_n718));
  OR3_X1    g293(.A1(new_n715), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n716), .B1(new_n715), .B2(new_n718), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT92), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G4), .B2(G16), .ZN(new_n722));
  OR3_X1    g297(.A1(new_n721), .A2(G4), .A3(G16), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n722), .B(new_n723), .C1(new_n606), .C2(new_n690), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G1348), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n632), .A2(G29), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT94), .ZN(new_n727));
  NOR2_X1   g302(.A1(G5), .A2(G16), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G171), .B2(G16), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G1961), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT30), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(G28), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(G28), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n732), .A2(new_n733), .A3(new_n711), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n727), .A2(new_n730), .A3(new_n734), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT31), .B(G11), .Z(new_n736));
  NAND2_X1  g311(.A1(new_n690), .A2(G21), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G168), .B2(new_n690), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G1966), .ZN(new_n739));
  NOR3_X1   g314(.A1(new_n735), .A2(new_n736), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT95), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n561), .A2(G16), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G16), .B2(G19), .ZN(new_n743));
  INV_X1    g318(.A(G1341), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n711), .A2(G27), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G164), .B2(new_n711), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n743), .A2(new_n744), .B1(G2078), .B2(new_n746), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n711), .A2(G26), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n481), .A2(G128), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n488), .A2(G140), .ZN(new_n750));
  NOR2_X1   g325(.A1(G104), .A2(G2105), .ZN(new_n751));
  OAI21_X1  g326(.A(G2104), .B1(new_n476), .B2(G116), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n749), .B(new_n750), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n748), .B1(new_n753), .B2(G29), .ZN(new_n754));
  MUX2_X1   g329(.A(new_n748), .B(new_n754), .S(KEYINPUT28), .Z(new_n755));
  INV_X1    g330(.A(G2067), .ZN(new_n756));
  OR2_X1    g331(.A1(G29), .A2(G32), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n481), .A2(G129), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n488), .A2(G141), .ZN(new_n759));
  NAND3_X1  g334(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT26), .Z(new_n761));
  NAND3_X1  g336(.A1(new_n472), .A2(G105), .A3(new_n476), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT93), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n758), .A2(new_n759), .A3(new_n761), .A4(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n757), .B1(new_n764), .B2(new_n711), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT27), .B(G1996), .ZN(new_n766));
  OAI22_X1  g341(.A1(new_n755), .A2(new_n756), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  NOR2_X1   g343(.A1(G160), .A2(new_n711), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT24), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n770), .A2(G34), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(G34), .ZN(new_n772));
  AOI21_X1  g347(.A(G29), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(G2084), .B1(new_n769), .B2(new_n773), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n768), .B(new_n774), .C1(G1961), .C2(new_n729), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n767), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n741), .A2(new_n747), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n711), .A2(G35), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G162), .B2(new_n711), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT29), .ZN(new_n780));
  OAI22_X1  g355(.A1(new_n780), .A2(G2090), .B1(new_n744), .B2(new_n743), .ZN(new_n781));
  NOR3_X1   g356(.A1(new_n769), .A2(G2084), .A3(new_n773), .ZN(new_n782));
  OAI21_X1  g357(.A(G127), .B1(new_n503), .B2(new_n504), .ZN(new_n783));
  INV_X1    g358(.A(G115), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(new_n460), .ZN(new_n785));
  AOI22_X1  g360(.A1(G139), .A2(new_n488), .B1(new_n785), .B2(G2105), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n476), .A2(G103), .A3(G2104), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT25), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  MUX2_X1   g364(.A(G33), .B(new_n789), .S(G29), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G2072), .ZN(new_n791));
  NOR4_X1   g366(.A1(new_n777), .A2(new_n781), .A3(new_n782), .A4(new_n791), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n719), .A2(new_n720), .A3(new_n725), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n755), .A2(new_n756), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n780), .A2(G2090), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT96), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n690), .A2(KEYINPUT23), .A3(G20), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT23), .ZN(new_n799));
  INV_X1    g374(.A(G20), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(G16), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n798), .B(new_n801), .C1(new_n583), .C2(new_n690), .ZN(new_n802));
  INV_X1    g377(.A(G1956), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n797), .A2(new_n804), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT97), .Z(new_n806));
  NOR2_X1   g381(.A1(new_n746), .A2(G2078), .ZN(new_n807));
  NOR4_X1   g382(.A1(new_n793), .A2(new_n795), .A3(new_n806), .A4(new_n807), .ZN(G311));
  INV_X1    g383(.A(G311), .ZN(G150));
  AOI22_X1  g384(.A1(new_n528), .A2(G93), .B1(G55), .B2(new_n541), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT98), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n810), .B1(new_n531), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(G860), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT37), .Z(new_n815));
  OR2_X1    g390(.A1(new_n561), .A2(new_n813), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n561), .A2(new_n813), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n606), .A2(new_n613), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n815), .B1(new_n822), .B2(G860), .ZN(G145));
  XNOR2_X1  g398(.A(G160), .B(KEYINPUT99), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n492), .B(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(new_n632), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(new_n764), .ZN(new_n827));
  AOI21_X1  g402(.A(KEYINPUT4), .B1(new_n620), .B2(G138), .ZN(new_n828));
  NOR3_X1   g403(.A1(new_n828), .A2(new_n510), .A3(new_n511), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n789), .B(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n753), .B(new_n622), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n481), .A2(G130), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n488), .A2(G142), .ZN(new_n834));
  NOR2_X1   g409(.A1(G106), .A2(G2105), .ZN(new_n835));
  OAI21_X1  g410(.A(G2104), .B1(new_n476), .B2(G118), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n833), .B(new_n834), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n710), .B(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n832), .B(new_n838), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n827), .B(new_n839), .Z(new_n840));
  NOR2_X1   g415(.A1(new_n840), .A2(G37), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT40), .Z(G395));
  NOR2_X1   g417(.A1(new_n813), .A2(G868), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT100), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n606), .B1(new_n583), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(new_n844), .B2(new_n583), .ZN(new_n846));
  NAND3_X1  g421(.A1(G299), .A2(KEYINPUT100), .A3(new_n606), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT41), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n818), .B(new_n616), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(new_n850), .B2(new_n848), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT102), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XOR2_X1   g429(.A(G303), .B(G305), .Z(new_n855));
  XNOR2_X1  g430(.A(G290), .B(G288), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n855), .B1(new_n857), .B2(KEYINPUT101), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n857), .A2(KEYINPUT101), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n854), .B1(KEYINPUT42), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(KEYINPUT42), .B2(new_n860), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n852), .A2(new_n853), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n862), .B(new_n863), .Z(new_n864));
  AOI21_X1  g439(.A(new_n843), .B1(new_n864), .B2(G868), .ZN(G295));
  AOI21_X1  g440(.A(new_n843), .B1(new_n864), .B2(G868), .ZN(G331));
  INV_X1    g441(.A(KEYINPUT44), .ZN(new_n867));
  INV_X1    g442(.A(new_n860), .ZN(new_n868));
  NAND2_X1  g443(.A1(G171), .A2(KEYINPUT103), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT104), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(G286), .B1(G171), .B2(KEYINPUT103), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n871), .B(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n818), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n871), .B(new_n872), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(new_n818), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n849), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT105), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n876), .A2(new_n878), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n877), .A2(KEYINPUT105), .A3(new_n818), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n848), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n868), .B1(new_n880), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n849), .A2(new_n883), .A3(new_n882), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n879), .A2(new_n848), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n886), .A2(new_n887), .A3(new_n860), .ZN(new_n888));
  INV_X1    g463(.A(G37), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n885), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n867), .B1(new_n890), .B2(KEYINPUT43), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n886), .A2(new_n887), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n868), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT43), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n893), .A2(new_n894), .A3(new_n889), .A4(new_n888), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT106), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n888), .A2(new_n889), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n898), .A2(KEYINPUT106), .A3(new_n894), .A4(new_n893), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n891), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(KEYINPUT107), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT107), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n891), .A2(new_n897), .A3(new_n899), .A4(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n898), .A2(new_n893), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT43), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n906), .B1(KEYINPUT43), .B2(new_n890), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n867), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(KEYINPUT108), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT108), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n904), .A2(new_n911), .A3(new_n908), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(G397));
  NAND3_X1  g488(.A1(new_n471), .A2(new_n477), .A3(G40), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT109), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n471), .A2(new_n477), .A3(KEYINPUT109), .A4(G40), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT45), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n919), .B1(new_n829), .B2(G1384), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n710), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n923), .A2(new_n713), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n753), .B(new_n756), .ZN(new_n925));
  INV_X1    g500(.A(G1996), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n764), .B(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n924), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  OR2_X1    g503(.A1(new_n753), .A2(G2067), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n922), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n925), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n921), .B1(new_n931), .B2(new_n764), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT46), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n933), .B1(new_n922), .B2(G1996), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n921), .A2(KEYINPUT46), .A3(new_n926), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n932), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  XOR2_X1   g511(.A(new_n936), .B(KEYINPUT47), .Z(new_n937));
  INV_X1    g512(.A(new_n924), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n923), .A2(new_n713), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n938), .A2(new_n939), .A3(new_n925), .A4(new_n927), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n921), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n922), .A2(G1986), .A3(G290), .ZN(new_n942));
  XNOR2_X1  g517(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n942), .B(new_n943), .ZN(new_n944));
  AOI211_X1 g519(.A(new_n930), .B(new_n937), .C1(new_n941), .C2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(G286), .A2(G8), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n946), .A2(KEYINPUT120), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n947), .A2(KEYINPUT51), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT116), .ZN(new_n949));
  INV_X1    g524(.A(G1384), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT45), .B1(new_n508), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n949), .B1(new_n918), .B2(new_n951), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n920), .A2(KEYINPUT116), .A3(new_n916), .A4(new_n917), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n509), .A2(new_n514), .A3(KEYINPUT45), .A4(new_n950), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(G1966), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n508), .A2(new_n950), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n916), .B(new_n917), .C1(new_n958), .C2(KEYINPUT50), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n509), .A2(new_n950), .A3(new_n514), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n959), .B1(KEYINPUT50), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(G2084), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n957), .A2(new_n963), .ZN(new_n964));
  OAI211_X1 g539(.A(G8), .B(new_n948), .C1(new_n964), .C2(G286), .ZN(new_n965));
  INV_X1    g540(.A(new_n948), .ZN(new_n966));
  AOI22_X1  g541(.A1(new_n955), .A2(new_n956), .B1(new_n961), .B2(new_n962), .ZN(new_n967));
  INV_X1    g542(.A(G8), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n946), .B(new_n966), .C1(new_n967), .C2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n964), .A2(G8), .A3(G286), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n965), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT121), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n965), .A2(new_n969), .A3(KEYINPUT121), .A4(new_n970), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(KEYINPUT122), .B(KEYINPUT54), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n508), .A2(KEYINPUT45), .A3(new_n950), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n977), .A2(new_n916), .A3(new_n917), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n978), .B1(new_n919), .B2(new_n960), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT110), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n960), .A2(new_n919), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n977), .A2(new_n916), .A3(new_n917), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT110), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G2078), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n980), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT53), .ZN(new_n988));
  INV_X1    g563(.A(G1961), .ZN(new_n989));
  INV_X1    g564(.A(new_n961), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n987), .A2(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n914), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n988), .A2(G2078), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n920), .A2(new_n992), .A3(new_n977), .A4(new_n993), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n991), .A2(G301), .A3(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n952), .A2(new_n953), .A3(new_n954), .A4(new_n993), .ZN(new_n996));
  AOI21_X1  g571(.A(G301), .B1(new_n991), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n976), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n991), .A2(G301), .A3(new_n996), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n987), .A2(new_n988), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n990), .A2(new_n989), .ZN(new_n1001));
  AND3_X1   g576(.A1(new_n1000), .A2(new_n1001), .A3(new_n994), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n999), .B(KEYINPUT54), .C1(new_n1002), .C2(G301), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n582), .B1(new_n572), .B2(new_n574), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT57), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT118), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n577), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n572), .A2(new_n574), .A3(new_n575), .ZN(new_n1008));
  OAI211_X1 g583(.A(KEYINPUT57), .B(new_n582), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n578), .A2(KEYINPUT118), .A3(KEYINPUT57), .A4(new_n582), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OR2_X1    g587(.A1(new_n960), .A2(KEYINPUT50), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n918), .B1(KEYINPUT50), .B2(new_n958), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n803), .ZN(new_n1016));
  XNOR2_X1  g591(.A(KEYINPUT56), .B(G2072), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n979), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1012), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1012), .B1(new_n1018), .B2(new_n1016), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n918), .A2(new_n958), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n756), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n959), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n960), .A2(KEYINPUT50), .ZN(new_n1025));
  AOI21_X1  g600(.A(G1348), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1027), .A2(new_n606), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1019), .B1(new_n1020), .B2(new_n1028), .ZN(new_n1029));
  OR2_X1    g604(.A1(new_n918), .A2(new_n958), .ZN(new_n1030));
  XOR2_X1   g605(.A(KEYINPUT58), .B(G1341), .Z(new_n1031));
  AOI22_X1  g606(.A1(new_n979), .A2(new_n926), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT59), .B1(new_n1032), .B2(new_n560), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(new_n983), .B2(G1996), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT59), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(new_n1036), .A3(new_n561), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1033), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT60), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1039), .B1(new_n1023), .B2(new_n1026), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT119), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n606), .A2(new_n1041), .ZN(new_n1042));
  OAI211_X1 g617(.A(KEYINPUT60), .B(new_n1022), .C1(new_n961), .C2(G1348), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n606), .A2(new_n1041), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1040), .B(new_n1042), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  OR2_X1    g620(.A1(new_n1043), .A2(new_n1042), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1038), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1019), .A2(KEYINPUT61), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT61), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1012), .A2(new_n1016), .A3(new_n1049), .A4(new_n1018), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1029), .B1(new_n1047), .B2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n975), .A2(new_n998), .A3(new_n1003), .A4(new_n1052), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n967), .A2(new_n968), .A3(G286), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT63), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1053), .A2(new_n1056), .ZN(new_n1057));
  XOR2_X1   g632(.A(KEYINPUT111), .B(G1971), .Z(new_n1058));
  AOI21_X1  g633(.A(new_n1058), .B1(new_n980), .B2(new_n985), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n990), .A2(G2090), .ZN(new_n1060));
  OAI21_X1  g635(.A(G8), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(G303), .A2(G8), .ZN(new_n1062));
  XOR2_X1   g637(.A(new_n1062), .B(KEYINPUT55), .Z(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1061), .A2(new_n1064), .ZN(new_n1065));
  OR2_X1    g640(.A1(G305), .A2(G1981), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT113), .ZN(new_n1067));
  XOR2_X1   g642(.A(KEYINPUT112), .B(G86), .Z(new_n1068));
  NAND2_X1  g643(.A1(new_n528), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1067), .B1(new_n1069), .B2(new_n591), .ZN(new_n1070));
  AOI211_X1 g645(.A(KEYINPUT113), .B(new_n590), .C1(new_n528), .C2(new_n1068), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n592), .A2(new_n531), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G1981), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1066), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT49), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1021), .A2(new_n968), .ZN(new_n1078));
  OAI211_X1 g653(.A(KEYINPUT49), .B(new_n1066), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G1976), .ZN(new_n1081));
  NOR2_X1   g656(.A1(G288), .A2(new_n1081), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1021), .A2(new_n968), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT52), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1083), .B(new_n1084), .C1(G1976), .C2(new_n695), .ZN(new_n1085));
  OR2_X1    g660(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1080), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1015), .A2(G2090), .ZN(new_n1088));
  OR3_X1    g663(.A1(new_n1059), .A2(KEYINPUT115), .A3(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT115), .B1(new_n1059), .B2(new_n1088), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1089), .A2(new_n1090), .A3(G8), .ZN(new_n1091));
  AOI211_X1 g666(.A(new_n1065), .B(new_n1087), .C1(new_n1091), .C2(new_n1064), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1057), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1061), .A2(new_n1064), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1087), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n1054), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1096), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT63), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1065), .B1(new_n1095), .B2(KEYINPUT63), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1080), .A2(new_n1081), .A3(new_n695), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n1066), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n1078), .B(KEYINPUT114), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1100), .A2(new_n1101), .A3(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1093), .A2(KEYINPUT123), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT123), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1091), .A2(new_n1064), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1109), .B(new_n1095), .C1(new_n1064), .C2(new_n1061), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1110), .B1(new_n1053), .B2(new_n1056), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1100), .A2(new_n1101), .A3(new_n1105), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1108), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT124), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT62), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n973), .A2(new_n1115), .A3(new_n974), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n997), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1114), .B1(new_n1117), .B2(new_n1110), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n975), .A2(KEYINPUT62), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1092), .A2(KEYINPUT124), .A3(new_n997), .A4(new_n1116), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1107), .A2(new_n1113), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n940), .B1(G1986), .B2(G290), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(G1986), .B2(G290), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n921), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n1122), .A2(KEYINPUT125), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT125), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n945), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT127), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT127), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1130), .B(new_n945), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(new_n1131), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g707(.A1(new_n841), .A2(G401), .A3(G227), .ZN(new_n1134));
  INV_X1    g708(.A(G229), .ZN(new_n1135));
  NAND4_X1  g709(.A1(new_n1134), .A2(G319), .A3(new_n1135), .A4(new_n907), .ZN(G225));
  INV_X1    g710(.A(G225), .ZN(G308));
endmodule


