//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 0 1 1 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n806,
    new_n807, new_n808, new_n809, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n878, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT24), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G183gat), .ZN(new_n205));
  INV_X1    g004(.A(G190gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND3_X1  g006(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n208));
  AND3_X1   g007(.A1(new_n204), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210));
  INV_X1    g009(.A(G169gat), .ZN(new_n211));
  INV_X1    g010(.A(G176gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT23), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n210), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(KEYINPUT23), .B1(new_n211), .B2(new_n212), .ZN(new_n216));
  NOR4_X1   g015(.A1(new_n209), .A2(new_n215), .A3(KEYINPUT25), .A4(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT66), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n207), .B(new_n208), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n204), .A2(KEYINPUT65), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n218), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NOR3_X1   g022(.A1(new_n214), .A2(G169gat), .A3(G176gat), .ZN(new_n224));
  INV_X1    g023(.A(new_n210), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT64), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT64), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n227), .B(new_n210), .C1(new_n213), .C2(new_n214), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(G183gat), .A2(G190gat), .ZN(new_n230));
  AND2_X1   g029(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n230), .B1(new_n231), .B2(G190gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n204), .A2(KEYINPUT65), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n219), .A2(new_n220), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n232), .A2(new_n233), .A3(KEYINPUT66), .A4(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n216), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n223), .A2(new_n229), .A3(new_n235), .A4(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n217), .B1(new_n237), .B2(KEYINPUT25), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n239));
  AND3_X1   g038(.A1(new_n239), .A2(KEYINPUT68), .A3(new_n210), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT68), .B1(new_n239), .B2(new_n210), .ZN(new_n241));
  NOR3_X1   g040(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n242));
  NOR3_X1   g041(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n202), .ZN(new_n244));
  OAI21_X1  g043(.A(KEYINPUT69), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n241), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n239), .A2(KEYINPUT68), .A3(new_n210), .ZN(new_n247));
  INV_X1    g046(.A(new_n242), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n249), .A2(new_n250), .A3(new_n202), .ZN(new_n251));
  XNOR2_X1  g050(.A(KEYINPUT27), .B(G183gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(new_n206), .ZN(new_n253));
  XOR2_X1   g052(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n245), .A2(new_n251), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n238), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT29), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(G226gat), .A2(G233gat), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n259), .A2(KEYINPUT75), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT75), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT29), .B1(new_n238), .B2(new_n256), .ZN(new_n263));
  INV_X1    g062(.A(new_n260), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n261), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G197gat), .B(G204gat), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT22), .ZN(new_n268));
  INV_X1    g067(.A(G211gat), .ZN(new_n269));
  INV_X1    g068(.A(G218gat), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G211gat), .B(G218gat), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n273), .A2(new_n267), .A3(new_n271), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  XOR2_X1   g077(.A(new_n260), .B(KEYINPUT73), .Z(new_n279));
  AOI21_X1  g078(.A(new_n278), .B1(new_n257), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n266), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT74), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n260), .B1(new_n238), .B2(new_n256), .ZN(new_n283));
  OAI22_X1  g082(.A1(new_n282), .A2(new_n283), .B1(new_n263), .B2(new_n279), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n282), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n278), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G8gat), .B(G36gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n288), .B(G92gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT76), .B(G64gat), .ZN(new_n290));
  XOR2_X1   g089(.A(new_n289), .B(new_n290), .Z(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  AND2_X1   g091(.A1(new_n292), .A2(KEYINPUT30), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n281), .A2(new_n287), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(G155gat), .A2(G162gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT80), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n295), .B1(new_n296), .B2(KEYINPUT2), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT2), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n298), .A2(KEYINPUT80), .ZN(new_n299));
  INV_X1    g098(.A(G141gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n300), .A2(G148gat), .ZN(new_n301));
  INV_X1    g100(.A(G148gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n302), .A2(G141gat), .ZN(new_n303));
  OAI22_X1  g102(.A1(new_n297), .A2(new_n299), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  NOR2_X1   g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n295), .B1(new_n305), .B2(KEYINPUT79), .ZN(new_n306));
  INV_X1    g105(.A(G155gat), .ZN(new_n307));
  INV_X1    g106(.A(G162gat), .ZN(new_n308));
  OR3_X1    g107(.A1(new_n307), .A2(new_n308), .A3(KEYINPUT79), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n304), .A2(new_n306), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n298), .A2(new_n307), .A3(new_n308), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(new_n295), .ZN(new_n312));
  OR2_X1    g111(.A1(KEYINPUT81), .A2(G141gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(KEYINPUT81), .A2(G141gat), .ZN(new_n314));
  AND3_X1   g113(.A1(new_n313), .A2(G148gat), .A3(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(KEYINPUT82), .B1(new_n300), .B2(G148gat), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT82), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n317), .A2(new_n302), .A3(G141gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n312), .B1(new_n315), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n310), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT1), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n322), .B1(G113gat), .B2(G120gat), .ZN(new_n323));
  AND2_X1   g122(.A1(G113gat), .A2(G120gat), .ZN(new_n324));
  OAI21_X1  g123(.A(KEYINPUT70), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G127gat), .B(G134gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n325), .B(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT4), .B1(new_n321), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT83), .ZN(new_n329));
  XOR2_X1   g128(.A(G127gat), .B(G134gat), .Z(new_n330));
  XNOR2_X1  g129(.A(new_n325), .B(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT4), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n331), .A2(new_n332), .A3(new_n320), .A4(new_n310), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n328), .A2(new_n329), .A3(new_n333), .ZN(new_n334));
  AND2_X1   g133(.A1(new_n309), .A2(new_n306), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n313), .A2(new_n314), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n316), .B(new_n318), .C1(new_n336), .C2(new_n302), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n304), .A2(new_n335), .B1(new_n337), .B2(new_n312), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(new_n331), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n339), .A2(KEYINPUT83), .A3(KEYINPUT4), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n321), .A2(KEYINPUT3), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n310), .A2(new_n320), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n341), .A2(new_n327), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(G225gat), .A2(G233gat), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n334), .A2(new_n340), .A3(new_n344), .A4(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT85), .B(KEYINPUT5), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n321), .A2(new_n327), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n339), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n345), .ZN(new_n350));
  AND3_X1   g149(.A1(new_n349), .A2(KEYINPUT84), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT84), .B1(new_n349), .B2(new_n350), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n346), .B(new_n347), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n328), .A2(new_n333), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n347), .A2(new_n350), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n354), .A2(new_n344), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT87), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT87), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n354), .A2(new_n344), .A3(new_n358), .A4(new_n355), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n353), .A2(new_n360), .ZN(new_n361));
  XOR2_X1   g160(.A(G57gat), .B(G85gat), .Z(new_n362));
  XNOR2_X1  g161(.A(G1gat), .B(G29gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n362), .B(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(KEYINPUT86), .B(KEYINPUT0), .ZN(new_n365));
  XOR2_X1   g164(.A(new_n364), .B(new_n365), .Z(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n361), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT6), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n360), .A3(new_n366), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n361), .A2(KEYINPUT6), .A3(new_n367), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n294), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT77), .ZN(new_n374));
  INV_X1    g173(.A(new_n279), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n259), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n257), .A2(new_n264), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT74), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n376), .A2(new_n378), .A3(new_n285), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n278), .A2(new_n379), .B1(new_n266), .B2(new_n280), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n374), .B1(new_n380), .B2(new_n292), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n281), .A2(new_n287), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n382), .A2(KEYINPUT77), .A3(new_n291), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n380), .A2(new_n292), .ZN(new_n385));
  XNOR2_X1  g184(.A(KEYINPUT78), .B(KEYINPUT30), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n373), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n257), .A2(new_n331), .ZN(new_n389));
  INV_X1    g188(.A(G227gat), .ZN(new_n390));
  INV_X1    g189(.A(G233gat), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n238), .A2(new_n256), .A3(new_n327), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n389), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT32), .ZN(new_n395));
  XOR2_X1   g194(.A(KEYINPUT71), .B(KEYINPUT33), .Z(new_n396));
  NAND2_X1  g195(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  XOR2_X1   g196(.A(G71gat), .B(G99gat), .Z(new_n398));
  XNOR2_X1  g197(.A(G15gat), .B(G43gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n395), .A2(new_n397), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT72), .ZN(new_n402));
  OR2_X1    g201(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n400), .A2(new_n402), .ZN(new_n404));
  INV_X1    g203(.A(new_n396), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n394), .A2(KEYINPUT32), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n401), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT34), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n389), .A2(new_n393), .ZN(new_n410));
  INV_X1    g209(.A(new_n392), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n410), .A2(new_n409), .A3(new_n411), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n408), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n414), .A2(new_n412), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n416), .A2(new_n407), .A3(new_n401), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT88), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT29), .B1(new_n275), .B2(new_n276), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n321), .B1(new_n419), .B2(KEYINPUT3), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n277), .B1(new_n343), .B2(new_n258), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n418), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT29), .B1(new_n338), .B2(new_n342), .ZN(new_n424));
  OAI211_X1 g223(.A(KEYINPUT88), .B(new_n420), .C1(new_n424), .C2(new_n277), .ZN(new_n425));
  NAND2_X1  g224(.A1(G228gat), .A2(G233gat), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n423), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n426), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n418), .B(new_n428), .C1(new_n421), .C2(new_n422), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(G22gat), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n427), .A2(G22gat), .A3(new_n429), .ZN(new_n433));
  XNOR2_X1  g232(.A(G78gat), .B(G106gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(KEYINPUT31), .B(G50gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n434), .B(new_n435), .ZN(new_n436));
  AND4_X1   g235(.A1(KEYINPUT89), .A2(new_n432), .A3(new_n433), .A4(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT89), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n433), .A2(new_n438), .ZN(new_n439));
  AOI22_X1  g238(.A1(new_n439), .A2(new_n436), .B1(new_n432), .B2(new_n433), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n415), .B(new_n417), .C1(new_n437), .C2(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT35), .B1(new_n388), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT91), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT91), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n444), .B(KEYINPUT35), .C1(new_n388), .C2(new_n441), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT90), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT35), .B1(new_n371), .B2(new_n372), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n294), .B1(new_n385), .B2(new_n386), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(new_n448), .A3(new_n384), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n446), .B1(new_n449), .B2(new_n441), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n384), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n441), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n452), .A2(new_n453), .A3(KEYINPUT90), .A4(new_n447), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n443), .A2(new_n445), .A3(new_n450), .A4(new_n454), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n380), .A2(KEYINPUT37), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n281), .A2(KEYINPUT37), .A3(new_n287), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n291), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT38), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n371), .A2(new_n372), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n292), .A2(KEYINPUT38), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT37), .B1(new_n379), .B2(new_n278), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n257), .A2(new_n279), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n277), .B1(new_n266), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n462), .B1(new_n456), .B2(new_n466), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n459), .A2(new_n461), .A3(new_n385), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n354), .A2(new_n344), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n350), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n470), .A2(KEYINPUT39), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n471), .A2(new_n367), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n470), .B(KEYINPUT39), .C1(new_n350), .C2(new_n349), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n368), .B1(new_n474), .B2(KEYINPUT40), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n475), .B1(KEYINPUT40), .B2(new_n474), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n451), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n437), .A2(new_n440), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n468), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n415), .A2(new_n417), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT36), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT36), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n483), .A2(new_n485), .B1(new_n388), .B2(new_n478), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n480), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n455), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(G229gat), .A2(G233gat), .ZN(new_n489));
  XOR2_X1   g288(.A(new_n489), .B(KEYINPUT95), .Z(new_n490));
  XOR2_X1   g289(.A(new_n490), .B(KEYINPUT13), .Z(new_n491));
  INV_X1    g290(.A(G29gat), .ZN(new_n492));
  INV_X1    g291(.A(G36gat), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n492), .A2(new_n493), .A3(KEYINPUT14), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT14), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n495), .B1(G29gat), .B2(G36gat), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n494), .B(new_n496), .C1(new_n492), .C2(new_n493), .ZN(new_n497));
  INV_X1    g296(.A(G50gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(G43gat), .ZN(new_n499));
  INV_X1    g298(.A(G43gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(G50gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT92), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT15), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  OR3_X1    g303(.A1(new_n497), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n502), .B1(new_n497), .B2(new_n504), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT15), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n497), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n505), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT93), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT93), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n505), .A2(new_n506), .A3(new_n511), .A4(new_n508), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(G8gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(G15gat), .B(G22gat), .ZN(new_n515));
  OR2_X1    g314(.A1(new_n515), .A2(G1gat), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT94), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT16), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n515), .B1(new_n519), .B2(G1gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n518), .B(new_n521), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n513), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n513), .A2(new_n522), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n491), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n513), .A2(new_n522), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT17), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n510), .A2(new_n527), .A3(new_n512), .ZN(new_n528));
  INV_X1    g327(.A(new_n522), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n509), .A2(KEYINPUT17), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n526), .A2(new_n531), .A3(KEYINPUT18), .A4(new_n490), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n525), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n526), .A2(new_n531), .A3(new_n490), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT18), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT96), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G113gat), .B(G141gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(KEYINPUT11), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(new_n211), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n541), .A2(G197gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(G197gat), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n542), .A2(KEYINPUT12), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT12), .B1(new_n542), .B2(new_n543), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n534), .A2(KEYINPUT96), .A3(new_n535), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n533), .A2(new_n538), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n536), .A2(new_n532), .A3(new_n525), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n549), .B1(new_n545), .B2(new_n544), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G190gat), .B(G218gat), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  AND3_X1   g352(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(KEYINPUT99), .B(KEYINPUT7), .ZN(new_n555));
  NAND2_X1  g354(.A1(G85gat), .A2(G92gat), .ZN(new_n556));
  OR2_X1    g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n556), .ZN(new_n558));
  NAND2_X1  g357(.A1(G99gat), .A2(G106gat), .ZN(new_n559));
  INV_X1    g358(.A(G85gat), .ZN(new_n560));
  INV_X1    g359(.A(G92gat), .ZN(new_n561));
  AOI22_X1  g360(.A1(KEYINPUT8), .A2(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n557), .A2(new_n558), .A3(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G99gat), .B(G106gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT100), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n563), .B(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n554), .B1(new_n513), .B2(new_n566), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n563), .A2(new_n565), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n563), .A2(new_n565), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n528), .A2(new_n530), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n553), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n571), .A2(KEYINPUT102), .ZN(new_n572));
  XOR2_X1   g371(.A(G134gat), .B(G162gat), .Z(new_n573));
  AOI21_X1  g372(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  AND3_X1   g374(.A1(new_n567), .A2(new_n553), .A3(new_n570), .ZN(new_n576));
  NOR3_X1   g375(.A1(new_n572), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n571), .A2(KEYINPUT102), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n575), .B1(new_n576), .B2(new_n571), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(KEYINPUT101), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT101), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n582), .B(new_n575), .C1(new_n576), .C2(new_n571), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT9), .ZN(new_n586));
  INV_X1    g385(.A(G71gat), .ZN(new_n587));
  INV_X1    g386(.A(G78gat), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT97), .ZN(new_n590));
  XOR2_X1   g389(.A(G57gat), .B(G64gat), .Z(new_n591));
  INV_X1    g390(.A(KEYINPUT97), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n592), .B(new_n586), .C1(new_n587), .C2(new_n588), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n590), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G71gat), .B(G78gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n522), .B1(KEYINPUT21), .B2(new_n596), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n596), .A2(KEYINPUT21), .ZN(new_n598));
  XNOR2_X1  g397(.A(G127gat), .B(G155gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(G211gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n602));
  NAND2_X1  g401(.A1(G231gat), .A2(G233gat), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n602), .B(new_n603), .Z(new_n604));
  OR2_X1    g403(.A1(new_n598), .A2(new_n599), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n598), .A2(new_n599), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n605), .A2(new_n269), .A3(new_n606), .ZN(new_n607));
  AND3_X1   g406(.A1(new_n601), .A2(new_n604), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n604), .B1(new_n601), .B2(new_n607), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n597), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(KEYINPUT98), .B(G183gat), .ZN(new_n611));
  INV_X1    g410(.A(new_n604), .ZN(new_n612));
  INV_X1    g411(.A(new_n607), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n269), .B1(new_n605), .B2(new_n606), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n597), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n601), .A2(new_n604), .A3(new_n607), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  AND3_X1   g417(.A1(new_n610), .A2(new_n611), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n611), .B1(new_n610), .B2(new_n618), .ZN(new_n620));
  NOR3_X1   g419(.A1(new_n585), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n566), .A2(new_n596), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n594), .B(new_n595), .Z(new_n623));
  NAND3_X1  g422(.A1(new_n623), .A2(new_n568), .A3(new_n569), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT10), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n622), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n566), .A2(KEYINPUT10), .A3(new_n596), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(G230gat), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n629), .A2(new_n391), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n622), .A2(new_n624), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(new_n630), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G120gat), .B(G148gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(G176gat), .ZN(new_n637));
  INV_X1    g436(.A(G204gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n635), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n632), .A2(new_n634), .A3(new_n639), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  AND4_X1   g443(.A1(new_n488), .A2(new_n551), .A3(new_n621), .A4(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(new_n461), .ZN(new_n646));
  XOR2_X1   g445(.A(KEYINPUT103), .B(G1gat), .Z(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(G1324gat));
  AND2_X1   g447(.A1(new_n645), .A2(new_n451), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n649), .A2(new_n514), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT42), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT104), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(new_n514), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n645), .A2(new_n451), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n650), .B1(new_n651), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n655), .B1(new_n651), .B2(new_n654), .ZN(G1325gat));
  INV_X1    g455(.A(G15gat), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n645), .A2(new_n657), .A3(new_n482), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n483), .A2(new_n485), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n645), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n658), .B1(new_n661), .B2(new_n657), .ZN(G1326gat));
  NAND2_X1  g461(.A1(new_n645), .A2(new_n478), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT43), .B(G22gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(G1327gat));
  INV_X1    g464(.A(new_n585), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n666), .B1(new_n455), .B2(new_n487), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n619), .A2(new_n620), .ZN(new_n668));
  INV_X1    g467(.A(new_n551), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n668), .A2(new_n669), .A3(new_n643), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n672), .A2(new_n492), .A3(new_n461), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT45), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n667), .B(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(new_n670), .ZN(new_n677));
  OAI21_X1  g476(.A(G29gat), .B1(new_n677), .B2(new_n460), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n674), .A2(new_n678), .ZN(G1328gat));
  NOR3_X1   g478(.A1(new_n671), .A2(G36gat), .A3(new_n452), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT46), .ZN(new_n681));
  OAI21_X1  g480(.A(G36gat), .B1(new_n677), .B2(new_n452), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(G1329gat));
  NAND3_X1  g482(.A1(new_n672), .A2(new_n500), .A3(new_n482), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n684), .A2(KEYINPUT47), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n675), .B1(new_n488), .B2(new_n585), .ZN(new_n686));
  AOI211_X1 g485(.A(KEYINPUT44), .B(new_n666), .C1(new_n455), .C2(new_n487), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n660), .B(new_n670), .C1(new_n686), .C2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(KEYINPUT106), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(G43gat), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n688), .A2(KEYINPUT106), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n685), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n688), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n684), .B1(new_n693), .B2(new_n500), .ZN(new_n694));
  XNOR2_X1  g493(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n692), .A2(new_n696), .ZN(G1330gat));
  NAND2_X1  g496(.A1(new_n672), .A2(KEYINPUT107), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT107), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n671), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n698), .A2(new_n498), .A3(new_n478), .A4(new_n700), .ZN(new_n701));
  OAI211_X1 g500(.A(new_n478), .B(new_n670), .C1(new_n686), .C2(new_n687), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(G50gat), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT48), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n701), .A2(new_n703), .A3(KEYINPUT48), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(G1331gat));
  NAND3_X1  g507(.A1(new_n621), .A2(new_n669), .A3(new_n643), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n709), .B1(new_n455), .B2(new_n487), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n461), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g511(.A(new_n452), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT108), .ZN(new_n715));
  NOR2_X1   g514(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1333gat));
  NOR2_X1   g516(.A1(new_n659), .A2(new_n587), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n710), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT109), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n710), .A2(new_n482), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n587), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n478), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g526(.A1(new_n668), .A2(new_n551), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n643), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT110), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n676), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n560), .B1(new_n731), .B2(new_n461), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n667), .A2(new_n728), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT51), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n667), .A2(KEYINPUT51), .A3(new_n728), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AND4_X1   g536(.A1(new_n560), .A2(new_n737), .A3(new_n461), .A4(new_n643), .ZN(new_n738));
  OR2_X1    g537(.A1(new_n732), .A2(new_n738), .ZN(G1336gat));
  NAND3_X1  g538(.A1(new_n676), .A2(new_n451), .A3(new_n730), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(G92gat), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n737), .A2(new_n561), .A3(new_n451), .A4(new_n643), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT52), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  AND4_X1   g543(.A1(KEYINPUT51), .A2(new_n488), .A3(new_n585), .A4(new_n728), .ZN(new_n745));
  XOR2_X1   g544(.A(KEYINPUT111), .B(KEYINPUT51), .Z(new_n746));
  AOI21_X1  g545(.A(new_n746), .B1(new_n667), .B2(new_n728), .ZN(new_n747));
  OR2_X1    g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n452), .A2(G92gat), .A3(new_n644), .ZN(new_n749));
  AOI22_X1  g548(.A1(new_n740), .A2(G92gat), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n744), .B1(new_n743), .B2(new_n750), .ZN(G1337gat));
  INV_X1    g550(.A(G99gat), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n737), .A2(new_n482), .A3(new_n643), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n659), .A2(new_n752), .ZN(new_n754));
  AOI22_X1  g553(.A1(new_n752), .A2(new_n753), .B1(new_n731), .B2(new_n754), .ZN(G1338gat));
  NOR3_X1   g554(.A1(new_n479), .A2(G106gat), .A3(new_n644), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n756), .B1(new_n745), .B2(new_n747), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT112), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI211_X1 g558(.A(KEYINPUT112), .B(new_n756), .C1(new_n745), .C2(new_n747), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n478), .B(new_n730), .C1(new_n686), .C2(new_n687), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G106gat), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n759), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT53), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT113), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n676), .A2(new_n765), .A3(new_n478), .A4(new_n730), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n761), .A2(KEYINPUT113), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n766), .A2(new_n767), .A3(G106gat), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT53), .B1(new_n737), .B2(new_n756), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n764), .A2(new_n770), .ZN(G1339gat));
  INV_X1    g570(.A(new_n668), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n626), .A2(new_n627), .A3(new_n630), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n632), .A2(KEYINPUT54), .A3(new_n773), .ZN(new_n774));
  XOR2_X1   g573(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n775));
  NAND3_X1  g574(.A1(new_n628), .A2(new_n631), .A3(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT115), .ZN(new_n777));
  AND3_X1   g576(.A1(new_n776), .A2(new_n777), .A3(new_n640), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n777), .B1(new_n776), .B2(new_n640), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n774), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI211_X1 g581(.A(KEYINPUT55), .B(new_n774), .C1(new_n778), .C2(new_n779), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n782), .A2(new_n551), .A3(new_n642), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n542), .A2(new_n543), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n523), .A2(new_n524), .A3(new_n491), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n490), .B1(new_n526), .B2(new_n531), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n785), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n548), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n643), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n585), .B1(new_n784), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n585), .A2(new_n782), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n783), .A2(new_n548), .A3(new_n642), .A4(new_n788), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n772), .B1(new_n791), .B2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n621), .A2(new_n669), .A3(new_n644), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n451), .A2(new_n460), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n797), .A2(new_n453), .A3(new_n798), .ZN(new_n799));
  XOR2_X1   g598(.A(new_n799), .B(KEYINPUT117), .Z(new_n800));
  INV_X1    g599(.A(G113gat), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n800), .A2(new_n801), .A3(new_n551), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n799), .B(KEYINPUT116), .ZN(new_n803));
  OAI21_X1  g602(.A(G113gat), .B1(new_n803), .B2(new_n669), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(G1340gat));
  NOR2_X1   g604(.A1(new_n644), .A2(G120gat), .ZN(new_n806));
  XOR2_X1   g605(.A(new_n806), .B(KEYINPUT118), .Z(new_n807));
  NAND2_X1  g606(.A1(new_n800), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(G120gat), .B1(new_n803), .B2(new_n644), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(G1341gat));
  OAI21_X1  g609(.A(G127gat), .B1(new_n803), .B2(new_n772), .ZN(new_n811));
  OR3_X1    g610(.A1(new_n799), .A2(G127gat), .A3(new_n772), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT119), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT119), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n811), .A2(new_n815), .A3(new_n812), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(G1342gat));
  AND2_X1   g616(.A1(KEYINPUT120), .A2(KEYINPUT56), .ZN(new_n818));
  NOR2_X1   g617(.A1(KEYINPUT120), .A2(KEYINPUT56), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n799), .A2(G134gat), .A3(new_n666), .ZN(new_n821));
  MUX2_X1   g620(.A(new_n820), .B(new_n818), .S(new_n821), .Z(new_n822));
  OAI21_X1  g621(.A(G134gat), .B1(new_n803), .B2(new_n666), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(G1343gat));
  INV_X1    g623(.A(KEYINPUT57), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n797), .A2(new_n825), .A3(new_n478), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n659), .A2(new_n798), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g628(.A(KEYINPUT121), .B(KEYINPUT57), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  AND4_X1   g630(.A1(new_n669), .A2(new_n668), .A3(new_n666), .A4(new_n644), .ZN(new_n832));
  AOI22_X1  g631(.A1(new_n780), .A2(new_n781), .B1(new_n548), .B2(new_n550), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n783), .A2(new_n642), .ZN(new_n834));
  AOI22_X1  g633(.A1(new_n833), .A2(new_n834), .B1(new_n643), .B2(new_n789), .ZN(new_n835));
  OAI22_X1  g634(.A1(new_n835), .A2(new_n585), .B1(new_n792), .B2(new_n793), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n832), .B1(new_n836), .B2(new_n772), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n831), .B1(new_n837), .B2(new_n479), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n829), .A2(new_n551), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n336), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n797), .A2(new_n478), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(new_n827), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n842), .A2(new_n300), .A3(new_n551), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(KEYINPUT58), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT58), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n840), .A2(new_n846), .A3(new_n843), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(new_n847), .ZN(G1344gat));
  NAND3_X1  g647(.A1(new_n842), .A2(new_n302), .A3(new_n643), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT57), .B1(new_n797), .B2(new_n478), .ZN(new_n851));
  AOI211_X1 g650(.A(new_n479), .B(new_n830), .C1(new_n795), .C2(new_n796), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n643), .B(new_n828), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n850), .B1(new_n853), .B2(G148gat), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n838), .A2(new_n643), .A3(new_n826), .A4(new_n828), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n302), .A2(KEYINPUT59), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n849), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT122), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT122), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n860), .B(new_n849), .C1(new_n854), .C2(new_n857), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(G1345gat));
  NAND3_X1  g661(.A1(new_n829), .A2(new_n668), .A3(new_n838), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(G155gat), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n842), .A2(new_n307), .A3(new_n668), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(KEYINPUT123), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT123), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n864), .A2(new_n868), .A3(new_n865), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n869), .ZN(G1346gat));
  NAND3_X1  g669(.A1(new_n842), .A2(new_n308), .A3(new_n585), .ZN(new_n871));
  AND3_X1   g670(.A1(new_n829), .A2(new_n585), .A3(new_n838), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n871), .B1(new_n872), .B2(new_n308), .ZN(G1347gat));
  NOR2_X1   g672(.A1(new_n452), .A2(new_n461), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n797), .A2(new_n453), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n551), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n876), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n643), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n878), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g678(.A1(new_n875), .A2(new_n668), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n205), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n881), .B1(new_n252), .B2(new_n880), .ZN(new_n882));
  XOR2_X1   g681(.A(new_n882), .B(KEYINPUT60), .Z(G1350gat));
  AOI21_X1  g682(.A(new_n206), .B1(new_n875), .B2(new_n585), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT61), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(KEYINPUT124), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n885), .A2(KEYINPUT124), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n884), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n875), .A2(new_n206), .A3(new_n585), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n887), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT125), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n887), .A2(KEYINPUT125), .A3(new_n889), .A4(new_n890), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(G1351gat));
  NAND2_X1  g694(.A1(new_n874), .A2(new_n659), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n841), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(G197gat), .B1(new_n897), .B2(new_n551), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n851), .A2(new_n852), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n899), .A2(new_n896), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n551), .A2(G197gat), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(G1352gat));
  NAND3_X1  g701(.A1(new_n897), .A2(new_n638), .A3(new_n643), .ZN(new_n903));
  XOR2_X1   g702(.A(new_n903), .B(KEYINPUT62), .Z(new_n904));
  NOR3_X1   g703(.A1(new_n899), .A2(new_n644), .A3(new_n896), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n638), .B2(new_n905), .ZN(G1353gat));
  NAND3_X1  g705(.A1(new_n897), .A2(new_n269), .A3(new_n668), .ZN(new_n907));
  INV_X1    g706(.A(new_n896), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n668), .B(new_n908), .C1(new_n851), .C2(new_n852), .ZN(new_n909));
  OR2_X1    g708(.A1(new_n909), .A2(KEYINPUT126), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n269), .B1(new_n909), .B2(KEYINPUT126), .ZN(new_n911));
  AND3_X1   g710(.A1(new_n910), .A2(KEYINPUT63), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(KEYINPUT63), .B1(new_n910), .B2(new_n911), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n907), .B1(new_n912), .B2(new_n913), .ZN(G1354gat));
  AOI21_X1  g713(.A(G218gat), .B1(new_n897), .B2(new_n585), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n915), .A2(KEYINPUT127), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(KEYINPUT127), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n666), .A2(new_n270), .ZN(new_n918));
  AOI22_X1  g717(.A1(new_n916), .A2(new_n917), .B1(new_n900), .B2(new_n918), .ZN(G1355gat));
endmodule


