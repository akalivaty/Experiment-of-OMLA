

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U547 ( .A1(n965), .A2(n673), .ZN(n640) );
  INV_X1 U548 ( .A(KEYINPUT103), .ZN(n702) );
  BUF_X1 U549 ( .A(n652), .Z(n689) );
  XNOR2_X1 U550 ( .A(n698), .B(KEYINPUT32), .ZN(n699) );
  NOR2_X1 U551 ( .A1(G164), .A2(G1384), .ZN(n614) );
  XNOR2_X1 U552 ( .A(KEYINPUT78), .B(KEYINPUT13), .ZN(n646) );
  XNOR2_X1 U553 ( .A(n647), .B(n646), .ZN(n648) );
  NOR2_X2 U554 ( .A1(G2105), .A2(n516), .ZN(n858) );
  NOR2_X1 U555 ( .A1(n554), .A2(n529), .ZN(n771) );
  NOR2_X1 U556 ( .A1(G651), .A2(n554), .ZN(n779) );
  NAND2_X1 U557 ( .A1(n651), .A2(n650), .ZN(n975) );
  NOR2_X1 U558 ( .A1(G2104), .A2(G2105), .ZN(n512) );
  XOR2_X2 U559 ( .A(KEYINPUT17), .B(n512), .Z(n861) );
  NAND2_X1 U560 ( .A1(G138), .A2(n861), .ZN(n513) );
  XNOR2_X1 U561 ( .A(n513), .B(KEYINPUT92), .ZN(n522) );
  XNOR2_X1 U562 ( .A(KEYINPUT65), .B(G2104), .ZN(n516) );
  NAND2_X1 U563 ( .A1(G102), .A2(n858), .ZN(n514) );
  XNOR2_X1 U564 ( .A(KEYINPUT91), .B(n514), .ZN(n520) );
  AND2_X1 U565 ( .A1(G2104), .A2(G2105), .ZN(n852) );
  NAND2_X1 U566 ( .A1(n852), .A2(G114), .ZN(n515) );
  XNOR2_X1 U567 ( .A(n515), .B(KEYINPUT90), .ZN(n518) );
  AND2_X1 U568 ( .A1(n516), .A2(G2105), .ZN(n854) );
  NAND2_X1 U569 ( .A1(G126), .A2(n854), .ZN(n517) );
  NAND2_X1 U570 ( .A1(n518), .A2(n517), .ZN(n519) );
  NOR2_X1 U571 ( .A1(n520), .A2(n519), .ZN(n521) );
  AND2_X1 U572 ( .A1(n522), .A2(n521), .ZN(G164) );
  NOR2_X1 U573 ( .A1(G543), .A2(G651), .ZN(n523) );
  XNOR2_X1 U574 ( .A(n523), .B(KEYINPUT64), .ZN(n775) );
  NAND2_X1 U575 ( .A1(n775), .A2(G89), .ZN(n524) );
  XOR2_X1 U576 ( .A(KEYINPUT79), .B(n524), .Z(n525) );
  XNOR2_X1 U577 ( .A(n525), .B(KEYINPUT4), .ZN(n527) );
  XOR2_X1 U578 ( .A(KEYINPUT0), .B(G543), .Z(n554) );
  INV_X1 U579 ( .A(G651), .ZN(n529) );
  NAND2_X1 U580 ( .A1(G76), .A2(n771), .ZN(n526) );
  NAND2_X1 U581 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U582 ( .A(n528), .B(KEYINPUT5), .ZN(n537) );
  NOR2_X1 U583 ( .A1(G543), .A2(n529), .ZN(n530) );
  XOR2_X1 U584 ( .A(KEYINPUT68), .B(n530), .Z(n531) );
  XNOR2_X1 U585 ( .A(KEYINPUT1), .B(n531), .ZN(n772) );
  NAND2_X1 U586 ( .A1(G63), .A2(n772), .ZN(n532) );
  XNOR2_X1 U587 ( .A(n532), .B(KEYINPUT80), .ZN(n534) );
  NAND2_X1 U588 ( .A1(G51), .A2(n779), .ZN(n533) );
  NAND2_X1 U589 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U590 ( .A(KEYINPUT6), .B(n535), .Z(n536) );
  NAND2_X1 U591 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U592 ( .A(n538), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U593 ( .A1(n771), .A2(G77), .ZN(n539) );
  XOR2_X1 U594 ( .A(KEYINPUT71), .B(n539), .Z(n541) );
  NAND2_X1 U595 ( .A1(G90), .A2(n775), .ZN(n540) );
  NAND2_X1 U596 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U597 ( .A(n542), .B(KEYINPUT9), .ZN(n544) );
  NAND2_X1 U598 ( .A1(G64), .A2(n772), .ZN(n543) );
  NAND2_X1 U599 ( .A1(n544), .A2(n543), .ZN(n547) );
  NAND2_X1 U600 ( .A1(n779), .A2(G52), .ZN(n545) );
  XOR2_X1 U601 ( .A(KEYINPUT70), .B(n545), .Z(n546) );
  NOR2_X1 U602 ( .A1(n547), .A2(n546), .ZN(G171) );
  INV_X1 U603 ( .A(G171), .ZN(G301) );
  XOR2_X1 U604 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U605 ( .A1(n771), .A2(G75), .ZN(n549) );
  NAND2_X1 U606 ( .A1(G88), .A2(n775), .ZN(n548) );
  NAND2_X1 U607 ( .A1(n549), .A2(n548), .ZN(n553) );
  NAND2_X1 U608 ( .A1(n779), .A2(G50), .ZN(n551) );
  NAND2_X1 U609 ( .A1(G62), .A2(n772), .ZN(n550) );
  NAND2_X1 U610 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U611 ( .A1(n553), .A2(n552), .ZN(G166) );
  INV_X1 U612 ( .A(G166), .ZN(G303) );
  NAND2_X1 U613 ( .A1(G87), .A2(n554), .ZN(n556) );
  NAND2_X1 U614 ( .A1(G74), .A2(G651), .ZN(n555) );
  NAND2_X1 U615 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U616 ( .A1(n772), .A2(n557), .ZN(n559) );
  NAND2_X1 U617 ( .A1(n779), .A2(G49), .ZN(n558) );
  NAND2_X1 U618 ( .A1(n559), .A2(n558), .ZN(G288) );
  XOR2_X1 U619 ( .A(KEYINPUT84), .B(KEYINPUT2), .Z(n561) );
  NAND2_X1 U620 ( .A1(G73), .A2(n771), .ZN(n560) );
  XNOR2_X1 U621 ( .A(n561), .B(n560), .ZN(n565) );
  NAND2_X1 U622 ( .A1(G61), .A2(n772), .ZN(n563) );
  NAND2_X1 U623 ( .A1(G86), .A2(n775), .ZN(n562) );
  NAND2_X1 U624 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U625 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U626 ( .A(KEYINPUT85), .B(n566), .Z(n568) );
  NAND2_X1 U627 ( .A1(n779), .A2(G48), .ZN(n567) );
  NAND2_X1 U628 ( .A1(n568), .A2(n567), .ZN(G305) );
  NAND2_X1 U629 ( .A1(n779), .A2(G47), .ZN(n570) );
  NAND2_X1 U630 ( .A1(G60), .A2(n772), .ZN(n569) );
  NAND2_X1 U631 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U632 ( .A(KEYINPUT69), .B(n571), .Z(n574) );
  NAND2_X1 U633 ( .A1(G85), .A2(n775), .ZN(n572) );
  XNOR2_X1 U634 ( .A(KEYINPUT67), .B(n572), .ZN(n573) );
  NOR2_X1 U635 ( .A1(n574), .A2(n573), .ZN(n576) );
  NAND2_X1 U636 ( .A1(n771), .A2(G72), .ZN(n575) );
  NAND2_X1 U637 ( .A1(n576), .A2(n575), .ZN(G290) );
  AND2_X1 U638 ( .A1(G125), .A2(n854), .ZN(n580) );
  NAND2_X1 U639 ( .A1(G137), .A2(n861), .ZN(n578) );
  NAND2_X1 U640 ( .A1(G113), .A2(n852), .ZN(n577) );
  NAND2_X1 U641 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U642 ( .A1(n580), .A2(n579), .ZN(n744) );
  AND2_X1 U643 ( .A1(G40), .A2(n744), .ZN(n584) );
  INV_X1 U644 ( .A(KEYINPUT66), .ZN(n582) );
  NAND2_X1 U645 ( .A1(G101), .A2(n858), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(n583), .B(KEYINPUT23), .ZN(n745) );
  NAND2_X1 U648 ( .A1(n584), .A2(n745), .ZN(n615) );
  NOR2_X1 U649 ( .A1(n614), .A2(n615), .ZN(n739) );
  NAND2_X1 U650 ( .A1(G116), .A2(n852), .ZN(n586) );
  NAND2_X1 U651 ( .A1(G128), .A2(n854), .ZN(n585) );
  NAND2_X1 U652 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n587), .B(KEYINPUT35), .ZN(n592) );
  NAND2_X1 U654 ( .A1(G140), .A2(n861), .ZN(n589) );
  NAND2_X1 U655 ( .A1(G104), .A2(n858), .ZN(n588) );
  NAND2_X1 U656 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U657 ( .A(KEYINPUT34), .B(n590), .Z(n591) );
  NAND2_X1 U658 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U659 ( .A(n593), .B(KEYINPUT36), .Z(n871) );
  XNOR2_X1 U660 ( .A(G2067), .B(KEYINPUT37), .ZN(n737) );
  OR2_X1 U661 ( .A1(n871), .A2(n737), .ZN(n594) );
  XNOR2_X1 U662 ( .A(n594), .B(KEYINPUT93), .ZN(n926) );
  NAND2_X1 U663 ( .A1(n739), .A2(n926), .ZN(n735) );
  NAND2_X1 U664 ( .A1(G107), .A2(n852), .ZN(n596) );
  NAND2_X1 U665 ( .A1(G119), .A2(n854), .ZN(n595) );
  NAND2_X1 U666 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U667 ( .A(KEYINPUT94), .B(n597), .Z(n601) );
  NAND2_X1 U668 ( .A1(G131), .A2(n861), .ZN(n599) );
  NAND2_X1 U669 ( .A1(G95), .A2(n858), .ZN(n598) );
  AND2_X1 U670 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U671 ( .A1(n601), .A2(n600), .ZN(n866) );
  XOR2_X1 U672 ( .A(KEYINPUT95), .B(G1991), .Z(n935) );
  AND2_X1 U673 ( .A1(n866), .A2(n935), .ZN(n611) );
  XOR2_X1 U674 ( .A(KEYINPUT38), .B(KEYINPUT96), .Z(n603) );
  NAND2_X1 U675 ( .A1(G105), .A2(n858), .ZN(n602) );
  XNOR2_X1 U676 ( .A(n603), .B(n602), .ZN(n607) );
  NAND2_X1 U677 ( .A1(G141), .A2(n861), .ZN(n605) );
  NAND2_X1 U678 ( .A1(G117), .A2(n852), .ZN(n604) );
  NAND2_X1 U679 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U680 ( .A1(n607), .A2(n606), .ZN(n609) );
  NAND2_X1 U681 ( .A1(n854), .A2(G129), .ZN(n608) );
  NAND2_X1 U682 ( .A1(n609), .A2(n608), .ZN(n870) );
  AND2_X1 U683 ( .A1(G1996), .A2(n870), .ZN(n610) );
  NOR2_X1 U684 ( .A1(n611), .A2(n610), .ZN(n915) );
  XNOR2_X1 U685 ( .A(KEYINPUT97), .B(n739), .ZN(n612) );
  NOR2_X1 U686 ( .A1(n915), .A2(n612), .ZN(n732) );
  INV_X1 U687 ( .A(n732), .ZN(n613) );
  NAND2_X1 U688 ( .A1(n735), .A2(n613), .ZN(n727) );
  INV_X1 U689 ( .A(n614), .ZN(n616) );
  NOR2_X2 U690 ( .A1(n616), .A2(n615), .ZN(n633) );
  INV_X1 U691 ( .A(n633), .ZN(n652) );
  NOR2_X1 U692 ( .A1(G2084), .A2(n689), .ZN(n617) );
  NAND2_X1 U693 ( .A1(G8), .A2(n617), .ZN(n687) );
  NAND2_X1 U694 ( .A1(G8), .A2(n652), .ZN(n721) );
  NOR2_X1 U695 ( .A1(G1966), .A2(n721), .ZN(n685) );
  NOR2_X1 U696 ( .A1(n685), .A2(n617), .ZN(n618) );
  NAND2_X1 U697 ( .A1(G8), .A2(n618), .ZN(n619) );
  XNOR2_X1 U698 ( .A(n619), .B(KEYINPUT30), .ZN(n620) );
  NOR2_X1 U699 ( .A1(n620), .A2(G168), .ZN(n621) );
  XNOR2_X1 U700 ( .A(n621), .B(KEYINPUT99), .ZN(n625) );
  XOR2_X1 U701 ( .A(G2078), .B(KEYINPUT25), .Z(n936) );
  NOR2_X1 U702 ( .A1(n936), .A2(n689), .ZN(n623) );
  INV_X1 U703 ( .A(n689), .ZN(n665) );
  NOR2_X1 U704 ( .A1(n665), .A2(G1961), .ZN(n622) );
  NOR2_X1 U705 ( .A1(n623), .A2(n622), .ZN(n679) );
  NAND2_X1 U706 ( .A1(n679), .A2(G301), .ZN(n624) );
  NAND2_X1 U707 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U708 ( .A(n626), .B(KEYINPUT31), .ZN(n683) );
  NAND2_X1 U709 ( .A1(n779), .A2(G53), .ZN(n628) );
  NAND2_X1 U710 ( .A1(G65), .A2(n772), .ZN(n627) );
  NAND2_X1 U711 ( .A1(n628), .A2(n627), .ZN(n632) );
  NAND2_X1 U712 ( .A1(n771), .A2(G78), .ZN(n630) );
  NAND2_X1 U713 ( .A1(G91), .A2(n775), .ZN(n629) );
  NAND2_X1 U714 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U715 ( .A1(n632), .A2(n631), .ZN(n965) );
  NAND2_X1 U716 ( .A1(n633), .A2(G2072), .ZN(n635) );
  INV_X1 U717 ( .A(KEYINPUT27), .ZN(n634) );
  XNOR2_X1 U718 ( .A(n635), .B(n634), .ZN(n637) );
  NAND2_X1 U719 ( .A1(G1956), .A2(n652), .ZN(n636) );
  NAND2_X1 U720 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U721 ( .A(n638), .B(KEYINPUT98), .Z(n673) );
  INV_X1 U722 ( .A(KEYINPUT28), .ZN(n639) );
  XNOR2_X1 U723 ( .A(n640), .B(n639), .ZN(n677) );
  NAND2_X1 U724 ( .A1(G56), .A2(n772), .ZN(n641) );
  XOR2_X1 U725 ( .A(KEYINPUT14), .B(n641), .Z(n649) );
  NAND2_X1 U726 ( .A1(n771), .A2(G68), .ZN(n642) );
  XNOR2_X1 U727 ( .A(KEYINPUT77), .B(n642), .ZN(n645) );
  NAND2_X1 U728 ( .A1(G81), .A2(n775), .ZN(n643) );
  XOR2_X1 U729 ( .A(n643), .B(KEYINPUT12), .Z(n644) );
  NOR2_X1 U730 ( .A1(n645), .A2(n644), .ZN(n647) );
  NOR2_X1 U731 ( .A1(n649), .A2(n648), .ZN(n651) );
  NAND2_X1 U732 ( .A1(n779), .A2(G43), .ZN(n650) );
  INV_X1 U733 ( .A(G1996), .ZN(n821) );
  NOR2_X1 U734 ( .A1(n652), .A2(n821), .ZN(n654) );
  INV_X1 U735 ( .A(KEYINPUT26), .ZN(n653) );
  XNOR2_X1 U736 ( .A(n654), .B(n653), .ZN(n656) );
  NAND2_X1 U737 ( .A1(n689), .A2(G1341), .ZN(n655) );
  NAND2_X1 U738 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U739 ( .A1(n975), .A2(n657), .ZN(n669) );
  NAND2_X1 U740 ( .A1(G54), .A2(n779), .ZN(n659) );
  NAND2_X1 U741 ( .A1(G92), .A2(n775), .ZN(n658) );
  NAND2_X1 U742 ( .A1(n659), .A2(n658), .ZN(n663) );
  NAND2_X1 U743 ( .A1(n771), .A2(G79), .ZN(n661) );
  NAND2_X1 U744 ( .A1(G66), .A2(n772), .ZN(n660) );
  NAND2_X1 U745 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U746 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U747 ( .A(n664), .B(KEYINPUT15), .Z(n956) );
  INV_X1 U748 ( .A(n956), .ZN(n766) );
  NAND2_X1 U749 ( .A1(G1348), .A2(n689), .ZN(n667) );
  NAND2_X1 U750 ( .A1(G2067), .A2(n665), .ZN(n666) );
  NAND2_X1 U751 ( .A1(n667), .A2(n666), .ZN(n670) );
  NOR2_X1 U752 ( .A1(n766), .A2(n670), .ZN(n668) );
  OR2_X1 U753 ( .A1(n669), .A2(n668), .ZN(n672) );
  NAND2_X1 U754 ( .A1(n766), .A2(n670), .ZN(n671) );
  NAND2_X1 U755 ( .A1(n672), .A2(n671), .ZN(n675) );
  NAND2_X1 U756 ( .A1(n965), .A2(n673), .ZN(n674) );
  NAND2_X1 U757 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U758 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U759 ( .A(KEYINPUT29), .B(n678), .Z(n681) );
  OR2_X1 U760 ( .A1(n679), .A2(G301), .ZN(n680) );
  NAND2_X1 U761 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U762 ( .A1(n683), .A2(n682), .ZN(n688) );
  XOR2_X1 U763 ( .A(n688), .B(KEYINPUT100), .Z(n684) );
  NOR2_X1 U764 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U765 ( .A1(n687), .A2(n686), .ZN(n700) );
  NAND2_X1 U766 ( .A1(n688), .A2(G286), .ZN(n696) );
  NOR2_X1 U767 ( .A1(G2090), .A2(n689), .ZN(n690) );
  XOR2_X1 U768 ( .A(KEYINPUT101), .B(n690), .Z(n692) );
  NOR2_X1 U769 ( .A1(G1971), .A2(n721), .ZN(n691) );
  NOR2_X1 U770 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U771 ( .A(n693), .B(KEYINPUT102), .ZN(n694) );
  NAND2_X1 U772 ( .A1(n694), .A2(G303), .ZN(n695) );
  NAND2_X1 U773 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U774 ( .A1(n697), .A2(G8), .ZN(n698) );
  NAND2_X1 U775 ( .A1(n700), .A2(n699), .ZN(n715) );
  NOR2_X1 U776 ( .A1(G1976), .A2(G288), .ZN(n708) );
  NOR2_X1 U777 ( .A1(G1971), .A2(G303), .ZN(n701) );
  NOR2_X1 U778 ( .A1(n708), .A2(n701), .ZN(n969) );
  NAND2_X1 U779 ( .A1(n715), .A2(n969), .ZN(n703) );
  XNOR2_X1 U780 ( .A(n703), .B(n702), .ZN(n706) );
  NAND2_X1 U781 ( .A1(G1976), .A2(G288), .ZN(n964) );
  INV_X1 U782 ( .A(n964), .ZN(n704) );
  NOR2_X1 U783 ( .A1(n721), .A2(n704), .ZN(n705) );
  AND2_X1 U784 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U785 ( .A1(n707), .A2(KEYINPUT33), .ZN(n711) );
  NAND2_X1 U786 ( .A1(n708), .A2(KEYINPUT33), .ZN(n709) );
  NOR2_X1 U787 ( .A1(n709), .A2(n721), .ZN(n710) );
  NOR2_X1 U788 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U789 ( .A(G1981), .B(G305), .Z(n960) );
  NAND2_X1 U790 ( .A1(n712), .A2(n960), .ZN(n725) );
  NOR2_X1 U791 ( .A1(G2090), .A2(G303), .ZN(n713) );
  XNOR2_X1 U792 ( .A(n713), .B(KEYINPUT104), .ZN(n714) );
  NAND2_X1 U793 ( .A1(n714), .A2(G8), .ZN(n716) );
  NAND2_X1 U794 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U795 ( .A(KEYINPUT105), .B(n717), .Z(n718) );
  AND2_X1 U796 ( .A1(n718), .A2(n721), .ZN(n723) );
  NOR2_X1 U797 ( .A1(G1981), .A2(G305), .ZN(n719) );
  XOR2_X1 U798 ( .A(n719), .B(KEYINPUT24), .Z(n720) );
  NOR2_X1 U799 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U800 ( .A1(n723), .A2(n722), .ZN(n724) );
  AND2_X1 U801 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U802 ( .A1(n727), .A2(n726), .ZN(n729) );
  XNOR2_X1 U803 ( .A(G1986), .B(G290), .ZN(n971) );
  NAND2_X1 U804 ( .A1(n971), .A2(n739), .ZN(n728) );
  NAND2_X1 U805 ( .A1(n729), .A2(n728), .ZN(n742) );
  NOR2_X1 U806 ( .A1(G1996), .A2(n870), .ZN(n905) );
  NOR2_X1 U807 ( .A1(n935), .A2(n866), .ZN(n908) );
  NOR2_X1 U808 ( .A1(G1986), .A2(G290), .ZN(n730) );
  NOR2_X1 U809 ( .A1(n908), .A2(n730), .ZN(n731) );
  NOR2_X1 U810 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U811 ( .A1(n905), .A2(n733), .ZN(n734) );
  XNOR2_X1 U812 ( .A(n734), .B(KEYINPUT39), .ZN(n736) );
  NAND2_X1 U813 ( .A1(n736), .A2(n735), .ZN(n738) );
  NAND2_X1 U814 ( .A1(n737), .A2(n871), .ZN(n914) );
  NAND2_X1 U815 ( .A1(n738), .A2(n914), .ZN(n740) );
  NAND2_X1 U816 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U817 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U818 ( .A(n743), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U819 ( .A1(n745), .A2(n744), .ZN(G160) );
  AND2_X1 U820 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U821 ( .A1(G99), .A2(n858), .ZN(n752) );
  NAND2_X1 U822 ( .A1(G135), .A2(n861), .ZN(n747) );
  NAND2_X1 U823 ( .A1(G111), .A2(n852), .ZN(n746) );
  NAND2_X1 U824 ( .A1(n747), .A2(n746), .ZN(n750) );
  NAND2_X1 U825 ( .A1(n854), .A2(G123), .ZN(n748) );
  XOR2_X1 U826 ( .A(KEYINPUT18), .B(n748), .Z(n749) );
  NOR2_X1 U827 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U828 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U829 ( .A(n753), .B(KEYINPUT82), .ZN(n910) );
  XNOR2_X1 U830 ( .A(n910), .B(G2096), .ZN(n754) );
  OR2_X1 U831 ( .A1(G2100), .A2(n754), .ZN(G156) );
  INV_X1 U832 ( .A(n965), .ZN(G299) );
  INV_X1 U833 ( .A(G82), .ZN(G220) );
  XOR2_X1 U834 ( .A(KEYINPUT75), .B(KEYINPUT10), .Z(n756) );
  NAND2_X1 U835 ( .A1(G7), .A2(G661), .ZN(n755) );
  XNOR2_X1 U836 ( .A(n756), .B(n755), .ZN(n757) );
  XNOR2_X1 U837 ( .A(KEYINPUT74), .B(n757), .ZN(G223) );
  XOR2_X1 U838 ( .A(KEYINPUT76), .B(G223), .Z(n812) );
  NAND2_X1 U839 ( .A1(n812), .A2(G567), .ZN(n758) );
  XOR2_X1 U840 ( .A(KEYINPUT11), .B(n758), .Z(G234) );
  INV_X1 U841 ( .A(G860), .ZN(n763) );
  OR2_X1 U842 ( .A1(n975), .A2(n763), .ZN(G153) );
  NAND2_X1 U843 ( .A1(G868), .A2(G301), .ZN(n760) );
  INV_X1 U844 ( .A(G868), .ZN(n793) );
  NAND2_X1 U845 ( .A1(n766), .A2(n793), .ZN(n759) );
  NAND2_X1 U846 ( .A1(n760), .A2(n759), .ZN(G284) );
  NOR2_X1 U847 ( .A1(G286), .A2(n793), .ZN(n762) );
  NOR2_X1 U848 ( .A1(G868), .A2(G299), .ZN(n761) );
  NOR2_X1 U849 ( .A1(n762), .A2(n761), .ZN(G297) );
  NAND2_X1 U850 ( .A1(n763), .A2(G559), .ZN(n764) );
  NAND2_X1 U851 ( .A1(n764), .A2(n956), .ZN(n765) );
  XNOR2_X1 U852 ( .A(n765), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U853 ( .A1(n766), .A2(n793), .ZN(n767) );
  XNOR2_X1 U854 ( .A(n767), .B(KEYINPUT81), .ZN(n768) );
  NOR2_X1 U855 ( .A1(G559), .A2(n768), .ZN(n770) );
  NOR2_X1 U856 ( .A1(G868), .A2(n975), .ZN(n769) );
  NOR2_X1 U857 ( .A1(n770), .A2(n769), .ZN(G282) );
  NAND2_X1 U858 ( .A1(n771), .A2(G80), .ZN(n774) );
  NAND2_X1 U859 ( .A1(G67), .A2(n772), .ZN(n773) );
  NAND2_X1 U860 ( .A1(n774), .A2(n773), .ZN(n778) );
  NAND2_X1 U861 ( .A1(G93), .A2(n775), .ZN(n776) );
  XNOR2_X1 U862 ( .A(KEYINPUT83), .B(n776), .ZN(n777) );
  NOR2_X1 U863 ( .A1(n778), .A2(n777), .ZN(n781) );
  NAND2_X1 U864 ( .A1(n779), .A2(G55), .ZN(n780) );
  NAND2_X1 U865 ( .A1(n781), .A2(n780), .ZN(n795) );
  NAND2_X1 U866 ( .A1(n956), .A2(G559), .ZN(n792) );
  XNOR2_X1 U867 ( .A(n975), .B(n792), .ZN(n782) );
  NOR2_X1 U868 ( .A1(G860), .A2(n782), .ZN(n783) );
  XOR2_X1 U869 ( .A(n795), .B(n783), .Z(G145) );
  XNOR2_X1 U870 ( .A(KEYINPUT19), .B(G288), .ZN(n784) );
  XNOR2_X1 U871 ( .A(n784), .B(n795), .ZN(n787) );
  XOR2_X1 U872 ( .A(G299), .B(G290), .Z(n785) );
  XOR2_X1 U873 ( .A(n785), .B(G166), .Z(n786) );
  XNOR2_X1 U874 ( .A(n787), .B(n786), .ZN(n789) );
  XNOR2_X1 U875 ( .A(G305), .B(KEYINPUT86), .ZN(n788) );
  XNOR2_X1 U876 ( .A(n789), .B(n788), .ZN(n790) );
  XNOR2_X1 U877 ( .A(n790), .B(n975), .ZN(n882) );
  XOR2_X1 U878 ( .A(n882), .B(KEYINPUT87), .Z(n791) );
  XNOR2_X1 U879 ( .A(n792), .B(n791), .ZN(n794) );
  NOR2_X1 U880 ( .A1(n794), .A2(n793), .ZN(n797) );
  NOR2_X1 U881 ( .A1(G868), .A2(n795), .ZN(n796) );
  NOR2_X1 U882 ( .A1(n797), .A2(n796), .ZN(G295) );
  NAND2_X1 U883 ( .A1(G2084), .A2(G2078), .ZN(n799) );
  XOR2_X1 U884 ( .A(KEYINPUT88), .B(KEYINPUT20), .Z(n798) );
  XNOR2_X1 U885 ( .A(n799), .B(n798), .ZN(n800) );
  NAND2_X1 U886 ( .A1(G2090), .A2(n800), .ZN(n801) );
  XNOR2_X1 U887 ( .A(KEYINPUT21), .B(n801), .ZN(n802) );
  NAND2_X1 U888 ( .A1(n802), .A2(G2072), .ZN(G158) );
  XOR2_X1 U889 ( .A(KEYINPUT72), .B(G57), .Z(G237) );
  XNOR2_X1 U890 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U891 ( .A(KEYINPUT73), .B(G132), .ZN(G219) );
  NAND2_X1 U892 ( .A1(G108), .A2(G120), .ZN(n803) );
  NOR2_X1 U893 ( .A1(G237), .A2(n803), .ZN(n804) );
  NAND2_X1 U894 ( .A1(G69), .A2(n804), .ZN(n816) );
  NAND2_X1 U895 ( .A1(n816), .A2(G567), .ZN(n809) );
  NOR2_X1 U896 ( .A1(G220), .A2(G219), .ZN(n805) );
  XOR2_X1 U897 ( .A(KEYINPUT22), .B(n805), .Z(n806) );
  NOR2_X1 U898 ( .A1(G218), .A2(n806), .ZN(n807) );
  NAND2_X1 U899 ( .A1(G96), .A2(n807), .ZN(n817) );
  NAND2_X1 U900 ( .A1(n817), .A2(G2106), .ZN(n808) );
  NAND2_X1 U901 ( .A1(n809), .A2(n808), .ZN(n818) );
  NAND2_X1 U902 ( .A1(G661), .A2(G483), .ZN(n810) );
  XOR2_X1 U903 ( .A(KEYINPUT89), .B(n810), .Z(n811) );
  NOR2_X1 U904 ( .A1(n818), .A2(n811), .ZN(n815) );
  NAND2_X1 U905 ( .A1(n815), .A2(G36), .ZN(G176) );
  NAND2_X1 U906 ( .A1(G2106), .A2(n812), .ZN(G217) );
  AND2_X1 U907 ( .A1(G15), .A2(G2), .ZN(n813) );
  NAND2_X1 U908 ( .A1(G661), .A2(n813), .ZN(G259) );
  NAND2_X1 U909 ( .A1(G3), .A2(G1), .ZN(n814) );
  NAND2_X1 U910 ( .A1(n815), .A2(n814), .ZN(G188) );
  INV_X1 U912 ( .A(G120), .ZN(G236) );
  INV_X1 U913 ( .A(G108), .ZN(G238) );
  INV_X1 U914 ( .A(G96), .ZN(G221) );
  INV_X1 U915 ( .A(G69), .ZN(G235) );
  NOR2_X1 U916 ( .A1(n817), .A2(n816), .ZN(G325) );
  INV_X1 U917 ( .A(G325), .ZN(G261) );
  INV_X1 U918 ( .A(n818), .ZN(G319) );
  XNOR2_X1 U919 ( .A(G1961), .B(KEYINPUT41), .ZN(n829) );
  XOR2_X1 U920 ( .A(G1976), .B(G1971), .Z(n820) );
  XNOR2_X1 U921 ( .A(G1986), .B(G1956), .ZN(n819) );
  XNOR2_X1 U922 ( .A(n820), .B(n819), .ZN(n825) );
  XOR2_X1 U923 ( .A(G1981), .B(G1966), .Z(n823) );
  XOR2_X1 U924 ( .A(n821), .B(G1991), .Z(n822) );
  XNOR2_X1 U925 ( .A(n823), .B(n822), .ZN(n824) );
  XOR2_X1 U926 ( .A(n825), .B(n824), .Z(n827) );
  XNOR2_X1 U927 ( .A(G2474), .B(KEYINPUT108), .ZN(n826) );
  XNOR2_X1 U928 ( .A(n827), .B(n826), .ZN(n828) );
  XNOR2_X1 U929 ( .A(n829), .B(n828), .ZN(G229) );
  XOR2_X1 U930 ( .A(G2100), .B(G2096), .Z(n831) );
  XNOR2_X1 U931 ( .A(KEYINPUT42), .B(G2678), .ZN(n830) );
  XNOR2_X1 U932 ( .A(n831), .B(n830), .ZN(n835) );
  XOR2_X1 U933 ( .A(KEYINPUT43), .B(G2090), .Z(n833) );
  XNOR2_X1 U934 ( .A(G2067), .B(G2072), .ZN(n832) );
  XNOR2_X1 U935 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U936 ( .A(n835), .B(n834), .Z(n837) );
  XNOR2_X1 U937 ( .A(G2084), .B(G2078), .ZN(n836) );
  XNOR2_X1 U938 ( .A(n837), .B(n836), .ZN(G227) );
  NAND2_X1 U939 ( .A1(G136), .A2(n861), .ZN(n839) );
  NAND2_X1 U940 ( .A1(G112), .A2(n852), .ZN(n838) );
  NAND2_X1 U941 ( .A1(n839), .A2(n838), .ZN(n844) );
  NAND2_X1 U942 ( .A1(G124), .A2(n854), .ZN(n840) );
  XNOR2_X1 U943 ( .A(n840), .B(KEYINPUT44), .ZN(n842) );
  NAND2_X1 U944 ( .A1(n858), .A2(G100), .ZN(n841) );
  NAND2_X1 U945 ( .A1(n842), .A2(n841), .ZN(n843) );
  NOR2_X1 U946 ( .A1(n844), .A2(n843), .ZN(G162) );
  NAND2_X1 U947 ( .A1(G118), .A2(n852), .ZN(n846) );
  NAND2_X1 U948 ( .A1(G130), .A2(n854), .ZN(n845) );
  NAND2_X1 U949 ( .A1(n846), .A2(n845), .ZN(n851) );
  NAND2_X1 U950 ( .A1(G142), .A2(n861), .ZN(n848) );
  NAND2_X1 U951 ( .A1(G106), .A2(n858), .ZN(n847) );
  NAND2_X1 U952 ( .A1(n848), .A2(n847), .ZN(n849) );
  XOR2_X1 U953 ( .A(KEYINPUT45), .B(n849), .Z(n850) );
  NOR2_X1 U954 ( .A1(n851), .A2(n850), .ZN(n865) );
  NAND2_X1 U955 ( .A1(n852), .A2(G115), .ZN(n853) );
  XNOR2_X1 U956 ( .A(n853), .B(KEYINPUT112), .ZN(n856) );
  NAND2_X1 U957 ( .A1(G127), .A2(n854), .ZN(n855) );
  NAND2_X1 U958 ( .A1(n856), .A2(n855), .ZN(n857) );
  XNOR2_X1 U959 ( .A(n857), .B(KEYINPUT47), .ZN(n860) );
  NAND2_X1 U960 ( .A1(G103), .A2(n858), .ZN(n859) );
  NAND2_X1 U961 ( .A1(n860), .A2(n859), .ZN(n864) );
  NAND2_X1 U962 ( .A1(G139), .A2(n861), .ZN(n862) );
  XNOR2_X1 U963 ( .A(KEYINPUT111), .B(n862), .ZN(n863) );
  NOR2_X1 U964 ( .A1(n864), .A2(n863), .ZN(n916) );
  XOR2_X1 U965 ( .A(n865), .B(n916), .Z(n868) );
  XOR2_X1 U966 ( .A(G164), .B(n866), .Z(n867) );
  XNOR2_X1 U967 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U968 ( .A(n869), .B(G162), .Z(n873) );
  XNOR2_X1 U969 ( .A(n871), .B(n870), .ZN(n872) );
  XNOR2_X1 U970 ( .A(n873), .B(n872), .ZN(n880) );
  XOR2_X1 U971 ( .A(KEYINPUT46), .B(KEYINPUT109), .Z(n875) );
  XNOR2_X1 U972 ( .A(n910), .B(KEYINPUT48), .ZN(n874) );
  XNOR2_X1 U973 ( .A(n875), .B(n874), .ZN(n876) );
  XOR2_X1 U974 ( .A(n876), .B(KEYINPUT110), .Z(n878) );
  XNOR2_X1 U975 ( .A(G160), .B(KEYINPUT113), .ZN(n877) );
  XNOR2_X1 U976 ( .A(n878), .B(n877), .ZN(n879) );
  XNOR2_X1 U977 ( .A(n880), .B(n879), .ZN(n881) );
  NOR2_X1 U978 ( .A1(G37), .A2(n881), .ZN(G395) );
  XNOR2_X1 U979 ( .A(n882), .B(KEYINPUT114), .ZN(n884) );
  XOR2_X1 U980 ( .A(n956), .B(G286), .Z(n883) );
  XNOR2_X1 U981 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U982 ( .A(n885), .B(G301), .Z(n886) );
  NOR2_X1 U983 ( .A1(G37), .A2(n886), .ZN(G397) );
  XNOR2_X1 U984 ( .A(G2451), .B(G2443), .ZN(n896) );
  XOR2_X1 U985 ( .A(G2446), .B(G2430), .Z(n888) );
  XNOR2_X1 U986 ( .A(KEYINPUT107), .B(G2438), .ZN(n887) );
  XNOR2_X1 U987 ( .A(n888), .B(n887), .ZN(n892) );
  XOR2_X1 U988 ( .A(G2435), .B(G2454), .Z(n890) );
  XNOR2_X1 U989 ( .A(G1341), .B(G1348), .ZN(n889) );
  XNOR2_X1 U990 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U991 ( .A(n892), .B(n891), .Z(n894) );
  XNOR2_X1 U992 ( .A(KEYINPUT106), .B(G2427), .ZN(n893) );
  XNOR2_X1 U993 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U994 ( .A(n896), .B(n895), .ZN(n897) );
  NAND2_X1 U995 ( .A1(n897), .A2(G14), .ZN(n903) );
  NAND2_X1 U996 ( .A1(G319), .A2(n903), .ZN(n900) );
  NOR2_X1 U997 ( .A1(G229), .A2(G227), .ZN(n898) );
  XNOR2_X1 U998 ( .A(KEYINPUT49), .B(n898), .ZN(n899) );
  NOR2_X1 U999 ( .A1(n900), .A2(n899), .ZN(n902) );
  NOR2_X1 U1000 ( .A1(G395), .A2(G397), .ZN(n901) );
  NAND2_X1 U1001 ( .A1(n902), .A2(n901), .ZN(G225) );
  INV_X1 U1002 ( .A(G225), .ZN(G308) );
  INV_X1 U1003 ( .A(n903), .ZN(G401) );
  XOR2_X1 U1004 ( .A(G2090), .B(G162), .Z(n904) );
  NOR2_X1 U1005 ( .A1(n905), .A2(n904), .ZN(n906) );
  XNOR2_X1 U1006 ( .A(n906), .B(KEYINPUT51), .ZN(n907) );
  NOR2_X1 U1007 ( .A1(n908), .A2(n907), .ZN(n909) );
  NAND2_X1 U1008 ( .A1(n910), .A2(n909), .ZN(n913) );
  XNOR2_X1 U1009 ( .A(G2084), .B(G160), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(KEYINPUT115), .B(n911), .ZN(n912) );
  NOR2_X1 U1011 ( .A1(n913), .A2(n912), .ZN(n924) );
  NAND2_X1 U1012 ( .A1(n915), .A2(n914), .ZN(n922) );
  XOR2_X1 U1013 ( .A(G2072), .B(n916), .Z(n918) );
  XOR2_X1 U1014 ( .A(G164), .B(G2078), .Z(n917) );
  NOR2_X1 U1015 ( .A1(n918), .A2(n917), .ZN(n919) );
  XOR2_X1 U1016 ( .A(KEYINPUT116), .B(n919), .Z(n920) );
  XNOR2_X1 U1017 ( .A(KEYINPUT50), .B(n920), .ZN(n921) );
  NOR2_X1 U1018 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1019 ( .A1(n924), .A2(n923), .ZN(n925) );
  NOR2_X1 U1020 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1021 ( .A(KEYINPUT52), .B(n927), .ZN(n928) );
  XNOR2_X1 U1022 ( .A(KEYINPUT55), .B(KEYINPUT117), .ZN(n952) );
  NAND2_X1 U1023 ( .A1(n928), .A2(n952), .ZN(n929) );
  NAND2_X1 U1024 ( .A1(n929), .A2(G29), .ZN(n1012) );
  XOR2_X1 U1025 ( .A(G32), .B(G1996), .Z(n930) );
  NAND2_X1 U1026 ( .A1(n930), .A2(G28), .ZN(n942) );
  XOR2_X1 U1027 ( .A(G2072), .B(G33), .Z(n931) );
  XNOR2_X1 U1028 ( .A(KEYINPUT119), .B(n931), .ZN(n933) );
  XNOR2_X1 U1029 ( .A(G26), .B(G2067), .ZN(n932) );
  NOR2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1031 ( .A(KEYINPUT120), .B(n934), .ZN(n940) );
  XNOR2_X1 U1032 ( .A(n935), .B(G25), .ZN(n938) );
  XNOR2_X1 U1033 ( .A(n936), .B(G27), .ZN(n937) );
  NOR2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  NOR2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n944) );
  XNOR2_X1 U1037 ( .A(KEYINPUT53), .B(KEYINPUT121), .ZN(n943) );
  XNOR2_X1 U1038 ( .A(n944), .B(n943), .ZN(n950) );
  XNOR2_X1 U1039 ( .A(G2084), .B(G34), .ZN(n945) );
  XNOR2_X1 U1040 ( .A(n945), .B(KEYINPUT54), .ZN(n948) );
  XNOR2_X1 U1041 ( .A(G2090), .B(KEYINPUT118), .ZN(n946) );
  XNOR2_X1 U1042 ( .A(n946), .B(G35), .ZN(n947) );
  NOR2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1045 ( .A(n952), .B(n951), .ZN(n954) );
  INV_X1 U1046 ( .A(G29), .ZN(n953) );
  NAND2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1048 ( .A1(G11), .A2(n955), .ZN(n1010) );
  XNOR2_X1 U1049 ( .A(KEYINPUT56), .B(G16), .ZN(n981) );
  XOR2_X1 U1050 ( .A(G171), .B(G1961), .Z(n958) );
  XOR2_X1 U1051 ( .A(n956), .B(G1348), .Z(n957) );
  NOR2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1053 ( .A(KEYINPUT122), .B(n959), .ZN(n979) );
  XNOR2_X1 U1054 ( .A(G1966), .B(G168), .ZN(n961) );
  NAND2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1056 ( .A(n962), .B(KEYINPUT57), .ZN(n974) );
  NAND2_X1 U1057 ( .A1(G1971), .A2(G303), .ZN(n963) );
  NAND2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n967) );
  XOR2_X1 U1059 ( .A(G1956), .B(n965), .Z(n966) );
  NOR2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n970) );
  NOR2_X1 U1062 ( .A1(n971), .A2(n970), .ZN(n972) );
  XOR2_X1 U1063 ( .A(KEYINPUT123), .B(n972), .Z(n973) );
  NAND2_X1 U1064 ( .A1(n974), .A2(n973), .ZN(n977) );
  XNOR2_X1 U1065 ( .A(G1341), .B(n975), .ZN(n976) );
  NOR2_X1 U1066 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1067 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1068 ( .A1(n981), .A2(n980), .ZN(n1008) );
  XOR2_X1 U1069 ( .A(G16), .B(KEYINPUT124), .Z(n1006) );
  XNOR2_X1 U1070 ( .A(G1966), .B(G21), .ZN(n983) );
  XNOR2_X1 U1071 ( .A(G5), .B(G1961), .ZN(n982) );
  NOR2_X1 U1072 ( .A1(n983), .A2(n982), .ZN(n993) );
  XOR2_X1 U1073 ( .A(G1348), .B(KEYINPUT59), .Z(n984) );
  XNOR2_X1 U1074 ( .A(G4), .B(n984), .ZN(n986) );
  XNOR2_X1 U1075 ( .A(G20), .B(G1956), .ZN(n985) );
  NOR2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n990) );
  XNOR2_X1 U1077 ( .A(G1341), .B(G19), .ZN(n988) );
  XNOR2_X1 U1078 ( .A(G1981), .B(G6), .ZN(n987) );
  NOR2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1081 ( .A(KEYINPUT60), .B(n991), .Z(n992) );
  NAND2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n1003) );
  XOR2_X1 U1083 ( .A(G1986), .B(G24), .Z(n999) );
  XOR2_X1 U1084 ( .A(G1976), .B(KEYINPUT125), .Z(n994) );
  XNOR2_X1 U1085 ( .A(G23), .B(n994), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(G22), .B(G1971), .ZN(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1088 ( .A(n997), .B(KEYINPUT126), .ZN(n998) );
  NAND2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1090 ( .A(KEYINPUT58), .B(n1000), .Z(n1001) );
  XNOR2_X1 U1091 ( .A(KEYINPUT127), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(n1004), .B(KEYINPUT61), .ZN(n1005) );
  NAND2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1097 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1098 ( .A(KEYINPUT62), .B(n1013), .ZN(G150) );
  INV_X1 U1099 ( .A(G150), .ZN(G311) );
endmodule

