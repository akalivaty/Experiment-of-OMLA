//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 1 0 0 0 0 1 0 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 0 0 1 1 1 0 0 0 0 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1292, new_n1293, new_n1294, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  XNOR2_X1  g0012(.A(KEYINPUT64), .B(G20), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  INV_X1    g0025(.A(G58), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  INV_X1    g0027(.A(G97), .ZN(new_n228));
  INV_X1    g0028(.A(G257), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n225), .B1(new_n226), .B2(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n209), .B1(new_n224), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n212), .B(new_n218), .C1(KEYINPUT1), .C2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n202), .A2(G68), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n220), .A2(G50), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n244), .B(new_n249), .ZN(G351));
  NAND2_X1  g0050(.A1(new_n213), .A2(G33), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT70), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n213), .A2(KEYINPUT70), .A3(G33), .ZN(new_n254));
  XOR2_X1   g0054(.A(KEYINPUT8), .B(G58), .Z(new_n255));
  NAND3_X1  g0055(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G20), .A2(G33), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n214), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(new_n261), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n202), .B1(new_n206), .B2(G20), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n265), .A2(new_n266), .B1(new_n202), .B2(new_n264), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n268), .B(KEYINPUT9), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT66), .ZN(new_n270));
  INV_X1    g0070(.A(G274), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n214), .B1(KEYINPUT65), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT65), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G33), .A3(G41), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n271), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G41), .A2(G45), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(G1), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n270), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n272), .A2(KEYINPUT65), .ZN(new_n280));
  AND2_X1   g0080(.A1(G1), .A2(G13), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n280), .A2(new_n275), .A3(new_n281), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n282), .A2(new_n270), .A3(G274), .A4(new_n278), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n279), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT67), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n286), .B1(new_n277), .B2(G1), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n206), .B(KEYINPUT67), .C1(G41), .C2(G45), .ZN(new_n288));
  AND3_X1   g0088(.A1(new_n282), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n285), .B1(G226), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n281), .A2(new_n272), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT3), .B(G33), .ZN(new_n293));
  INV_X1    g0093(.A(G77), .ZN(new_n294));
  OAI21_X1  g0094(.A(KEYINPUT68), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G1698), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n293), .A2(G222), .A3(new_n296), .ZN(new_n297));
  MUX2_X1   g0097(.A(KEYINPUT68), .B(new_n295), .S(new_n297), .Z(new_n298));
  INV_X1    g0098(.A(G223), .ZN(new_n299));
  INV_X1    g0099(.A(G33), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT3), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT3), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G33), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n301), .A2(new_n303), .A3(G1698), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT69), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n293), .A2(KEYINPUT69), .A3(G1698), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n299), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n292), .B1(new_n298), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n290), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G200), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n290), .A2(new_n309), .A3(G190), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n269), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT10), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT10), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n269), .A2(new_n315), .A3(new_n311), .A4(new_n312), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G169), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n310), .A2(new_n318), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n319), .B(new_n268), .C1(G179), .C2(new_n310), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G226), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n296), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n227), .A2(G1698), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n301), .A2(new_n323), .A3(new_n303), .A4(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(G33), .A2(G97), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT73), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(KEYINPUT73), .A2(G33), .A3(G97), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n282), .A2(new_n287), .A3(new_n288), .ZN(new_n332));
  OAI22_X1  g0132(.A1(new_n331), .A2(new_n291), .B1(new_n332), .B2(new_n221), .ZN(new_n333));
  NOR3_X1   g0133(.A1(new_n285), .A2(new_n333), .A3(KEYINPUT13), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT13), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n291), .B1(new_n325), .B2(new_n330), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n336), .B1(new_n289), .B2(G238), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n282), .A2(G274), .A3(new_n278), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT66), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n283), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n335), .B1(new_n337), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n334), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(KEYINPUT14), .B1(new_n342), .B2(new_n318), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT14), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n344), .B(G169), .C1(new_n334), .C2(new_n341), .ZN(new_n345));
  OAI21_X1  g0145(.A(KEYINPUT74), .B1(new_n285), .B2(new_n333), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT74), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n337), .A2(new_n340), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n346), .A2(KEYINPUT13), .A3(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G179), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n285), .A2(new_n333), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n350), .B1(new_n351), .B2(new_n335), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT76), .ZN(new_n353));
  AND3_X1   g0153(.A1(new_n349), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n353), .B1(new_n349), .B2(new_n352), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n343), .B(new_n345), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n261), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n253), .A2(G77), .A3(new_n254), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n257), .A2(G50), .B1(G20), .B2(new_n220), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n360), .A2(KEYINPUT11), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n206), .A2(G20), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n265), .A2(G68), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT75), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n363), .B(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n264), .A2(new_n220), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n366), .B(KEYINPUT12), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n360), .A2(KEYINPUT11), .ZN(new_n369));
  NOR3_X1   g0169(.A1(new_n361), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n356), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(G200), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n370), .B1(new_n373), .B2(new_n342), .ZN(new_n374));
  INV_X1    g0174(.A(G190), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n334), .A2(new_n375), .ZN(new_n376));
  AND2_X1   g0176(.A1(new_n376), .A2(new_n349), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n372), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n301), .A2(new_n303), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n381), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n382));
  AOI21_X1  g0182(.A(KEYINPUT7), .B1(new_n381), .B2(new_n213), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT77), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AOI211_X1 g0185(.A(KEYINPUT77), .B(KEYINPUT7), .C1(new_n381), .C2(new_n213), .ZN(new_n386));
  OAI21_X1  g0186(.A(G68), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n226), .A2(new_n220), .ZN(new_n388));
  OAI21_X1  g0188(.A(G20), .B1(new_n388), .B2(new_n201), .ZN(new_n389));
  INV_X1    g0189(.A(G159), .ZN(new_n390));
  INV_X1    g0190(.A(new_n257), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(KEYINPUT78), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT78), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n389), .B(new_n394), .C1(new_n390), .C2(new_n391), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n387), .A2(KEYINPUT16), .A3(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT16), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n301), .A2(KEYINPUT79), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT79), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n400), .A2(new_n300), .A3(KEYINPUT3), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n399), .A2(new_n303), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n402), .A2(KEYINPUT7), .A3(new_n213), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT7), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(new_n293), .B2(G20), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n220), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n398), .B1(new_n406), .B2(new_n392), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n397), .A2(new_n261), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n299), .A2(new_n296), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n322), .A2(G1698), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n301), .A2(new_n409), .A3(new_n303), .A4(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G33), .A2(G87), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n291), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n413), .B1(new_n289), .B2(G232), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n414), .A2(new_n340), .A3(new_n375), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n414), .A2(new_n340), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n415), .B1(new_n416), .B2(G200), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n255), .A2(new_n362), .ZN(new_n418));
  INV_X1    g0218(.A(new_n255), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n418), .A2(new_n265), .B1(new_n264), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n408), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT80), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n422), .A2(KEYINPUT17), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g0225(.A(KEYINPUT80), .B(KEYINPUT17), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n408), .A2(new_n417), .A3(new_n420), .A4(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n408), .A2(new_n420), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n318), .B1(new_n414), .B2(new_n340), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n431), .B1(G179), .B2(new_n416), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT18), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT18), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n430), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n429), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n339), .A2(new_n283), .B1(new_n289), .B2(G244), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n221), .B1(new_n306), .B2(new_n307), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n227), .A2(G1698), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n441), .A2(new_n301), .A3(new_n303), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT71), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n293), .A2(KEYINPUT71), .A3(new_n441), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n381), .A2(G107), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n292), .B1(new_n440), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT72), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n439), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n449), .B1(new_n439), .B2(new_n448), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n350), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  AND3_X1   g0252(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT69), .B1(new_n293), .B2(G1698), .ZN(new_n454));
  AND4_X1   g0254(.A1(KEYINPUT69), .A2(new_n301), .A3(new_n303), .A4(G1698), .ZN(new_n455));
  OAI21_X1  g0255(.A(G238), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n291), .B1(new_n453), .B2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n282), .A2(G244), .A3(new_n287), .A4(new_n288), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n458), .B1(new_n279), .B2(new_n284), .ZN(new_n459));
  OAI21_X1  g0259(.A(KEYINPUT72), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n439), .A2(new_n448), .A3(new_n449), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n460), .A2(new_n318), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n207), .A2(KEYINPUT64), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT64), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G20), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n255), .A2(new_n257), .B1(new_n466), .B2(G77), .ZN(new_n467));
  XNOR2_X1  g0267(.A(KEYINPUT15), .B(G87), .ZN(new_n468));
  OR2_X1    g0268(.A1(new_n251), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n357), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n265), .A2(G77), .A3(new_n362), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n471), .B1(G77), .B2(new_n263), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n452), .A2(new_n462), .A3(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(G190), .B1(new_n450), .B2(new_n451), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n460), .A2(G200), .A3(new_n461), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n476), .A2(new_n473), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  NOR4_X1   g0279(.A1(new_n321), .A2(new_n380), .A3(new_n438), .A4(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT81), .ZN(new_n481));
  INV_X1    g0281(.A(G41), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(KEYINPUT5), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n206), .A2(G45), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT5), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G41), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n487), .A2(KEYINPUT81), .A3(new_n206), .A4(G45), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n482), .A2(KEYINPUT5), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n485), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT82), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n490), .A2(new_n491), .A3(G257), .A4(new_n282), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n276), .A2(new_n488), .A3(new_n489), .A4(new_n485), .ZN(new_n493));
  AND2_X1   g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n490), .A2(G257), .A3(new_n282), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(KEYINPUT82), .ZN(new_n496));
  INV_X1    g0296(.A(G244), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n497), .A2(G1698), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n498), .A2(new_n301), .A3(new_n303), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n293), .A2(G250), .A3(G1698), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n293), .A2(KEYINPUT4), .A3(new_n498), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G33), .A2(G283), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n501), .A2(new_n502), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(G179), .B1(new_n505), .B2(new_n292), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n494), .A2(new_n496), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(KEYINPUT84), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n505), .A2(new_n292), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n496), .A2(new_n509), .A3(new_n493), .A4(new_n492), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n318), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT84), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n494), .A2(new_n512), .A3(new_n496), .A4(new_n506), .ZN(new_n513));
  AND3_X1   g0313(.A1(new_n508), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT83), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n399), .A2(new_n303), .A3(new_n401), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n213), .A2(KEYINPUT7), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n405), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G107), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT6), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n520), .A2(new_n228), .A3(G107), .ZN(new_n521));
  XNOR2_X1  g0321(.A(G97), .B(G107), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n521), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  OAI22_X1  g0323(.A1(new_n523), .A2(new_n213), .B1(new_n294), .B2(new_n391), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n357), .B1(new_n519), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n263), .A2(G97), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n206), .A2(G33), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n263), .A2(new_n528), .A3(new_n214), .A4(new_n260), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n527), .B1(new_n530), .B2(G97), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n515), .B1(new_n526), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(G107), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n534), .B1(new_n403), .B2(new_n405), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n261), .B1(new_n535), .B2(new_n524), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n536), .A2(KEYINPUT83), .A3(new_n531), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n494), .A2(new_n496), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n539), .A2(G190), .A3(new_n509), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n536), .A2(new_n531), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n541), .B1(G200), .B2(new_n510), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n514), .A2(new_n538), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(G116), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n260), .A2(new_n214), .B1(G20), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n504), .B1(new_n228), .B2(G33), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n545), .B1(new_n466), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT20), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n545), .B(KEYINPUT20), .C1(new_n466), .C2(new_n546), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n263), .A2(new_n544), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n530), .B2(new_n544), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n490), .A2(G270), .A3(new_n282), .ZN(new_n555));
  INV_X1    g0355(.A(G303), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n291), .B1(new_n381), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(G257), .A2(G1698), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n296), .A2(G264), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n293), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n555), .A2(new_n493), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n554), .B1(G200), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(new_n375), .B2(new_n562), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n318), .B1(new_n551), .B2(new_n553), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n562), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT21), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(KEYINPUT21), .A2(G169), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n569), .B1(new_n551), .B2(new_n553), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n350), .B1(new_n557), .B2(new_n560), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n555), .A2(new_n571), .A3(new_n493), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n562), .A2(new_n570), .B1(new_n572), .B2(new_n554), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n564), .A2(new_n568), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(KEYINPUT89), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n570), .A2(new_n562), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n572), .A2(new_n554), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT21), .B1(new_n565), .B2(new_n562), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT89), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n580), .A2(new_n581), .A3(new_n564), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n575), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n529), .A2(new_n222), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n463), .A2(new_n465), .A3(G33), .A4(G97), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT19), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n213), .A2(new_n293), .A3(G68), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n328), .A2(KEYINPUT19), .A3(new_n329), .ZN(new_n590));
  NOR2_X1   g0390(.A1(G97), .A2(G107), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n590), .A2(new_n213), .B1(new_n222), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n261), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n468), .A2(new_n264), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT86), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n593), .A2(KEYINPUT86), .A3(new_n594), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n584), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT88), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n484), .A2(G274), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n601), .B1(new_n223), .B2(new_n484), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n221), .A2(new_n296), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n497), .A2(G1698), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI22_X1  g0405(.A1(new_n381), .A2(new_n605), .B1(new_n300), .B2(new_n544), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n282), .A2(new_n602), .B1(new_n606), .B2(new_n292), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n600), .B1(new_n607), .B2(G190), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n484), .A2(new_n223), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n282), .B(new_n609), .C1(G274), .C2(new_n484), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n300), .A2(new_n544), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n603), .A2(new_n604), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n611), .B1(new_n612), .B2(new_n293), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n610), .B1(new_n613), .B2(new_n291), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(G200), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n375), .B2(new_n614), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n608), .B1(new_n616), .B2(new_n600), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n599), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n614), .A2(G169), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT85), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n610), .B(G179), .C1(new_n613), .C2(new_n291), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n620), .B1(new_n619), .B2(new_n621), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g0424(.A(new_n468), .B(KEYINPUT87), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n530), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n593), .A2(KEYINPUT86), .A3(new_n594), .ZN(new_n627));
  AOI21_X1  g0427(.A(KEYINPUT86), .B1(new_n593), .B2(new_n594), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n223), .A2(new_n296), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n229), .A2(G1698), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n293), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(G294), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n633), .B1(new_n300), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n292), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n490), .A2(G264), .A3(new_n282), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n638), .A2(new_n350), .A3(new_n493), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n636), .A2(new_n493), .A3(new_n637), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n318), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n213), .A2(new_n293), .A3(G87), .ZN(new_n642));
  NOR2_X1   g0442(.A1(KEYINPUT90), .A2(KEYINPUT22), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g0444(.A(KEYINPUT91), .B(KEYINPUT23), .Z(new_n645));
  NAND2_X1  g0445(.A1(new_n534), .A2(G20), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n645), .A2(new_n646), .B1(new_n207), .B2(new_n611), .ZN(new_n647));
  XOR2_X1   g0447(.A(KEYINPUT90), .B(KEYINPUT22), .Z(new_n648));
  NAND4_X1  g0448(.A1(new_n648), .A2(G87), .A3(new_n213), .A4(new_n293), .ZN(new_n649));
  NOR2_X1   g0449(.A1(KEYINPUT23), .A2(G107), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n466), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n644), .A2(new_n647), .A3(new_n649), .A4(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(KEYINPUT24), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n645), .A2(new_n646), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n611), .A2(new_n207), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n654), .A2(new_n651), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT24), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n656), .A2(new_n657), .A3(new_n644), .A4(new_n649), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n357), .B1(new_n653), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n264), .A2(new_n534), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n660), .A2(KEYINPUT92), .A3(KEYINPUT25), .ZN(new_n661));
  XNOR2_X1  g0461(.A(KEYINPUT92), .B(KEYINPUT25), .ZN(new_n662));
  OAI221_X1 g0462(.A(new_n661), .B1(new_n529), .B2(new_n534), .C1(new_n660), .C2(new_n662), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n639), .B(new_n641), .C1(new_n659), .C2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n653), .A2(new_n658), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n261), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n640), .A2(new_n373), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n636), .A2(new_n375), .A3(new_n493), .A4(new_n637), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n663), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n666), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  AND4_X1   g0471(.A1(new_n618), .A2(new_n630), .A3(new_n664), .A4(new_n671), .ZN(new_n672));
  AND4_X1   g0472(.A1(new_n480), .A2(new_n543), .A3(new_n583), .A4(new_n672), .ZN(G372));
  INV_X1    g0473(.A(new_n431), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n414), .A2(new_n340), .A3(G179), .ZN(new_n675));
  AOI221_X4 g0475(.A(KEYINPUT18), .B1(new_n674), .B2(new_n675), .C1(new_n408), .C2(new_n420), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n436), .B1(new_n430), .B2(new_n433), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n475), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n379), .A2(new_n679), .B1(new_n356), .B2(new_n371), .ZN(new_n680));
  INV_X1    g0480(.A(new_n429), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n678), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n317), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n683), .A2(new_n320), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n508), .A2(new_n511), .A3(new_n513), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n533), .A2(new_n537), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n629), .A2(new_n624), .B1(new_n599), .B2(new_n617), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(new_n688), .A3(KEYINPUT26), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT26), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n619), .A2(new_n621), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n629), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n614), .A2(new_n375), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n693), .B1(G200), .B2(new_n614), .ZN(new_n694));
  INV_X1    g0494(.A(new_n584), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n694), .B(new_n695), .C1(new_n628), .C2(new_n627), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n508), .A2(new_n511), .A3(new_n513), .A4(new_n541), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n690), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n689), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n692), .A2(new_n696), .A3(new_n671), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT93), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n578), .A2(new_n703), .A3(new_n579), .ZN(new_n704));
  AOI21_X1  g0504(.A(KEYINPUT93), .B1(new_n568), .B2(new_n573), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n664), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n543), .A2(new_n702), .A3(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n700), .A2(new_n707), .A3(new_n692), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n480), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n684), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT94), .ZN(G369));
  INV_X1    g0511(.A(G330), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n568), .A2(new_n573), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n703), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n568), .A2(new_n573), .A3(KEYINPUT93), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n213), .A2(new_n206), .A3(G13), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n716), .A2(KEYINPUT27), .ZN(new_n717));
  OAI21_X1  g0517(.A(G213), .B1(new_n716), .B2(KEYINPUT27), .ZN(new_n718));
  OR2_X1    g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(G343), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n554), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n714), .A2(new_n715), .A3(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT95), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n723), .B1(new_n575), .B2(new_n582), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n724), .A2(new_n725), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  OR2_X1    g0529(.A1(new_n729), .A2(KEYINPUT96), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(KEYINPUT96), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n712), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n721), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n664), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n721), .B1(new_n659), .B2(new_n663), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n671), .A2(new_n664), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n732), .A2(new_n737), .ZN(new_n738));
  AND4_X1   g0538(.A1(new_n713), .A2(new_n671), .A3(new_n664), .A4(new_n733), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n664), .A2(new_n721), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n738), .A2(new_n741), .ZN(G399));
  INV_X1    g0542(.A(new_n210), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G41), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(new_n206), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n591), .A2(new_n222), .A3(new_n544), .ZN(new_n747));
  INV_X1    g0547(.A(new_n744), .ZN(new_n748));
  OAI22_X1  g0548(.A1(new_n746), .A2(new_n747), .B1(new_n216), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT28), .ZN(new_n750));
  INV_X1    g0550(.A(new_n692), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n714), .A2(new_n715), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n701), .B1(new_n752), .B2(new_n664), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n751), .B1(new_n753), .B2(new_n543), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n721), .B1(new_n754), .B2(new_n700), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n755), .A2(KEYINPUT29), .ZN(new_n756));
  NOR3_X1   g0556(.A1(new_n697), .A2(new_n690), .A3(new_n698), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(KEYINPUT99), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT99), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n514), .A2(new_n538), .A3(new_n630), .A4(new_n618), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n759), .B1(new_n760), .B2(new_n690), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n758), .B1(new_n761), .B2(new_n757), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT100), .ZN(new_n763));
  AND3_X1   g0563(.A1(new_n580), .A2(new_n763), .A3(new_n664), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n763), .B1(new_n580), .B2(new_n664), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n764), .A2(new_n765), .A3(new_n701), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n751), .B1(new_n766), .B2(new_n543), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n721), .B1(new_n762), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(KEYINPUT29), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n756), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n562), .A2(new_n350), .A3(new_n614), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(KEYINPUT97), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT97), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n562), .A2(new_n773), .A3(new_n350), .A4(new_n614), .ZN(new_n774));
  NAND4_X1  g0574(.A1(new_n772), .A2(new_n510), .A3(new_n640), .A4(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT30), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n638), .A2(new_n572), .A3(new_n607), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n776), .B1(new_n777), .B2(new_n510), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(KEYINPUT98), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT98), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n775), .A2(new_n778), .A3(new_n781), .ZN(new_n782));
  OR3_X1    g0582(.A1(new_n777), .A2(new_n776), .A3(new_n510), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n780), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n784), .A2(KEYINPUT31), .A3(new_n721), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n583), .A2(new_n672), .A3(new_n543), .A4(new_n733), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n783), .A2(new_n778), .A3(new_n775), .ZN(new_n787));
  AND2_X1   g0587(.A1(new_n787), .A2(new_n721), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n785), .B(new_n786), .C1(KEYINPUT31), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G330), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n770), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n750), .B1(new_n792), .B2(G1), .ZN(G364));
  INV_X1    g0593(.A(new_n732), .ZN(new_n794));
  INV_X1    g0594(.A(G13), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n466), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G45), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n745), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n730), .A2(new_n712), .A3(new_n731), .ZN(new_n799));
  AND3_X1   g0599(.A1(new_n794), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n743), .A2(new_n381), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n801), .A2(G355), .B1(new_n544), .B2(new_n743), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n743), .A2(new_n293), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(G45), .B2(new_n216), .ZN(new_n804));
  INV_X1    g0604(.A(G45), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n249), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n802), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(G13), .A2(G33), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(G20), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n214), .B1(G20), .B2(new_n318), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n798), .B1(new_n807), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(G179), .A2(G190), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n466), .A2(G200), .A3(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(new_n534), .ZN(new_n816));
  NOR4_X1   g0616(.A1(new_n207), .A2(new_n375), .A3(new_n373), .A4(G179), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n381), .B(new_n816), .C1(G87), .C2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n375), .A2(G200), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n213), .B1(new_n350), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n818), .B1(new_n228), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n466), .A2(G179), .ZN(new_n822));
  NOR3_X1   g0622(.A1(new_n822), .A2(G190), .A3(G200), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT102), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n823), .A2(new_n824), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(new_n294), .ZN(new_n829));
  INV_X1    g0629(.A(new_n822), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n819), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT101), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n821), .B(new_n829), .C1(G58), .C2(new_n832), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n466), .A2(new_n373), .A3(new_n814), .ZN(new_n834));
  XOR2_X1   g0634(.A(KEYINPUT103), .B(KEYINPUT32), .Z(new_n835));
  NOR3_X1   g0635(.A1(new_n834), .A2(new_n390), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n835), .B1(new_n834), .B2(new_n390), .ZN(new_n837));
  NOR3_X1   g0637(.A1(new_n822), .A2(G190), .A3(new_n373), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n837), .B1(new_n839), .B2(new_n220), .ZN(new_n840));
  NOR3_X1   g0640(.A1(new_n822), .A2(new_n375), .A3(new_n373), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n836), .B(new_n840), .C1(G50), .C2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n820), .ZN(new_n843));
  AOI22_X1  g0643(.A1(G311), .A2(new_n823), .B1(new_n843), .B2(G294), .ZN(new_n844));
  INV_X1    g0644(.A(G326), .ZN(new_n845));
  INV_X1    g0645(.A(new_n841), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n847), .B(KEYINPUT104), .Z(new_n848));
  INV_X1    g0648(.A(new_n815), .ZN(new_n849));
  INV_X1    g0649(.A(new_n834), .ZN(new_n850));
  AOI22_X1  g0650(.A1(G283), .A2(new_n849), .B1(new_n850), .B2(G329), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n293), .B1(new_n817), .B2(G303), .ZN(new_n852));
  INV_X1    g0652(.A(G322), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n851), .B(new_n852), .C1(new_n853), .C2(new_n831), .ZN(new_n854));
  XNOR2_X1  g0654(.A(KEYINPUT105), .B(KEYINPUT33), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(G317), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n854), .B1(new_n838), .B2(new_n856), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n833), .A2(new_n842), .B1(new_n848), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n811), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n813), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(new_n729), .B2(new_n810), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n800), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(G396));
  INV_X1    g0663(.A(new_n798), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n474), .A2(new_n721), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n475), .A2(new_n478), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(KEYINPUT108), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT108), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n475), .A2(new_n478), .A3(new_n868), .A4(new_n865), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n452), .A2(new_n462), .A3(new_n474), .A4(new_n721), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n871), .B(KEYINPUT109), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n755), .B(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n864), .B1(new_n874), .B2(new_n790), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(new_n790), .B2(new_n874), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n811), .A2(new_n808), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n798), .B1(new_n294), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(G283), .ZN(new_n879));
  OAI22_X1  g0679(.A1(new_n828), .A2(new_n544), .B1(new_n879), .B2(new_n839), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT106), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n880), .A2(new_n881), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n815), .A2(new_n222), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(G311), .B2(new_n850), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n634), .B2(new_n831), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n293), .B1(new_n817), .B2(G107), .ZN(new_n887));
  OAI221_X1 g0687(.A(new_n887), .B1(new_n820), .B2(new_n228), .C1(new_n846), .C2(new_n556), .ZN(new_n888));
  NOR4_X1   g0688(.A1(new_n882), .A2(new_n883), .A3(new_n886), .A4(new_n888), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n843), .A2(G58), .B1(new_n849), .B2(G68), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n381), .B1(new_n817), .B2(G50), .ZN(new_n891));
  INV_X1    g0691(.A(G132), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n890), .B(new_n891), .C1(new_n892), .C2(new_n834), .ZN(new_n893));
  XOR2_X1   g0693(.A(new_n893), .B(KEYINPUT107), .Z(new_n894));
  INV_X1    g0694(.A(KEYINPUT34), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n832), .A2(G143), .ZN(new_n896));
  AOI22_X1  g0696(.A1(G137), .A2(new_n841), .B1(new_n838), .B2(G150), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n896), .B(new_n897), .C1(new_n390), .C2(new_n828), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n894), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  OR2_X1    g0699(.A1(new_n898), .A2(new_n895), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n889), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI221_X1 g0701(.A(new_n878), .B1(new_n901), .B2(new_n859), .C1(new_n873), .C2(new_n809), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n876), .A2(new_n902), .ZN(G384));
  NOR2_X1   g0703(.A1(new_n796), .A2(new_n206), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT38), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n397), .A2(new_n261), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT16), .B1(new_n387), .B2(new_n396), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n420), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT110), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI211_X1 g0710(.A(KEYINPUT110), .B(new_n420), .C1(new_n906), .C2(new_n907), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI211_X1 g0712(.A(new_n719), .B(new_n912), .C1(new_n678), .C2(new_n429), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n432), .A2(new_n719), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n910), .A2(new_n914), .A3(new_n911), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n421), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT111), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT37), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n421), .A2(new_n918), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n432), .A2(new_n719), .B1(new_n408), .B2(new_n420), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n917), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n914), .A2(new_n430), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n922), .A2(KEYINPUT111), .A3(new_n918), .A4(new_n421), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n916), .A2(KEYINPUT37), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n905), .B1(new_n913), .B2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n719), .ZN(new_n926));
  INV_X1    g0726(.A(new_n912), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n438), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n921), .A2(new_n923), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n918), .B1(new_n915), .B2(new_n421), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n928), .B(KEYINPUT38), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT40), .B1(new_n925), .B2(new_n932), .ZN(new_n933));
  AND3_X1   g0733(.A1(new_n787), .A2(KEYINPUT31), .A3(new_n721), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT31), .B1(new_n787), .B2(new_n721), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n786), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n371), .A2(new_n721), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n372), .A2(new_n379), .A3(new_n938), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n371), .B(new_n721), .C1(new_n378), .C2(new_n356), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AND3_X1   g0741(.A1(new_n937), .A2(new_n941), .A3(new_n873), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n933), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n937), .A2(new_n941), .A3(new_n873), .ZN(new_n944));
  AND3_X1   g0744(.A1(new_n438), .A2(new_n430), .A3(new_n926), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n421), .A2(KEYINPUT112), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n946), .A2(new_n918), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n922), .A2(KEYINPUT112), .A3(new_n421), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n921), .A2(new_n923), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n905), .B1(new_n945), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n944), .B1(new_n932), .B2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT40), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n943), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n480), .A2(new_n937), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n712), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n954), .B2(new_n953), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT39), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n913), .A2(new_n924), .A3(new_n905), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n947), .A2(new_n948), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n929), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n438), .A2(new_n430), .A3(new_n926), .ZN(new_n961));
  AOI21_X1  g0761(.A(KEYINPUT38), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n957), .B1(new_n958), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n372), .A2(new_n721), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n925), .A2(KEYINPUT39), .A3(new_n932), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n678), .A2(new_n926), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n939), .A2(new_n940), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n873), .A2(new_n708), .A3(new_n733), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n475), .A2(new_n721), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n968), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n925), .A2(new_n932), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n967), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n966), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n756), .A2(new_n480), .A3(new_n769), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n684), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n975), .B(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n904), .B1(new_n956), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n978), .B2(new_n956), .ZN(new_n980));
  INV_X1    g0780(.A(new_n523), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n981), .A2(KEYINPUT35), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(KEYINPUT35), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n982), .A2(G116), .A3(new_n215), .A4(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT36), .ZN(new_n985));
  OAI21_X1  g0785(.A(G77), .B1(new_n226), .B2(new_n220), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n245), .B1(new_n986), .B2(new_n216), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n987), .A2(G1), .A3(new_n795), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n980), .A2(new_n985), .A3(new_n988), .ZN(G367));
  INV_X1    g0789(.A(new_n828), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(G50), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n849), .A2(G77), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n381), .B1(new_n817), .B2(G58), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(new_n839), .C2(new_n390), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n994), .B1(G143), .B2(new_n841), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n843), .A2(G68), .ZN(new_n996));
  INV_X1    g0796(.A(new_n831), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n997), .A2(G150), .B1(G137), .B2(new_n850), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n991), .A2(new_n995), .A3(new_n996), .A4(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n832), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n1000), .A2(new_n556), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n828), .A2(new_n879), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n815), .A2(new_n228), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(G317), .B2(new_n850), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n534), .B2(new_n820), .ZN(new_n1005));
  OR3_X1    g0805(.A1(new_n1001), .A2(new_n1002), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n838), .A2(G294), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n841), .A2(G311), .ZN(new_n1008));
  AOI21_X1  g0808(.A(KEYINPUT46), .B1(new_n817), .B2(G116), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1009), .A2(new_n293), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n817), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1007), .A2(new_n1008), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n999), .B1(new_n1006), .B2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT116), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT47), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n811), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n599), .A2(new_n733), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n751), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n697), .B2(new_n1017), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n810), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n803), .A2(new_n240), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n210), .A2(new_n468), .ZN(new_n1023));
  NOR3_X1   g0823(.A1(new_n1023), .A2(new_n810), .A3(new_n811), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n798), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1016), .A2(new_n1021), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n541), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n543), .B1(new_n1027), .B2(new_n733), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n514), .A2(new_n541), .A3(new_n721), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n739), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT42), .Z(new_n1032));
  INV_X1    g0832(.A(new_n1030), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1033), .A2(new_n664), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n733), .B1(new_n1034), .B2(new_n687), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT43), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1020), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(KEYINPUT113), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1019), .A2(KEYINPUT43), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1036), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  OR3_X1    g0842(.A1(new_n1036), .A2(KEYINPUT113), .A3(new_n1038), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n738), .A2(new_n1033), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(KEYINPUT114), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT114), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1042), .A2(new_n1048), .A3(new_n1045), .A4(new_n1043), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1047), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n797), .A2(G1), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1030), .A2(new_n741), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT44), .Z(new_n1054));
  NAND2_X1  g0854(.A1(new_n1030), .A2(new_n741), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT45), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n738), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n732), .B(new_n737), .C1(new_n1054), .C2(new_n1056), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n737), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n713), .A2(new_n733), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n739), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n732), .A2(new_n1064), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n712), .B(new_n1063), .C1(new_n730), .C2(new_n731), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n792), .B1(new_n1060), .B2(new_n1067), .ZN(new_n1068));
  XOR2_X1   g0868(.A(KEYINPUT115), .B(KEYINPUT41), .Z(new_n1069));
  XNOR2_X1  g0869(.A(new_n744), .B(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1052), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1026), .B1(new_n1051), .B2(new_n1071), .ZN(G387));
  INV_X1    g0872(.A(KEYINPUT117), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1052), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1073), .B1(new_n1067), .B2(new_n1074), .ZN(new_n1075));
  OAI211_X1 g0875(.A(KEYINPUT117), .B(new_n1052), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n990), .A2(G303), .B1(G317), .B2(new_n832), .ZN(new_n1077));
  OR2_X1    g0877(.A1(new_n1077), .A2(KEYINPUT118), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(KEYINPUT118), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G311), .A2(new_n838), .B1(new_n841), .B2(G322), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT48), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n843), .A2(G283), .B1(new_n817), .B2(G294), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT49), .Z(new_n1087));
  OAI221_X1 g0887(.A(new_n381), .B1(new_n834), .B2(new_n845), .C1(new_n544), .C2(new_n815), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n823), .A2(G68), .B1(G150), .B2(new_n850), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n625), .A2(new_n843), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1089), .B(new_n1090), .C1(new_n202), .C2(new_n831), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n381), .B(new_n1003), .C1(G77), .C2(new_n817), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1092), .B1(new_n390), .B2(new_n846), .C1(new_n419), .C2(new_n839), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n1087), .A2(new_n1088), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n811), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1061), .A2(new_n810), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n801), .A2(new_n747), .B1(new_n534), .B2(new_n743), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n237), .A2(new_n805), .ZN(new_n1098));
  AOI211_X1 g0898(.A(G45), .B(new_n747), .C1(G68), .C2(G77), .ZN(new_n1099));
  AOI21_X1  g0899(.A(KEYINPUT50), .B1(new_n255), .B2(new_n202), .ZN(new_n1100));
  AND3_X1   g0900(.A1(new_n255), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1099), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n803), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1097), .B1(new_n1098), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n798), .B1(new_n1104), .B2(new_n812), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n1096), .A2(new_n1105), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1075), .A2(new_n1076), .B1(new_n1095), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT119), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n792), .B1(new_n1066), .B2(new_n1065), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1067), .A2(new_n791), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1109), .A2(new_n1110), .A3(new_n744), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1107), .A2(new_n1108), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1108), .B1(new_n1107), .B2(new_n1111), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(G393));
  INV_X1    g0916(.A(new_n1060), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1109), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n748), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n1118), .B2(new_n1117), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1117), .A2(new_n1052), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1033), .A2(new_n810), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n997), .A2(G311), .B1(G317), .B2(new_n841), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1123), .B(KEYINPUT52), .Z(new_n1124));
  OAI22_X1  g0924(.A1(new_n820), .A2(new_n544), .B1(new_n834), .B2(new_n853), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(G294), .B2(new_n823), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n817), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n381), .B1(new_n1127), .B2(new_n879), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n816), .B(new_n1128), .C1(G303), .C2(new_n838), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1124), .A2(new_n1126), .A3(new_n1129), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n381), .B(new_n884), .C1(G68), .C2(new_n817), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n843), .A2(G77), .B1(new_n850), .B2(G143), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n1133), .B1(new_n202), .B2(new_n839), .C1(new_n419), .C2(new_n828), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n997), .A2(G159), .B1(G150), .B2(new_n841), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT51), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1130), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n811), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n803), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n812), .B1(new_n228), .B2(new_n210), .C1(new_n1139), .C2(new_n244), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1122), .A2(new_n864), .A3(new_n1138), .A4(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1120), .A2(new_n1121), .A3(new_n1141), .ZN(G390));
  INV_X1    g0942(.A(new_n873), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n968), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n712), .B1(new_n936), .B2(new_n786), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n925), .A2(KEYINPUT39), .A3(new_n932), .ZN(new_n1147));
  AOI21_X1  g0947(.A(KEYINPUT39), .B1(new_n950), .B2(new_n932), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n1147), .A2(new_n1148), .B1(new_n964), .B2(new_n972), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n964), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n950), .A2(new_n932), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n970), .B1(new_n768), .B2(new_n873), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1150), .B(new_n1151), .C1(new_n1152), .C2(new_n968), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1146), .B1(new_n1149), .B2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n789), .A2(G330), .A3(new_n873), .ZN(new_n1155));
  OR2_X1    g0955(.A1(new_n1155), .A2(new_n968), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1149), .A2(new_n1153), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(KEYINPUT120), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1155), .A2(new_n968), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n963), .A2(new_n965), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n970), .B1(new_n755), .B2(new_n873), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1150), .B1(new_n1161), .B2(new_n968), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1159), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT120), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1163), .A2(new_n1164), .A3(new_n1153), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1154), .B1(new_n1158), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n1052), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1160), .A2(new_n808), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n293), .B1(new_n817), .B2(G87), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1169), .B1(new_n220), .B2(new_n815), .C1(new_n839), .C2(new_n534), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n843), .A2(G77), .B1(new_n850), .B2(G294), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1171), .B1(new_n544), .B2(new_n831), .C1(new_n828), .C2(new_n228), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1170), .B(new_n1172), .C1(G283), .C2(new_n841), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n817), .A2(G150), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1174), .A2(KEYINPUT53), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n381), .B1(new_n1174), .B2(KEYINPUT53), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(G128), .ZN(new_n1178));
  INV_X1    g0978(.A(G137), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1177), .B1(new_n1178), .B2(new_n846), .C1(new_n1179), .C2(new_n839), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(KEYINPUT54), .B(G143), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n828), .A2(new_n1181), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(G50), .A2(new_n849), .B1(new_n850), .B2(G125), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1183), .B1(new_n892), .B2(new_n831), .C1(new_n390), .C2(new_n820), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n1180), .A2(new_n1182), .A3(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1173), .A2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1186), .A2(new_n859), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n798), .B(new_n1187), .C1(new_n419), .C2(new_n877), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1168), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n480), .A2(new_n1145), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n976), .A2(new_n684), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1155), .A2(new_n968), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1146), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1161), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n937), .A2(G330), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1196), .A2(KEYINPUT121), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT121), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n873), .B1(new_n1145), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n968), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1200), .A2(new_n1152), .A3(new_n1156), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1191), .B1(new_n1195), .B2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n744), .B1(new_n1166), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1154), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1164), .B1(new_n1163), .B2(new_n1153), .ZN(new_n1205));
  AND4_X1   g1005(.A1(new_n1164), .A2(new_n1149), .A3(new_n1153), .A4(new_n1156), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1204), .B(new_n1202), .C1(new_n1205), .C2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1167), .B(new_n1189), .C1(new_n1203), .C2(new_n1208), .ZN(G378));
  NAND2_X1  g1009(.A1(new_n268), .A2(new_n926), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n321), .B(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1214));
  AND2_X1   g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1151), .A2(new_n942), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n1216), .A2(KEYINPUT40), .B1(new_n933), .B2(new_n942), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(new_n1215), .A2(new_n1217), .A3(new_n712), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n953), .B2(G330), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n975), .B1(new_n1218), .B2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1215), .B1(new_n1217), .B2(new_n712), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n953), .A2(new_n1219), .A3(G330), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n975), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1221), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1215), .A2(new_n808), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n381), .A2(new_n482), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(G77), .B2(new_n817), .ZN(new_n1229));
  AND2_X1   g1029(.A1(new_n996), .A2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n228), .B2(new_n839), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n997), .A2(G107), .B1(new_n625), .B2(new_n823), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1232), .B1(new_n226), .B2(new_n815), .C1(new_n879), .C2(new_n834), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1231), .B(new_n1233), .C1(G116), .C2(new_n841), .ZN(new_n1234));
  AOI21_X1  g1034(.A(G50), .B1(new_n300), .B2(new_n482), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1234), .A2(KEYINPUT58), .B1(new_n1228), .B2(new_n1235), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(G137), .A2(new_n823), .B1(new_n843), .B2(G150), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n892), .B2(new_n839), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n831), .A2(new_n1178), .B1(new_n1127), .B2(new_n1181), .ZN(new_n1239));
  XOR2_X1   g1039(.A(new_n1239), .B(KEYINPUT122), .Z(new_n1240));
  AOI211_X1 g1040(.A(new_n1238), .B(new_n1240), .C1(G125), .C2(new_n841), .ZN(new_n1241));
  XOR2_X1   g1041(.A(new_n1241), .B(KEYINPUT123), .Z(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1243), .A2(KEYINPUT59), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n300), .B(new_n482), .C1(new_n815), .C2(new_n390), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(G124), .B2(new_n850), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT59), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1246), .B1(new_n1242), .B2(new_n1247), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n1236), .B1(KEYINPUT58), .B2(new_n1234), .C1(new_n1244), .C2(new_n1248), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1249), .A2(new_n811), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n798), .B(new_n1250), .C1(new_n202), .C2(new_n877), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n1226), .A2(new_n1052), .B1(new_n1227), .B2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1191), .B1(new_n1166), .B2(new_n1202), .ZN(new_n1253));
  AND3_X1   g1053(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1224), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1255));
  OAI21_X1  g1055(.A(KEYINPUT57), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n744), .B1(new_n1253), .B2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1191), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1207), .A2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT57), .B1(new_n1259), .B2(new_n1226), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1252), .B1(new_n1257), .B2(new_n1260), .ZN(G375));
  AND2_X1   g1061(.A1(new_n1201), .A2(new_n1195), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1191), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1202), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1263), .A2(new_n1264), .A3(new_n1070), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1201), .A2(new_n1195), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n1052), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n798), .B1(new_n220), .B2(new_n877), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n828), .A2(new_n534), .B1(new_n544), .B2(new_n839), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(new_n1269), .B(KEYINPUT124), .ZN(new_n1270));
  OAI221_X1 g1070(.A(new_n1090), .B1(new_n556), .B2(new_n834), .C1(new_n879), .C2(new_n831), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n293), .B1(new_n817), .B2(G97), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n992), .B(new_n1272), .C1(new_n846), .C2(new_n634), .ZN(new_n1273));
  OR3_X1    g1073(.A1(new_n1270), .A2(new_n1271), .A3(new_n1273), .ZN(new_n1274));
  OAI221_X1 g1074(.A(new_n293), .B1(new_n815), .B2(new_n226), .C1(new_n1127), .C2(new_n390), .ZN(new_n1275));
  OAI22_X1  g1075(.A1(new_n892), .A2(new_n846), .B1(new_n839), .B2(new_n1181), .ZN(new_n1276));
  AOI211_X1 g1076(.A(new_n1275), .B(new_n1276), .C1(G128), .C2(new_n850), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(G150), .A2(new_n823), .B1(new_n843), .B2(G50), .ZN(new_n1278));
  XOR2_X1   g1078(.A(new_n1278), .B(KEYINPUT125), .Z(new_n1279));
  OAI211_X1 g1079(.A(new_n1277), .B(new_n1279), .C1(new_n1179), .C2(new_n1000), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1274), .A2(new_n1280), .ZN(new_n1281));
  OAI221_X1 g1081(.A(new_n1268), .B1(new_n1281), .B2(new_n859), .C1(new_n809), .C2(new_n941), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1265), .A2(new_n1267), .A3(new_n1282), .ZN(G381));
  NOR4_X1   g1083(.A1(G387), .A2(G384), .A3(G390), .A4(G381), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1204), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1189), .B1(new_n1285), .B2(new_n1074), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n748), .B1(new_n1285), .B2(new_n1264), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1286), .B1(new_n1207), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(G375), .ZN(new_n1289));
  NOR3_X1   g1089(.A1(new_n1113), .A2(new_n1114), .A3(G396), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1284), .A2(new_n1288), .A3(new_n1289), .A4(new_n1290), .ZN(G407));
  NAND2_X1  g1091(.A1(new_n720), .A2(G213), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1289), .A2(new_n1288), .A3(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(G407), .A2(G213), .A3(new_n1294), .ZN(G409));
  OAI211_X1 g1095(.A(G378), .B(new_n1252), .C1(new_n1257), .C2(new_n1260), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1259), .A2(new_n1070), .A3(new_n1226), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1226), .A2(new_n1052), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1251), .A2(new_n1227), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1288), .B1(new_n1297), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1296), .A2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1292), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT60), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1263), .B1(new_n1304), .B2(new_n1202), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1262), .A2(KEYINPUT60), .A3(new_n1191), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1305), .A2(new_n744), .A3(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n876), .A2(KEYINPUT126), .A3(new_n902), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1308), .A2(new_n1267), .A3(new_n1282), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT126), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(G384), .A2(new_n1310), .ZN(new_n1311));
  AND3_X1   g1111(.A1(new_n1307), .A2(new_n1309), .A3(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1311), .B1(new_n1307), .B2(new_n1309), .ZN(new_n1313));
  INV_X1    g1113(.A(G2897), .ZN(new_n1314));
  OAI22_X1  g1114(.A1(new_n1312), .A2(new_n1313), .B1(new_n1314), .B2(new_n1292), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1307), .A2(new_n1309), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1311), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1307), .A2(new_n1309), .A3(new_n1311), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1292), .A2(new_n1314), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1318), .A2(new_n1319), .A3(new_n1320), .ZN(new_n1321));
  AND2_X1   g1121(.A1(new_n1315), .A2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(KEYINPUT61), .B1(new_n1303), .B2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT63), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1324), .B1(new_n1303), .B2(new_n1325), .ZN(new_n1326));
  OAI21_X1  g1126(.A(G396), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(KEYINPUT119), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1329), .A2(new_n862), .A3(new_n1112), .ZN(new_n1330));
  AND3_X1   g1130(.A1(new_n1327), .A2(new_n1330), .A3(G390), .ZN(new_n1331));
  AOI21_X1  g1131(.A(G390), .B1(new_n1327), .B2(new_n1330), .ZN(new_n1332));
  NOR3_X1   g1132(.A1(new_n1331), .A2(new_n1332), .A3(G387), .ZN(new_n1333));
  INV_X1    g1133(.A(G387), .ZN(new_n1334));
  INV_X1    g1134(.A(G390), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n862), .B1(new_n1329), .B2(new_n1112), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1335), .B1(new_n1290), .B2(new_n1336), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1327), .A2(new_n1330), .A3(G390), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1334), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1333), .A2(new_n1339), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1293), .B1(new_n1296), .B2(new_n1301), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1325), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1341), .A2(KEYINPUT63), .A3(new_n1342), .ZN(new_n1343));
  NAND4_X1  g1143(.A1(new_n1323), .A2(new_n1326), .A3(new_n1340), .A4(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT62), .ZN(new_n1345));
  AND3_X1   g1145(.A1(new_n1341), .A2(new_n1345), .A3(new_n1342), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT61), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1315), .A2(new_n1321), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1347), .B1(new_n1341), .B2(new_n1348), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1345), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1350));
  NOR3_X1   g1150(.A1(new_n1346), .A2(new_n1349), .A3(new_n1350), .ZN(new_n1351));
  OAI21_X1  g1151(.A(KEYINPUT127), .B1(new_n1333), .B2(new_n1339), .ZN(new_n1352));
  OAI21_X1  g1152(.A(G387), .B1(new_n1331), .B2(new_n1332), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1337), .A2(new_n1334), .A3(new_n1338), .ZN(new_n1354));
  INV_X1    g1154(.A(KEYINPUT127), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1353), .A2(new_n1354), .A3(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1352), .A2(new_n1356), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1344), .B1(new_n1351), .B2(new_n1357), .ZN(G405));
  NAND2_X1  g1158(.A1(G375), .A2(new_n1288), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1359), .A2(new_n1296), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1360), .A2(new_n1325), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1342), .A2(new_n1359), .A3(new_n1296), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1361), .A2(new_n1362), .ZN(new_n1363));
  XNOR2_X1  g1163(.A(new_n1363), .B(new_n1340), .ZN(G402));
endmodule


