//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 1 0 0 1 1 0 0 0 0 1 0 0 1 0 1 1 1 0 1 0 0 0 1 1 0 1 1 0 0 1 0 0 1 1 0 0 0 1 1 0 0 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009;
  INV_X1    g000(.A(KEYINPUT73), .ZN(new_n187));
  NOR2_X1   g001(.A1(G472), .A2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  NOR2_X1   g003(.A1(G237), .A2(G953), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G210), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n191), .B(KEYINPUT27), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT26), .B(G101), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT11), .ZN(new_n195));
  INV_X1    g009(.A(G134), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n195), .B1(new_n196), .B2(G137), .ZN(new_n197));
  INV_X1    g011(.A(G137), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(KEYINPUT11), .A3(G134), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n196), .A2(G137), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n197), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G131), .ZN(new_n202));
  INV_X1    g016(.A(G131), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n197), .A2(new_n199), .A3(new_n203), .A4(new_n200), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G143), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(KEYINPUT0), .A2(G128), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g026(.A1(KEYINPUT0), .A2(G128), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n210), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(G143), .B(G146), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(new_n211), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n205), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT1), .ZN(new_n219));
  AND4_X1   g033(.A1(new_n219), .A2(new_n207), .A3(new_n209), .A4(G128), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT1), .B1(new_n208), .B2(G146), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT65), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n223), .B(KEYINPUT1), .C1(new_n208), .C2(G146), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n222), .A2(G128), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n220), .B1(new_n225), .B2(new_n210), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT64), .ZN(new_n227));
  XNOR2_X1  g041(.A(G134), .B(G137), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n227), .B1(new_n228), .B2(new_n203), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n196), .A2(G137), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n198), .A2(G134), .ZN(new_n231));
  OAI211_X1 g045(.A(KEYINPUT64), .B(G131), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n229), .A2(new_n204), .A3(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n218), .B1(new_n226), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n235));
  INV_X1    g049(.A(G116), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n235), .B1(new_n236), .B2(G119), .ZN(new_n237));
  INV_X1    g051(.A(G119), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(KEYINPUT67), .A3(G116), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n236), .A2(G119), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n237), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G113), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT2), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT2), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G113), .ZN(new_n245));
  AND2_X1   g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n241), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n243), .A2(new_n245), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n248), .A2(new_n237), .A3(new_n239), .A4(new_n240), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n247), .A2(new_n249), .A3(KEYINPUT68), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n194), .B1(new_n234), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT31), .ZN(new_n257));
  AOI22_X1  g071(.A1(new_n202), .A2(new_n204), .B1(new_n214), .B2(new_n216), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n229), .A2(new_n204), .A3(new_n232), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n224), .A2(G128), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n223), .B1(new_n207), .B2(KEYINPUT1), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n210), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n220), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n258), .B1(new_n265), .B2(KEYINPUT66), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT66), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n259), .A2(new_n264), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT30), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n218), .B(KEYINPUT30), .C1(new_n226), .C2(new_n233), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n254), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n256), .B(new_n257), .C1(new_n269), .C2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT70), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(KEYINPUT66), .B1(new_n226), .B2(new_n233), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(new_n268), .A3(new_n218), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT30), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AND3_X1   g092(.A1(new_n247), .A2(new_n249), .A3(KEYINPUT68), .ZN(new_n279));
  AOI21_X1  g093(.A(KEYINPUT68), .B1(new_n247), .B2(new_n249), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n258), .B1(new_n264), .B2(new_n259), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n281), .B1(new_n282), .B2(KEYINPUT30), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n255), .B1(new_n278), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(KEYINPUT70), .A3(new_n257), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT69), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n286), .B1(new_n284), .B2(new_n257), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n271), .B1(new_n277), .B2(new_n276), .ZN(new_n288));
  OAI211_X1 g102(.A(KEYINPUT69), .B(KEYINPUT31), .C1(new_n288), .C2(new_n255), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n274), .A2(new_n285), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n194), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT72), .ZN(new_n292));
  AOI211_X1 g106(.A(new_n292), .B(KEYINPUT28), .C1(new_n282), .C2(new_n281), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n265), .A2(new_n252), .A3(new_n253), .A4(new_n218), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT28), .ZN(new_n295));
  AOI21_X1  g109(.A(KEYINPUT72), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n276), .A2(new_n254), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n295), .B1(new_n298), .B2(new_n294), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n297), .B1(new_n299), .B2(KEYINPUT71), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT71), .ZN(new_n301));
  AOI211_X1 g115(.A(new_n301), .B(new_n295), .C1(new_n298), .C2(new_n294), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n291), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n189), .B1(new_n290), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n187), .B1(new_n304), .B2(KEYINPUT32), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n274), .A2(new_n285), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n287), .A2(new_n289), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n295), .B1(new_n234), .B2(new_n254), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n292), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n294), .A2(KEYINPUT72), .A3(new_n295), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n281), .B1(new_n266), .B2(new_n268), .ZN(new_n313));
  INV_X1    g127(.A(new_n294), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT28), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n312), .B1(new_n315), .B2(new_n301), .ZN(new_n316));
  INV_X1    g130(.A(new_n302), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n194), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n188), .B1(new_n308), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT32), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(KEYINPUT73), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n304), .A2(KEYINPUT32), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n194), .B1(new_n300), .B2(new_n302), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n288), .A2(new_n314), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n291), .ZN(new_n325));
  AOI21_X1  g139(.A(KEYINPUT29), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G902), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n234), .A2(new_n254), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(new_n329), .A3(new_n294), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n234), .A2(KEYINPUT74), .A3(new_n254), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n297), .B1(new_n295), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n194), .A2(KEYINPUT29), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n327), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(G472), .B1(new_n326), .B2(new_n335), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n305), .A2(new_n321), .A3(new_n322), .A4(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G217), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n338), .B1(G234), .B2(new_n327), .ZN(new_n339));
  OAI21_X1  g153(.A(KEYINPUT75), .B1(new_n238), .B2(G128), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT75), .ZN(new_n341));
  INV_X1    g155(.A(G128), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n341), .A2(new_n342), .A3(G119), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n238), .A2(G128), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n340), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT24), .B(G110), .ZN(new_n346));
  AND3_X1   g160(.A1(new_n345), .A2(KEYINPUT77), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(KEYINPUT77), .B1(new_n345), .B2(new_n346), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT23), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n349), .B1(new_n238), .B2(G128), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n342), .A2(KEYINPUT23), .A3(G119), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n344), .A3(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n352), .A2(G110), .ZN(new_n353));
  NOR3_X1   g167(.A1(new_n347), .A2(new_n348), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G140), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G125), .ZN(new_n356));
  INV_X1    g170(.A(G125), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G140), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n356), .A2(new_n358), .A3(KEYINPUT16), .ZN(new_n359));
  OR3_X1    g173(.A1(new_n357), .A2(KEYINPUT16), .A3(G140), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n360), .A3(G146), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT78), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT78), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n359), .A2(new_n360), .A3(new_n363), .A4(G146), .ZN(new_n364));
  XNOR2_X1  g178(.A(G125), .B(G140), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n206), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n362), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n354), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n352), .A2(G110), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n369), .B1(new_n346), .B2(new_n345), .ZN(new_n370));
  AOI21_X1  g184(.A(G146), .B1(new_n359), .B2(new_n360), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT76), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n371), .B1(new_n372), .B2(new_n361), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n359), .A2(new_n360), .A3(KEYINPUT76), .A4(G146), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n370), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT79), .B1(new_n368), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n361), .A2(new_n372), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n359), .A2(new_n360), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n377), .B(new_n374), .C1(G146), .C2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n370), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT79), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n381), .B(new_n382), .C1(new_n354), .C2(new_n367), .ZN(new_n383));
  XNOR2_X1  g197(.A(KEYINPUT22), .B(G137), .ZN(new_n384));
  INV_X1    g198(.A(G953), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n385), .A2(G221), .A3(G234), .ZN(new_n386));
  XOR2_X1   g200(.A(new_n384), .B(new_n386), .Z(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n376), .A2(new_n383), .A3(new_n388), .ZN(new_n389));
  OAI211_X1 g203(.A(KEYINPUT79), .B(new_n387), .C1(new_n368), .C2(new_n375), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(KEYINPUT25), .B1(new_n391), .B2(new_n327), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT25), .ZN(new_n393));
  AOI211_X1 g207(.A(new_n393), .B(G902), .C1(new_n389), .C2(new_n390), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n339), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n339), .A2(G902), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n391), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G221), .ZN(new_n400));
  XNOR2_X1  g214(.A(KEYINPUT9), .B(G234), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n400), .B1(new_n402), .B2(new_n327), .ZN(new_n403));
  INV_X1    g217(.A(G469), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n404), .A2(new_n327), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n385), .A2(G227), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n406), .B(KEYINPUT80), .ZN(new_n407));
  XNOR2_X1  g221(.A(G110), .B(G140), .ZN(new_n408));
  XOR2_X1   g222(.A(new_n407), .B(new_n408), .Z(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT84), .ZN(new_n411));
  INV_X1    g225(.A(G104), .ZN(new_n412));
  OAI21_X1  g226(.A(KEYINPUT3), .B1(new_n412), .B2(G107), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT3), .ZN(new_n414));
  INV_X1    g228(.A(G107), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(new_n415), .A3(G104), .ZN(new_n416));
  INV_X1    g230(.A(G101), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n412), .A2(G107), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n413), .A2(new_n416), .A3(new_n417), .A4(new_n418), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n412), .A2(G107), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n415), .A2(G104), .ZN(new_n421));
  OAI21_X1  g235(.A(G101), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  OAI211_X1 g237(.A(KEYINPUT83), .B(KEYINPUT1), .C1(new_n208), .C2(G146), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G128), .ZN(new_n425));
  AOI21_X1  g239(.A(KEYINPUT83), .B1(new_n207), .B2(KEYINPUT1), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n210), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n423), .B1(new_n427), .B2(new_n263), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n411), .B1(new_n428), .B2(KEYINPUT10), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT10), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT83), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n221), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(G128), .A3(new_n424), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n220), .B1(new_n433), .B2(new_n210), .ZN(new_n434));
  OAI211_X1 g248(.A(KEYINPUT84), .B(new_n430), .C1(new_n434), .C2(new_n423), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n429), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n419), .A2(new_n422), .A3(KEYINPUT10), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n226), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n413), .A2(new_n416), .A3(new_n418), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT82), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n413), .A2(new_n416), .A3(KEYINPUT82), .A4(new_n418), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n441), .A2(G101), .A3(new_n442), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n419), .A2(KEYINPUT4), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n443), .A2(new_n444), .B1(new_n214), .B2(new_n216), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT4), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n441), .A2(new_n446), .A3(G101), .A4(new_n442), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n438), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n205), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n436), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n449), .B1(new_n436), .B2(new_n448), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n410), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n436), .A2(new_n448), .A3(new_n449), .ZN(new_n453));
  AND3_X1   g267(.A1(new_n262), .A2(new_n423), .A3(new_n263), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n205), .B1(new_n454), .B2(new_n428), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT12), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI211_X1 g271(.A(KEYINPUT12), .B(new_n205), .C1(new_n454), .C2(new_n428), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n453), .A2(new_n459), .A3(new_n409), .ZN(new_n460));
  AOI21_X1  g274(.A(G902), .B1(new_n452), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n405), .B1(new_n461), .B2(new_n404), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n436), .A2(new_n448), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n205), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(new_n453), .A3(new_n409), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT85), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n453), .A2(new_n459), .A3(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n409), .B(KEYINPUT81), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n466), .B1(new_n453), .B2(new_n459), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n465), .B(G469), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n403), .B1(new_n462), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT20), .ZN(new_n473));
  NOR2_X1   g287(.A1(G475), .A2(G902), .ZN(new_n474));
  INV_X1    g288(.A(G237), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n475), .A2(new_n385), .A3(G214), .ZN(new_n476));
  OR2_X1    g290(.A1(KEYINPUT88), .A2(G143), .ZN(new_n477));
  NAND2_X1  g291(.A1(KEYINPUT88), .A2(G143), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n476), .A2(new_n478), .ZN(new_n480));
  OAI21_X1  g294(.A(G131), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n477), .A2(new_n478), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n482), .A2(G214), .A3(new_n190), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n476), .A2(new_n478), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(new_n203), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT17), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n481), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  OAI211_X1 g301(.A(KEYINPUT17), .B(G131), .C1(new_n479), .C2(new_n480), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n487), .A2(new_n488), .A3(new_n373), .A4(new_n374), .ZN(new_n489));
  XNOR2_X1  g303(.A(G113), .B(G122), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(new_n412), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n356), .A2(new_n358), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT89), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT89), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n365), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(new_n495), .A3(G146), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n366), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT18), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n483), .B(new_n484), .C1(new_n498), .C2(new_n203), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n497), .B(new_n499), .C1(new_n498), .C2(new_n481), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n489), .A2(new_n491), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n481), .A2(new_n485), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n493), .A2(new_n495), .A3(KEYINPUT19), .ZN(new_n503));
  OR2_X1    g317(.A1(new_n492), .A2(KEYINPUT19), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n503), .A2(new_n206), .A3(new_n504), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n502), .A2(new_n505), .A3(new_n362), .A4(new_n364), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n491), .B1(new_n506), .B2(new_n500), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n473), .B(new_n474), .C1(new_n501), .C2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT90), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n506), .A2(new_n500), .ZN(new_n510));
  INV_X1    g324(.A(new_n491), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n489), .A2(new_n491), .A3(new_n500), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT90), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n514), .A2(new_n515), .A3(new_n473), .A4(new_n474), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n474), .B1(new_n501), .B2(new_n507), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT20), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n509), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT15), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G478), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n208), .A2(G128), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n342), .A2(G143), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n523), .A2(new_n524), .A3(new_n196), .ZN(new_n525));
  INV_X1    g339(.A(G122), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G116), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n236), .A2(G122), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(G107), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n527), .A2(new_n528), .A3(new_n415), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n525), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT13), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n523), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n524), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n523), .A2(new_n533), .ZN(new_n536));
  OAI21_X1  g350(.A(G134), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n532), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n236), .A2(KEYINPUT14), .A3(G122), .ZN(new_n539));
  OAI211_X1 g353(.A(G107), .B(new_n539), .C1(new_n529), .C2(KEYINPUT14), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n196), .B1(new_n523), .B2(new_n524), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n540), .B(new_n531), .C1(new_n525), .C2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n401), .A2(new_n338), .A3(G953), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n538), .A2(new_n542), .A3(new_n544), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT92), .B1(new_n548), .B2(new_n327), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n538), .A2(new_n542), .A3(new_n544), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n544), .B1(new_n538), .B2(new_n542), .ZN(new_n551));
  OAI211_X1 g365(.A(KEYINPUT92), .B(new_n327), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n522), .B1(new_n549), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(G902), .B1(new_n546), .B2(new_n547), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n521), .B1(new_n555), .B2(KEYINPUT92), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n491), .B1(new_n489), .B2(new_n500), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n327), .B1(new_n501), .B2(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(KEYINPUT91), .B(G475), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n519), .A2(new_n557), .A3(new_n561), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n385), .A2(G952), .ZN(new_n563));
  NAND2_X1  g377(.A1(G234), .A2(G237), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n564), .A2(G902), .A3(G953), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(KEYINPUT21), .B(G898), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n566), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n562), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(G214), .B1(G237), .B2(G902), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n443), .A2(new_n444), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n574), .B(new_n447), .C1(new_n280), .C2(new_n279), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n237), .A2(new_n239), .A3(KEYINPUT5), .A4(new_n240), .ZN(new_n576));
  NOR3_X1   g390(.A1(new_n236), .A2(KEYINPUT5), .A3(G119), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n577), .A2(new_n242), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n249), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(new_n423), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n575), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(G110), .B(G122), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT86), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n526), .A2(G110), .ZN(new_n587));
  INV_X1    g401(.A(G110), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(G122), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n587), .A2(new_n589), .A3(new_n585), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n583), .A2(new_n591), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n575), .B(new_n582), .C1(new_n590), .C2(new_n586), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(KEYINPUT6), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n357), .B1(new_n214), .B2(new_n216), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n595), .B1(new_n264), .B2(new_n357), .ZN(new_n596));
  INV_X1    g410(.A(G224), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n597), .A2(G953), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n596), .B(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT6), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n583), .A2(new_n600), .A3(new_n591), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n594), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  OR2_X1    g416(.A1(new_n584), .A2(new_n585), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n584), .A2(new_n585), .ZN(new_n604));
  AOI21_X1  g418(.A(KEYINPUT8), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT8), .ZN(new_n606));
  NOR3_X1   g420(.A1(new_n586), .A2(new_n590), .A3(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  AOI22_X1  g422(.A1(new_n579), .A2(new_n249), .B1(new_n419), .B2(new_n422), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n608), .B1(new_n581), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(KEYINPUT7), .B1(new_n597), .B2(G953), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n596), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT87), .ZN(new_n614));
  OR3_X1    g428(.A1(new_n596), .A2(new_n614), .A3(new_n611), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n614), .B1(new_n596), .B2(new_n611), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n613), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(G902), .B1(new_n617), .B2(new_n593), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n602), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(G210), .B1(G237), .B2(G902), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n602), .A2(new_n618), .A3(new_n620), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n573), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n472), .A2(new_n571), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n337), .A2(new_n399), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G101), .ZN(G3));
  NAND3_X1  g441(.A1(new_n303), .A2(new_n306), .A3(new_n307), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n327), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n304), .B1(new_n629), .B2(G472), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n630), .A2(new_n399), .A3(new_n472), .ZN(new_n631));
  INV_X1    g445(.A(new_n570), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n624), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n519), .A2(new_n561), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n548), .A2(KEYINPUT33), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT33), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n546), .A2(new_n636), .A3(new_n547), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n635), .A2(G478), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(G478), .A2(G902), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n548), .A2(new_n327), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n638), .B(new_n639), .C1(G478), .C2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n634), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n633), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n631), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT34), .B(G104), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G6));
  NAND2_X1  g461(.A1(new_n622), .A2(new_n623), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n518), .A2(new_n508), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n554), .A2(new_n556), .ZN(new_n650));
  AND3_X1   g464(.A1(new_n649), .A2(new_n650), .A3(new_n561), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n648), .A2(new_n572), .A3(new_n651), .A4(new_n632), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n631), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT35), .B(G107), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G9));
  NOR2_X1   g470(.A1(new_n368), .A2(new_n375), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n388), .A2(KEYINPUT36), .ZN(new_n658));
  XOR2_X1   g472(.A(new_n657), .B(new_n658), .Z(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n396), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n395), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n571), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n648), .A2(new_n572), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n664), .A2(new_n472), .A3(new_n630), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT93), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT37), .B(G110), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G12));
  INV_X1    g482(.A(new_n403), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n409), .B1(new_n464), .B2(new_n453), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n453), .A2(new_n459), .A3(new_n409), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n404), .B(new_n327), .C1(new_n670), .C2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n405), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n471), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n661), .A2(new_n669), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT94), .B(G900), .Z(new_n676));
  AOI21_X1  g490(.A(new_n566), .B1(new_n568), .B2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n649), .A2(new_n650), .A3(new_n561), .A4(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(KEYINPUT95), .ZN(new_n680));
  AOI22_X1  g494(.A1(new_n518), .A2(new_n508), .B1(new_n559), .B2(new_n560), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT95), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n681), .A2(new_n682), .A3(new_n650), .A4(new_n678), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n675), .A2(new_n684), .A3(new_n663), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n337), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G128), .ZN(G30));
  XOR2_X1   g501(.A(new_n677), .B(KEYINPUT39), .Z(new_n688));
  NAND2_X1  g502(.A1(new_n472), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT97), .ZN(new_n690));
  OR2_X1    g504(.A1(new_n690), .A2(KEYINPUT40), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(KEYINPUT40), .ZN(new_n692));
  INV_X1    g506(.A(G472), .ZN(new_n693));
  AOI21_X1  g507(.A(G902), .B1(new_n332), .B2(new_n291), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n194), .B1(new_n288), .B2(new_n314), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n696), .B1(new_n304), .B2(KEYINPUT32), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n305), .A2(new_n697), .A3(new_n321), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n648), .B(new_n699), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n557), .B1(new_n519), .B2(new_n561), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NOR4_X1   g516(.A1(new_n700), .A2(new_n573), .A3(new_n661), .A4(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n691), .A2(new_n692), .A3(new_n698), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G143), .ZN(G45));
  NAND3_X1  g519(.A1(new_n634), .A2(new_n642), .A3(new_n678), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n675), .A2(new_n663), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n337), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G146), .ZN(G48));
  NOR2_X1   g523(.A1(new_n461), .A2(new_n404), .ZN(new_n710));
  AOI211_X1 g524(.A(G469), .B(G902), .C1(new_n452), .C2(new_n460), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g526(.A(KEYINPUT98), .B1(new_n712), .B2(new_n669), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n327), .B1(new_n670), .B2(new_n671), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(G469), .ZN(new_n715));
  AND4_X1   g529(.A1(KEYINPUT98), .A2(new_n715), .A3(new_n669), .A4(new_n672), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n337), .A2(new_n717), .A3(new_n399), .A4(new_n644), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT41), .B(G113), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G15));
  NOR3_X1   g534(.A1(new_n713), .A2(new_n652), .A3(new_n716), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n337), .A3(new_n399), .ZN(new_n722));
  XOR2_X1   g536(.A(KEYINPUT99), .B(G116), .Z(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G18));
  NAND2_X1  g538(.A1(new_n715), .A2(new_n672), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n403), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n624), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n727), .A2(new_n662), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n337), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G119), .ZN(G21));
  XOR2_X1   g544(.A(KEYINPUT100), .B(G472), .Z(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n732), .B1(new_n628), .B2(new_n327), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n284), .A2(new_n257), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n734), .B1(new_n333), .B2(new_n291), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n189), .B1(new_n735), .B2(new_n306), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n733), .A2(new_n398), .A3(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n663), .A2(new_n702), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n717), .A2(new_n737), .A3(new_n632), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(KEYINPUT101), .B(G122), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(G24));
  NAND2_X1  g555(.A1(new_n735), .A2(new_n306), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n188), .ZN(new_n743));
  AOI21_X1  g557(.A(G902), .B1(new_n290), .B2(new_n303), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n743), .B(new_n661), .C1(new_n744), .C2(new_n732), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  AOI211_X1 g560(.A(new_n677), .B(new_n641), .C1(new_n519), .C2(new_n561), .ZN(new_n747));
  AND4_X1   g561(.A1(new_n669), .A2(new_n747), .A3(new_n624), .A4(new_n712), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(KEYINPUT102), .B(G125), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G27));
  NAND2_X1  g565(.A1(new_n674), .A2(new_n669), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n622), .A2(new_n572), .A3(new_n623), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n337), .A2(new_n399), .A3(new_n747), .A4(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT42), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n336), .A2(new_n322), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n319), .A2(new_n320), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n398), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n752), .A2(new_n706), .A3(new_n753), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(KEYINPUT42), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n757), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G131), .ZN(G33));
  INV_X1    g578(.A(new_n684), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n337), .A2(new_n399), .A3(new_n765), .A4(new_n754), .ZN(new_n766));
  XOR2_X1   g580(.A(KEYINPUT103), .B(G134), .Z(new_n767));
  XNOR2_X1  g581(.A(new_n766), .B(new_n767), .ZN(G36));
  OAI21_X1  g582(.A(new_n465), .B1(new_n469), .B2(new_n470), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n404), .B1(new_n769), .B2(new_n770), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n405), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT104), .ZN(new_n775));
  OR3_X1    g589(.A1(new_n774), .A2(new_n775), .A3(KEYINPUT46), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n775), .B1(new_n774), .B2(KEYINPUT46), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n711), .B1(new_n774), .B2(KEYINPUT46), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n779), .A2(new_n669), .A3(new_n688), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n395), .A2(new_n660), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n630), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(KEYINPUT105), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n634), .A2(new_n641), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(KEYINPUT43), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT44), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n753), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n783), .A2(KEYINPUT44), .A3(new_n785), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n780), .A2(new_n788), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G137), .ZN(G39));
  NOR4_X1   g606(.A1(new_n337), .A2(new_n399), .A3(new_n706), .A4(new_n753), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n779), .A2(KEYINPUT47), .A3(new_n669), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT47), .B1(new_n779), .B2(new_n669), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n793), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G140), .ZN(G42));
  NAND3_X1  g611(.A1(new_n700), .A2(new_n573), .A3(new_n726), .ZN(new_n798));
  XOR2_X1   g612(.A(new_n798), .B(KEYINPUT113), .Z(new_n799));
  NAND3_X1  g613(.A1(new_n785), .A2(new_n737), .A3(new_n566), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT50), .ZN(new_n802));
  AOI211_X1 g616(.A(new_n795), .B(new_n794), .C1(new_n403), .C2(new_n712), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n800), .A2(new_n753), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n802), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  AND4_X1   g620(.A1(new_n566), .A2(new_n785), .A3(new_n726), .A4(new_n789), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n746), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n808), .B(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n698), .ZN(new_n811));
  AND4_X1   g625(.A1(new_n399), .A2(new_n726), .A3(new_n566), .A4(new_n789), .ZN(new_n812));
  INV_X1    g626(.A(new_n634), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n811), .A2(new_n812), .A3(new_n813), .A4(new_n641), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT115), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n810), .A2(KEYINPUT115), .A3(new_n814), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n817), .A2(KEYINPUT51), .A3(new_n818), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n806), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT51), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n821), .B1(new_n806), .B2(new_n815), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n807), .A2(new_n760), .ZN(new_n823));
  XOR2_X1   g637(.A(new_n823), .B(KEYINPUT48), .Z(new_n824));
  NAND2_X1  g638(.A1(new_n811), .A2(new_n812), .ZN(new_n825));
  OAI221_X1 g639(.A(new_n563), .B1(new_n800), .B2(new_n727), .C1(new_n825), .C2(new_n643), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n820), .A2(new_n822), .A3(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n701), .A2(new_n395), .A3(new_n660), .A4(new_n678), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n829), .A2(new_n663), .A3(new_n752), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n698), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n686), .A2(new_n708), .A3(new_n831), .A4(new_n749), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT52), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI22_X1  g648(.A1(new_n337), .A2(new_n685), .B1(new_n746), .B2(new_n748), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n835), .A2(KEYINPUT52), .A3(new_n708), .A4(new_n831), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n834), .B1(KEYINPUT110), .B2(new_n836), .ZN(new_n837));
  XOR2_X1   g651(.A(KEYINPUT110), .B(KEYINPUT111), .Z(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n834), .B(new_n838), .C1(KEYINPUT110), .C2(new_n836), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n562), .B1(new_n813), .B2(new_n642), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n633), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n843), .A2(new_n399), .A3(new_n472), .A4(new_n630), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n626), .A2(new_n665), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n681), .A2(new_n557), .A3(new_n678), .ZN(new_n846));
  OR3_X1    g660(.A1(new_n753), .A2(KEYINPUT108), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n675), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT108), .B1(new_n753), .B2(new_n846), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n746), .A2(KEYINPUT109), .A3(new_n761), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT109), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n789), .A2(new_n472), .A3(new_n747), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n852), .B1(new_n853), .B2(new_n745), .ZN(new_n854));
  AOI22_X1  g668(.A1(new_n337), .A2(new_n850), .B1(new_n851), .B2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n845), .A2(new_n855), .A3(KEYINPUT112), .A4(new_n766), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT112), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n851), .A2(new_n854), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n337), .A2(new_n848), .A3(new_n847), .A4(new_n849), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n858), .A2(new_n766), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n626), .A2(new_n665), .A3(new_n844), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n857), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n856), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n624), .A2(new_n632), .A3(new_n701), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n713), .A2(new_n864), .A3(new_n716), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n737), .A2(new_n865), .B1(new_n728), .B2(new_n337), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n866), .A2(KEYINPUT53), .A3(new_n718), .A4(new_n722), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n867), .B1(new_n757), .B2(new_n762), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n840), .A2(new_n841), .A3(new_n863), .A4(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT54), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n860), .A2(new_n861), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n718), .A2(new_n722), .A3(new_n729), .A4(new_n739), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT107), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n866), .A2(KEYINPUT107), .A3(new_n718), .A4(new_n722), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n872), .A2(new_n875), .A3(new_n763), .A4(new_n876), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n834), .A2(new_n836), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n871), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n869), .A2(new_n870), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(KEYINPUT53), .B1(new_n877), .B2(new_n878), .ZN(new_n881));
  OR2_X1    g695(.A1(new_n877), .A2(KEYINPUT53), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n840), .A2(new_n841), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n880), .B1(new_n884), .B2(new_n870), .ZN(new_n885));
  OAI22_X1  g699(.A1(new_n828), .A2(new_n885), .B1(G952), .B2(G953), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n399), .A2(new_n669), .A3(new_n572), .A4(new_n784), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n887), .B1(KEYINPUT49), .B2(new_n725), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT106), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n700), .B1(KEYINPUT49), .B2(new_n725), .ZN(new_n890));
  OR2_X1    g704(.A1(new_n890), .A2(new_n698), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n886), .B1(new_n889), .B2(new_n891), .ZN(G75));
  NOR2_X1   g706(.A1(new_n385), .A2(G952), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n327), .B1(new_n869), .B2(new_n879), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT56), .B1(new_n895), .B2(G210), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n594), .A2(new_n601), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(new_n599), .Z(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT55), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n894), .B1(new_n896), .B2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT116), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n869), .A2(new_n879), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n902), .B1(new_n903), .B2(G902), .ZN(new_n904));
  AOI211_X1 g718(.A(KEYINPUT116), .B(new_n327), .C1(new_n869), .C2(new_n879), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n621), .ZN(new_n907));
  XNOR2_X1  g721(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n899), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n901), .B1(new_n907), .B2(new_n909), .ZN(G51));
  NAND2_X1  g724(.A1(new_n903), .A2(KEYINPUT54), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT118), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n911), .A2(new_n912), .A3(new_n880), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n903), .A2(KEYINPUT118), .A3(KEYINPUT54), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n405), .B(KEYINPUT57), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n916), .B1(new_n670), .B2(new_n671), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n906), .A2(new_n773), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n893), .B1(new_n917), .B2(new_n918), .ZN(G54));
  NAND2_X1  g733(.A1(KEYINPUT58), .A2(G475), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n904), .A2(new_n905), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n894), .B1(new_n921), .B2(new_n514), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n903), .A2(G902), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(KEYINPUT116), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n895), .A2(new_n902), .ZN(new_n925));
  INV_X1    g739(.A(new_n920), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n514), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(KEYINPUT119), .B1(new_n922), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n893), .B1(new_n927), .B2(new_n928), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT119), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n921), .A2(new_n514), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n930), .A2(new_n934), .ZN(G60));
  AND2_X1   g749(.A1(new_n635), .A2(new_n637), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n639), .B(KEYINPUT59), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n913), .A2(new_n937), .A3(new_n914), .A4(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT120), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n939), .A2(new_n940), .A3(new_n894), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n940), .B1(new_n939), .B2(new_n894), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n937), .B1(new_n885), .B2(new_n938), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(G63));
  NAND2_X1  g758(.A1(G217), .A2(G902), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT60), .Z(new_n946));
  NAND3_X1  g760(.A1(new_n903), .A2(new_n659), .A3(new_n946), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n903), .A2(new_n946), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n894), .B(new_n947), .C1(new_n948), .C2(new_n391), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g764(.A(G953), .B1(new_n569), .B2(new_n597), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n875), .A2(new_n876), .A3(new_n845), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT121), .Z(new_n954));
  AOI21_X1  g768(.A(new_n952), .B1(new_n954), .B2(new_n385), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n897), .B1(G898), .B2(new_n385), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n955), .B(new_n956), .Z(G69));
  NAND2_X1  g771(.A1(G227), .A2(G900), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(G953), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n959), .A2(KEYINPUT124), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT125), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n690), .A2(new_n753), .A3(new_n842), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n962), .A2(new_n337), .A3(new_n399), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n791), .A2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT123), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n964), .B(new_n965), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n835), .A2(new_n708), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n704), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(KEYINPUT62), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n796), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT62), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n704), .A2(new_n971), .A3(new_n967), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT122), .ZN(new_n973));
  OR2_X1    g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n972), .A2(new_n973), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n970), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(G953), .B1(new_n966), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n278), .A2(new_n270), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n503), .A2(new_n504), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n978), .B(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n780), .A2(new_n738), .A3(new_n760), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n763), .A2(new_n766), .A3(new_n967), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n791), .A2(new_n796), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n983), .A2(G953), .ZN(new_n984));
  NAND2_X1  g798(.A1(G900), .A2(G953), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n980), .A2(new_n985), .ZN(new_n986));
  OAI22_X1  g800(.A1(new_n977), .A2(new_n980), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n959), .A2(KEYINPUT124), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n961), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(KEYINPUT123), .B1(new_n791), .B2(new_n963), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n964), .A2(new_n965), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n976), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n980), .B1(new_n992), .B2(new_n385), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n984), .A2(new_n986), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n988), .B(new_n961), .C1(new_n993), .C2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n989), .A2(new_n996), .ZN(G72));
  XOR2_X1   g811(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n998));
  NOR2_X1   g812(.A1(new_n693), .A2(new_n327), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n1000), .B1(new_n992), .B2(new_n954), .ZN(new_n1001));
  INV_X1    g815(.A(new_n695), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n325), .A2(new_n695), .A3(new_n1000), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n884), .A2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT127), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1000), .B1(new_n954), .B2(new_n983), .ZN(new_n1007));
  INV_X1    g821(.A(new_n325), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n893), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AND3_X1   g823(.A1(new_n1003), .A2(new_n1006), .A3(new_n1009), .ZN(G57));
endmodule


