//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0 1 0 1 1 1 1 1 1 1 1 1 0 1 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n783, new_n785, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT13), .Z(new_n203));
  XNOR2_X1  g002(.A(G15gat), .B(G22gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT91), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n205), .B1(new_n206), .B2(G1gat), .ZN(new_n207));
  OR2_X1    g006(.A1(new_n204), .A2(KEYINPUT91), .ZN(new_n208));
  INV_X1    g007(.A(G1gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n204), .A2(KEYINPUT91), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n207), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT92), .ZN(new_n213));
  AOI21_X1  g012(.A(G8gat), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  XOR2_X1   g014(.A(G43gat), .B(G50gat), .Z(new_n216));
  INV_X1    g015(.A(KEYINPUT15), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OR3_X1    g017(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n219));
  OAI21_X1  g018(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n221), .A2(KEYINPUT90), .ZN(new_n222));
  NAND2_X1  g021(.A1(G29gat), .A2(G36gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(new_n221), .B2(KEYINPUT90), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n218), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n218), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n216), .A2(new_n217), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n226), .A2(new_n221), .A3(new_n223), .A4(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n207), .B(new_n211), .C1(new_n213), .C2(G8gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n215), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n229), .B1(new_n215), .B2(new_n230), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n203), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT93), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT93), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n236), .B(new_n203), .C1(new_n232), .C2(new_n233), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n229), .B(KEYINPUT17), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n215), .A2(new_n230), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(new_n231), .A3(new_n202), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT18), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n241), .A2(KEYINPUT18), .A3(new_n231), .A4(new_n202), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n238), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G113gat), .B(G141gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(G169gat), .B(G197gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g050(.A(KEYINPUT89), .B(KEYINPUT12), .Z(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n246), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n238), .A2(new_n253), .A3(new_n244), .A4(new_n245), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT84), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT71), .ZN(new_n259));
  INV_X1    g058(.A(G127gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G134gat), .ZN(new_n261));
  INV_X1    g060(.A(G134gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(G127gat), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n259), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT71), .B1(new_n260), .B2(G134gat), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT72), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n265), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT72), .ZN(new_n268));
  XNOR2_X1  g067(.A(G127gat), .B(G134gat), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n267), .B(new_n268), .C1(new_n269), .C2(new_n259), .ZN(new_n270));
  XNOR2_X1  g069(.A(G113gat), .B(G120gat), .ZN(new_n271));
  OR2_X1    g070(.A1(new_n271), .A2(KEYINPUT1), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n266), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n271), .ZN(new_n274));
  XOR2_X1   g073(.A(KEYINPUT73), .B(KEYINPUT1), .Z(new_n275));
  NAND3_X1  g074(.A1(new_n274), .A2(new_n275), .A3(new_n269), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(G183gat), .ZN(new_n278));
  INV_X1    g077(.A(G190gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT65), .ZN(new_n280));
  AOI22_X1  g079(.A1(new_n278), .A2(new_n279), .B1(new_n280), .B2(KEYINPUT24), .ZN(new_n281));
  NAND2_X1  g080(.A1(G183gat), .A2(G190gat), .ZN(new_n282));
  NOR3_X1   g081(.A1(new_n282), .A2(new_n280), .A3(KEYINPUT24), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT24), .ZN(new_n284));
  AOI22_X1  g083(.A1(new_n284), .A2(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n281), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(G169gat), .A2(G176gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT23), .ZN(new_n288));
  OR2_X1    g087(.A1(G169gat), .A2(G176gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AND2_X1   g089(.A1(KEYINPUT66), .A2(G169gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(KEYINPUT66), .A2(G169gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G176gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT23), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n286), .A2(new_n290), .A3(new_n297), .ZN(new_n298));
  XOR2_X1   g097(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n299));
  NAND2_X1  g098(.A1(new_n278), .A2(KEYINPUT68), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT68), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G183gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n279), .A2(KEYINPUT69), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT69), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G190gat), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n300), .A2(new_n302), .A3(new_n303), .A4(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n282), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n307), .B1(KEYINPUT67), .B2(KEYINPUT24), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT67), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n282), .A2(new_n309), .A3(new_n284), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n306), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT25), .ZN(new_n312));
  NOR2_X1   g111(.A1(G169gat), .A2(G176gat), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n312), .B1(new_n313), .B2(KEYINPUT23), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n290), .A2(new_n314), .ZN(new_n315));
  AOI22_X1  g114(.A1(new_n298), .A2(new_n299), .B1(new_n311), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT27), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G183gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n278), .A2(KEYINPUT27), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n303), .A2(new_n305), .A3(new_n318), .A4(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n307), .B1(new_n320), .B2(KEYINPUT28), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT70), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n322), .B1(new_n278), .B2(KEYINPUT27), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n317), .A2(KEYINPUT70), .A3(G183gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n300), .A2(new_n302), .A3(KEYINPUT27), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT28), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT69), .B(G190gat), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n325), .A2(new_n326), .A3(new_n327), .A4(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT26), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n287), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(new_n289), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n332), .B1(KEYINPUT26), .B2(new_n289), .ZN(new_n333));
  AND3_X1   g132(.A1(new_n321), .A2(new_n329), .A3(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n277), .B1(new_n316), .B2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(KEYINPUT66), .B(G169gat), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n290), .B1(new_n336), .B2(new_n295), .ZN(new_n337));
  OAI22_X1  g136(.A1(new_n284), .A2(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n282), .B1(new_n280), .B2(KEYINPUT24), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n284), .A2(KEYINPUT65), .A3(G183gat), .A4(G190gat), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n299), .B1(new_n337), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n311), .A2(new_n315), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n321), .A2(new_n329), .A3(new_n333), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n344), .A2(new_n273), .A3(new_n276), .A4(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n335), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(G227gat), .ZN(new_n348));
  INV_X1    g147(.A(G233gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT74), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT74), .ZN(new_n352));
  INV_X1    g151(.A(new_n350), .ZN(new_n353));
  AOI211_X1 g152(.A(new_n352), .B(new_n353), .C1(new_n335), .C2(new_n346), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT32), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT33), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n356), .B1(new_n351), .B2(new_n354), .ZN(new_n357));
  XNOR2_X1  g156(.A(G15gat), .B(G43gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n358), .B(KEYINPUT75), .ZN(new_n359));
  XNOR2_X1  g158(.A(G71gat), .B(G99gat), .ZN(new_n360));
  XOR2_X1   g159(.A(new_n359), .B(new_n360), .Z(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n355), .A2(new_n357), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT76), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n335), .A2(new_n346), .A3(new_n353), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT77), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n365), .A2(new_n366), .A3(KEYINPUT34), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n367), .B1(KEYINPUT34), .B2(new_n365), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n366), .B1(new_n365), .B2(KEYINPUT34), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n364), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI221_X1 g169(.A(KEYINPUT32), .B1(new_n356), .B2(new_n361), .C1(new_n351), .C2(new_n354), .ZN(new_n371));
  AND3_X1   g170(.A1(new_n363), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n370), .B1(new_n363), .B2(new_n371), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT36), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT36), .ZN(new_n375));
  INV_X1    g174(.A(new_n369), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n376), .B(new_n367), .C1(KEYINPUT34), .C2(new_n365), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n363), .A2(new_n371), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n377), .B1(new_n363), .B2(new_n371), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n375), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n374), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(G78gat), .B(G106gat), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(G228gat), .A2(G233gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(G155gat), .A2(G162gat), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  AND2_X1   g185(.A1(G141gat), .A2(G148gat), .ZN(new_n387));
  NOR2_X1   g186(.A1(G141gat), .A2(G148gat), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n385), .A2(KEYINPUT2), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n386), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT79), .ZN(new_n392));
  INV_X1    g191(.A(G155gat), .ZN(new_n393));
  INV_X1    g192(.A(G162gat), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT79), .B1(G155gat), .B2(G162gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(G141gat), .B(G148gat), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT80), .B1(new_n385), .B2(KEYINPUT2), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n393), .A2(new_n394), .ZN(new_n401));
  AND2_X1   g200(.A1(KEYINPUT80), .A2(KEYINPUT2), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n385), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n391), .A2(new_n397), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT29), .ZN(new_n405));
  XOR2_X1   g204(.A(G211gat), .B(G218gat), .Z(new_n406));
  INV_X1    g205(.A(G204gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(G197gat), .ZN(new_n408));
  INV_X1    g207(.A(G197gat), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(G204gat), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n408), .A2(new_n410), .A3(KEYINPUT22), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT83), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n406), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(G211gat), .B(G218gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(G197gat), .B(G204gat), .ZN(new_n415));
  INV_X1    g214(.A(G211gat), .ZN(new_n416));
  INV_X1    g215(.A(G218gat), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n414), .B(new_n415), .C1(KEYINPUT22), .C2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n413), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n412), .B1(new_n406), .B2(new_n411), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n405), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT3), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n404), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n406), .A2(new_n411), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n419), .A2(new_n425), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n397), .B(new_n385), .C1(KEYINPUT2), .C2(new_n398), .ZN(new_n427));
  INV_X1    g226(.A(new_n399), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n403), .A2(new_n428), .A3(new_n389), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n427), .A2(new_n429), .A3(new_n423), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n426), .B1(new_n430), .B2(new_n405), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n384), .B1(new_n424), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n431), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n427), .A2(new_n429), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT29), .B1(new_n419), .B2(new_n425), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n434), .B1(new_n435), .B2(KEYINPUT3), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n433), .A2(G228gat), .A3(G233gat), .A4(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(G22gat), .ZN(new_n438));
  AND3_X1   g237(.A1(new_n432), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n438), .B1(new_n432), .B2(new_n437), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n383), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n432), .A2(new_n437), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(G22gat), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n432), .A2(new_n437), .A3(new_n438), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(new_n444), .A3(new_n382), .ZN(new_n445));
  XOR2_X1   g244(.A(KEYINPUT31), .B(G50gat), .Z(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n441), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n447), .B1(new_n441), .B2(new_n445), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n273), .A2(new_n404), .A3(new_n276), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT81), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT81), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n273), .A2(new_n404), .A3(new_n453), .A4(new_n276), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT4), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT4), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n451), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n434), .A2(KEYINPUT3), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n277), .A2(new_n430), .A3(new_n459), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(G225gat), .A2(G233gat), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n463), .A2(KEYINPUT5), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n456), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n452), .A2(new_n457), .A3(new_n454), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n273), .A2(new_n404), .A3(KEYINPUT4), .A4(new_n276), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n460), .A2(new_n462), .A3(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT5), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n452), .A2(new_n454), .ZN(new_n470));
  INV_X1    g269(.A(new_n276), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n271), .A2(KEYINPUT1), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n267), .B1(new_n269), .B2(new_n259), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n472), .B1(new_n473), .B2(KEYINPUT72), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n471), .B1(new_n474), .B2(new_n270), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT82), .B1(new_n475), .B2(new_n404), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT82), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n277), .A2(new_n477), .A3(new_n434), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n462), .B1(new_n470), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n465), .B1(new_n469), .B2(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(G1gat), .B(G29gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n482), .B(KEYINPUT0), .ZN(new_n483));
  XNOR2_X1  g282(.A(G57gat), .B(G85gat), .ZN(new_n484));
  XOR2_X1   g283(.A(new_n483), .B(new_n484), .Z(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n481), .A2(KEYINPUT6), .A3(new_n486), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n485), .B(new_n465), .C1(new_n469), .C2(new_n480), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT6), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR3_X1   g289(.A1(new_n475), .A2(KEYINPUT82), .A3(new_n404), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n477), .B1(new_n277), .B2(new_n434), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n463), .B1(new_n493), .B2(new_n455), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT5), .ZN(new_n495));
  AND3_X1   g294(.A1(new_n460), .A2(new_n462), .A3(new_n467), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n452), .A2(new_n457), .A3(new_n454), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n485), .B1(new_n499), .B2(new_n465), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n487), .B1(new_n490), .B2(new_n500), .ZN(new_n501));
  XOR2_X1   g300(.A(G8gat), .B(G36gat), .Z(new_n502));
  XNOR2_X1  g301(.A(new_n502), .B(KEYINPUT78), .ZN(new_n503));
  XOR2_X1   g302(.A(G64gat), .B(G92gat), .Z(new_n504));
  XNOR2_X1  g303(.A(new_n503), .B(new_n504), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n344), .A2(G226gat), .A3(G233gat), .A4(new_n345), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n316), .A2(new_n334), .ZN(new_n507));
  INV_X1    g306(.A(G226gat), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n405), .B1(new_n508), .B2(new_n349), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n506), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n426), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n506), .B(new_n426), .C1(new_n507), .C2(new_n509), .ZN(new_n513));
  AOI211_X1 g312(.A(KEYINPUT30), .B(new_n505), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT30), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n512), .A2(new_n513), .ZN(new_n516));
  INV_X1    g315(.A(new_n505), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n512), .A2(new_n505), .A3(new_n513), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n514), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n450), .B1(new_n501), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n258), .B1(new_n381), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n501), .A2(new_n521), .ZN(new_n524));
  OR2_X1    g323(.A1(new_n448), .A2(new_n449), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n526), .A2(KEYINPUT84), .A3(new_n374), .A4(new_n380), .ZN(new_n527));
  INV_X1    g326(.A(new_n490), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n481), .A2(KEYINPUT86), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT86), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n530), .B(new_n465), .C1(new_n469), .C2(new_n480), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT87), .B1(new_n532), .B2(new_n486), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT87), .ZN(new_n534));
  AOI211_X1 g333(.A(new_n534), .B(new_n485), .C1(new_n529), .C2(new_n531), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n528), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT38), .B1(new_n516), .B2(new_n517), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n516), .B(KEYINPUT37), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n537), .B1(new_n538), .B2(new_n505), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT38), .ZN(new_n540));
  AND2_X1   g339(.A1(new_n538), .A2(new_n505), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n536), .A2(new_n487), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n530), .B1(new_n499), .B2(new_n465), .ZN(new_n544));
  INV_X1    g343(.A(new_n531), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n486), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(new_n534), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n532), .A2(KEYINPUT87), .A3(new_n486), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n462), .B1(new_n456), .B2(new_n461), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT39), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n470), .A2(new_n462), .A3(new_n479), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT39), .ZN(new_n554));
  OAI211_X1 g353(.A(new_n552), .B(new_n485), .C1(new_n554), .C2(new_n550), .ZN(new_n555));
  NOR2_X1   g354(.A1(KEYINPUT85), .A2(KEYINPUT40), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(new_n520), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n555), .A2(new_n556), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n525), .B1(new_n549), .B2(new_n560), .ZN(new_n561));
  AOI22_X1  g360(.A1(new_n523), .A2(new_n527), .B1(new_n543), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n536), .A2(new_n487), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n520), .A2(KEYINPUT35), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n450), .B(new_n564), .C1(new_n378), .C2(new_n379), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n372), .A2(new_n373), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n567), .A2(new_n501), .A3(new_n521), .A4(new_n450), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n563), .A2(new_n566), .B1(KEYINPUT35), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n257), .B1(new_n562), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(KEYINPUT94), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT94), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n572), .B(new_n257), .C1(new_n562), .C2(new_n569), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(G183gat), .B(G211gat), .Z(new_n575));
  XNOR2_X1  g374(.A(G127gat), .B(G155gat), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n576), .B(KEYINPUT20), .Z(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  AND2_X1   g377(.A1(G71gat), .A2(G78gat), .ZN(new_n579));
  NOR2_X1   g378(.A1(G71gat), .A2(G78gat), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n579), .B1(KEYINPUT9), .B2(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(G57gat), .B(G64gat), .Z(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT95), .ZN(new_n583));
  XNOR2_X1  g382(.A(G57gat), .B(G64gat), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT95), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n581), .B1(new_n583), .B2(new_n586), .ZN(new_n587));
  AOI211_X1 g386(.A(new_n579), .B(new_n580), .C1(new_n582), .C2(KEYINPUT9), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(KEYINPUT96), .B1(new_n589), .B2(KEYINPUT21), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT96), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT21), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n591), .B(new_n592), .C1(new_n587), .C2(new_n588), .ZN(new_n593));
  NAND2_X1  g392(.A1(G231gat), .A2(G233gat), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n594), .B(KEYINPUT97), .Z(new_n595));
  NAND3_X1  g394(.A1(new_n590), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n595), .B1(new_n590), .B2(new_n593), .ZN(new_n598));
  XOR2_X1   g397(.A(KEYINPUT98), .B(KEYINPUT19), .Z(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NOR3_X1   g399(.A1(new_n597), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n590), .A2(new_n593), .ZN(new_n602));
  INV_X1    g401(.A(new_n595), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n599), .B1(new_n604), .B2(new_n596), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n578), .B1(new_n601), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n600), .B1(new_n597), .B2(new_n598), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n604), .A2(new_n596), .A3(new_n599), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n607), .A2(new_n608), .A3(new_n577), .ZN(new_n609));
  INV_X1    g408(.A(new_n589), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n240), .B1(new_n592), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n606), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n611), .B1(new_n606), .B2(new_n609), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n575), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n614), .ZN(new_n616));
  INV_X1    g415(.A(new_n575), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n616), .A2(new_n612), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT99), .ZN(new_n619));
  XOR2_X1   g418(.A(KEYINPUT102), .B(G92gat), .Z(new_n620));
  INV_X1    g419(.A(G85gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(G99gat), .A2(G106gat), .ZN(new_n622));
  AOI22_X1  g421(.A1(new_n620), .A2(new_n621), .B1(KEYINPUT8), .B2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(KEYINPUT101), .B(KEYINPUT7), .ZN(new_n624));
  NAND3_X1  g423(.A1(KEYINPUT100), .A2(G85gat), .A3(G92gat), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n623), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G99gat), .B(G106gat), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n623), .A2(new_n629), .A3(new_n626), .A4(new_n627), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n239), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n633), .ZN(new_n635));
  AND2_X1   g434(.A1(G232gat), .A2(G233gat), .ZN(new_n636));
  AOI22_X1  g435(.A1(new_n635), .A2(new_n229), .B1(KEYINPUT41), .B2(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(G190gat), .B(G218gat), .Z(new_n638));
  AND3_X1   g437(.A1(new_n634), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n638), .B1(new_n634), .B2(new_n637), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n619), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n636), .A2(KEYINPUT41), .ZN(new_n642));
  XNOR2_X1  g441(.A(G134gat), .B(G162gat), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n642), .B(new_n643), .Z(new_n644));
  NAND2_X1  g443(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n644), .ZN(new_n646));
  OAI211_X1 g445(.A(new_n619), .B(new_n646), .C1(new_n639), .C2(new_n640), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n615), .A2(new_n618), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(KEYINPUT103), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n615), .A2(new_n618), .A3(new_n648), .A4(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n633), .A2(new_n610), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT10), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n631), .A2(new_n589), .A3(new_n632), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n635), .A2(KEYINPUT10), .A3(new_n589), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(G230gat), .A2(G233gat), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n654), .A2(new_n656), .ZN(new_n662));
  INV_X1    g461(.A(new_n660), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(G120gat), .B(G148gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(G176gat), .B(G204gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  AND3_X1   g467(.A1(new_n661), .A2(new_n664), .A3(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT105), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n670), .B1(new_n659), .B2(new_n660), .ZN(new_n671));
  AOI211_X1 g470(.A(KEYINPUT105), .B(new_n663), .C1(new_n657), .C2(new_n658), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n664), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n667), .B(KEYINPUT104), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n669), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n653), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n574), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n501), .ZN(new_n679));
  OR2_X1    g478(.A1(new_n679), .A2(KEYINPUT106), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(KEYINPUT106), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n678), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g483(.A(KEYINPUT107), .B(G1gat), .Z(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1324gat));
  AND2_X1   g485(.A1(new_n574), .A2(new_n677), .ZN(new_n687));
  XOR2_X1   g486(.A(KEYINPUT16), .B(G8gat), .Z(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT108), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n687), .A2(new_n520), .A3(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n690), .A2(KEYINPUT42), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT42), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n687), .A2(new_n520), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n692), .B1(new_n693), .B2(G8gat), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n691), .B1(new_n690), .B2(new_n694), .ZN(G1325gat));
  NOR2_X1   g494(.A1(new_n378), .A2(new_n379), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g496(.A(G15gat), .B1(new_n687), .B2(new_n697), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n698), .A2(KEYINPUT109), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n698), .A2(KEYINPUT109), .ZN(new_n700));
  AND3_X1   g499(.A1(new_n687), .A2(G15gat), .A3(new_n381), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(G1326gat));
  OR3_X1    g501(.A1(new_n678), .A2(KEYINPUT110), .A3(new_n450), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT110), .B1(new_n678), .B2(new_n450), .ZN(new_n704));
  XOR2_X1   g503(.A(KEYINPUT43), .B(G22gat), .Z(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT111), .ZN(new_n706));
  AND3_X1   g505(.A1(new_n703), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n706), .B1(new_n703), .B2(new_n704), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(G1327gat));
  NAND2_X1  g508(.A1(new_n615), .A2(new_n618), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(new_n676), .ZN(new_n712));
  INV_X1    g511(.A(new_n648), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n523), .A2(new_n527), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n543), .A2(new_n561), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n563), .A2(new_n566), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n568), .A2(KEYINPUT35), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n572), .B1(new_n722), .B2(new_n257), .ZN(new_n723));
  INV_X1    g522(.A(new_n573), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n715), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OR3_X1    g524(.A1(new_n725), .A2(G29gat), .A3(new_n683), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT45), .ZN(new_n727));
  OR2_X1    g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n526), .A2(new_n374), .A3(new_n380), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n729), .B1(new_n543), .B2(new_n561), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n713), .B1(new_n730), .B2(new_n569), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n648), .A2(new_n732), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n734), .B1(new_n562), .B2(new_n569), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n712), .A2(new_n257), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(G29gat), .B1(new_n739), .B2(new_n683), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n726), .A2(new_n727), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n728), .A2(new_n740), .A3(new_n741), .ZN(G1328gat));
  NOR3_X1   g541(.A1(new_n725), .A2(G36gat), .A3(new_n521), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT46), .ZN(new_n744));
  OAI21_X1  g543(.A(G36gat), .B1(new_n739), .B2(new_n521), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(G1329gat));
  AOI21_X1  g545(.A(new_n714), .B1(new_n571), .B2(new_n573), .ZN(new_n747));
  AOI21_X1  g546(.A(G43gat), .B1(new_n747), .B2(new_n697), .ZN(new_n748));
  INV_X1    g547(.A(new_n739), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n381), .A2(G43gat), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n748), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  XOR2_X1   g550(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n752));
  XNOR2_X1  g551(.A(new_n751), .B(new_n752), .ZN(G1330gat));
  INV_X1    g552(.A(KEYINPUT113), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n450), .B1(new_n725), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n747), .A2(KEYINPUT113), .ZN(new_n756));
  AOI21_X1  g555(.A(G50gat), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(G50gat), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n739), .A2(new_n758), .A3(new_n450), .ZN(new_n759));
  OAI21_X1  g558(.A(KEYINPUT48), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n756), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n525), .B1(new_n747), .B2(KEYINPUT113), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n758), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT48), .ZN(new_n764));
  INV_X1    g563(.A(new_n759), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n760), .A2(new_n766), .ZN(G1331gat));
  AND2_X1   g566(.A1(new_n543), .A2(new_n561), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n721), .B1(new_n768), .B2(new_n729), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n653), .A2(new_n257), .A3(new_n675), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n682), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g573(.A(new_n521), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT114), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n778));
  XOR2_X1   g577(.A(new_n777), .B(new_n778), .Z(G1333gat));
  NAND2_X1  g578(.A1(new_n772), .A2(new_n381), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(G71gat), .ZN(new_n781));
  OR3_X1    g580(.A1(new_n771), .A2(G71gat), .A3(new_n696), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XOR2_X1   g582(.A(new_n783), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g583(.A1(new_n772), .A2(new_n525), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g585(.A1(new_n711), .A2(new_n257), .A3(new_n675), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n736), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(KEYINPUT115), .B1(new_n788), .B2(new_n683), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(G85gat), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n788), .A2(KEYINPUT115), .A3(new_n683), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n711), .A2(new_n257), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n769), .A2(KEYINPUT51), .A3(new_n713), .A4(new_n792), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n713), .B(new_n792), .C1(new_n730), .C2(new_n569), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT51), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n682), .A2(new_n621), .A3(new_n676), .ZN(new_n799));
  OAI22_X1  g598(.A1(new_n790), .A2(new_n791), .B1(new_n798), .B2(new_n799), .ZN(G1336gat));
  NAND4_X1  g599(.A1(new_n733), .A2(new_n520), .A3(new_n735), .A4(new_n787), .ZN(new_n801));
  INV_X1    g600(.A(new_n620), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n675), .A2(new_n521), .A3(G92gat), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n794), .A2(new_n795), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n794), .A2(new_n795), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT117), .ZN(new_n808));
  XNOR2_X1  g607(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n803), .A2(new_n807), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n811));
  AOI22_X1  g610(.A1(new_n802), .A2(new_n801), .B1(new_n797), .B2(new_n804), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n808), .B1(new_n812), .B2(new_n809), .ZN(new_n814));
  OAI21_X1  g613(.A(KEYINPUT118), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n803), .A2(new_n807), .A3(new_n809), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(KEYINPUT117), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n803), .A2(new_n807), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT52), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n817), .A2(new_n819), .A3(new_n820), .A4(new_n810), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n815), .A2(new_n821), .ZN(G1337gat));
  NAND3_X1  g621(.A1(new_n736), .A2(new_n381), .A3(new_n787), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(G99gat), .ZN(new_n824));
  OR3_X1    g623(.A1(new_n696), .A2(G99gat), .A3(new_n675), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n824), .B1(new_n798), .B2(new_n825), .ZN(G1338gat));
  OAI21_X1  g625(.A(G106gat), .B1(new_n788), .B2(new_n450), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT119), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n675), .A2(G106gat), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n797), .A2(new_n525), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n829), .A2(new_n832), .A3(KEYINPUT53), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n827), .B(new_n831), .C1(new_n828), .C2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(G1339gat));
  INV_X1    g635(.A(new_n257), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n650), .A2(new_n837), .A3(new_n652), .A4(new_n675), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n661), .A2(KEYINPUT105), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n659), .A2(new_n670), .A3(new_n660), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n840), .B1(new_n659), .B2(new_n660), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n657), .A2(new_n663), .A3(new_n658), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n668), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n842), .A2(KEYINPUT55), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(KEYINPUT120), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT120), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n842), .A2(new_n845), .A3(new_n848), .A4(KEYINPUT55), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n669), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n842), .A2(new_n845), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT121), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT55), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n851), .A2(new_n853), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(KEYINPUT121), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n202), .B1(new_n241), .B2(new_n231), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n232), .A2(new_n233), .A3(new_n203), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n251), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AND4_X1   g658(.A1(new_n256), .A2(new_n645), .A3(new_n647), .A4(new_n859), .ZN(new_n860));
  AND4_X1   g659(.A1(new_n850), .A2(new_n854), .A3(new_n856), .A4(new_n860), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n256), .A2(new_n859), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n676), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n856), .A2(new_n257), .A3(new_n854), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n847), .A2(new_n849), .ZN(new_n865));
  INV_X1    g664(.A(new_n669), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n863), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n861), .B1(new_n868), .B2(new_n648), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n838), .B1(new_n869), .B2(new_n711), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n682), .A2(new_n521), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n567), .A2(new_n450), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(G113gat), .B1(new_n875), .B2(new_n257), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n873), .A2(new_n525), .A3(new_n696), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n257), .A2(G113gat), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(G1340gat));
  AOI21_X1  g678(.A(G120gat), .B1(new_n875), .B2(new_n676), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n676), .A2(G120gat), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n880), .B1(new_n877), .B2(new_n881), .ZN(G1341gat));
  NAND3_X1  g681(.A1(new_n875), .A2(new_n260), .A3(new_n711), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n877), .A2(new_n711), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n883), .B1(new_n884), .B2(new_n260), .ZN(G1342gat));
  NOR4_X1   g684(.A1(new_n873), .A2(G134gat), .A3(new_n874), .A4(new_n648), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT56), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n877), .A2(new_n713), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n887), .B1(new_n262), .B2(new_n888), .ZN(G1343gat));
  NOR2_X1   g688(.A1(new_n381), .A2(new_n450), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n837), .A2(G141gat), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n873), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n838), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n850), .A2(new_n854), .A3(new_n856), .A4(new_n860), .ZN(new_n895));
  INV_X1    g694(.A(new_n863), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n671), .A2(new_n672), .A3(KEYINPUT54), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n661), .A2(KEYINPUT54), .A3(new_n844), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n667), .ZN(new_n899));
  OAI21_X1  g698(.A(KEYINPUT122), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT122), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n842), .A2(new_n901), .A3(new_n845), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n900), .A2(new_n853), .A3(new_n902), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n903), .A2(new_n257), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n896), .B1(new_n904), .B2(new_n850), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n895), .B1(new_n905), .B2(new_n713), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n894), .B1(new_n906), .B2(new_n710), .ZN(new_n907));
  OAI21_X1  g706(.A(KEYINPUT57), .B1(new_n907), .B2(new_n450), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT57), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n870), .A2(new_n909), .A3(new_n525), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n871), .A2(new_n381), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n908), .A2(new_n910), .A3(new_n257), .A4(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n893), .B1(new_n912), .B2(G141gat), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT58), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT123), .ZN(new_n916));
  AND3_X1   g715(.A1(new_n913), .A2(new_n916), .A3(new_n914), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n913), .B2(new_n914), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(G1344gat));
  NOR3_X1   g718(.A1(new_n675), .A2(G148gat), .A3(new_n520), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n870), .A2(new_n682), .A3(new_n890), .A4(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT59), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n865), .A2(new_n903), .A3(new_n257), .A4(new_n866), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n713), .B1(new_n923), .B2(new_n863), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n710), .B1(new_n924), .B2(new_n861), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(new_n838), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n450), .B1(new_n926), .B2(KEYINPUT124), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT124), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n907), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(KEYINPUT57), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n868), .A2(new_n648), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(new_n895), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n894), .B1(new_n932), .B2(new_n710), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n933), .A2(new_n909), .A3(new_n450), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n676), .B(new_n911), .C1(new_n930), .C2(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n922), .B1(new_n935), .B2(G148gat), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n908), .A2(new_n910), .A3(new_n911), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n937), .A2(new_n675), .ZN(new_n938));
  INV_X1    g737(.A(G148gat), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n938), .A2(KEYINPUT59), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n921), .B1(new_n936), .B2(new_n940), .ZN(G1345gat));
  OAI21_X1  g740(.A(G155gat), .B1(new_n937), .B2(new_n710), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n873), .A2(new_n891), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n943), .A2(new_n393), .A3(new_n711), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n942), .A2(new_n944), .ZN(G1346gat));
  OAI21_X1  g744(.A(G162gat), .B1(new_n937), .B2(new_n648), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n943), .A2(new_n394), .A3(new_n713), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(G1347gat));
  INV_X1    g747(.A(KEYINPUT125), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n682), .A2(new_n521), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n696), .A2(new_n525), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n949), .B1(new_n933), .B2(new_n952), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n870), .A2(KEYINPUT125), .A3(new_n951), .A4(new_n950), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g754(.A(G169gat), .B1(new_n955), .B2(new_n837), .ZN(new_n956));
  NOR4_X1   g755(.A1(new_n933), .A2(new_n521), .A3(new_n874), .A4(new_n682), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n957), .A2(new_n257), .A3(new_n293), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n956), .A2(new_n958), .ZN(G1348gat));
  OAI21_X1  g758(.A(G176gat), .B1(new_n955), .B2(new_n675), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n957), .A2(new_n294), .A3(new_n676), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(G1349gat));
  NAND2_X1  g761(.A1(new_n300), .A2(new_n302), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n963), .B1(new_n955), .B2(new_n710), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n957), .A2(new_n318), .A3(new_n319), .A4(new_n711), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(KEYINPUT60), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT60), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n964), .A2(new_n965), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n967), .A2(new_n969), .ZN(G1350gat));
  INV_X1    g769(.A(KEYINPUT61), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n953), .A2(new_n713), .A3(new_n954), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT126), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n972), .A2(new_n973), .A3(G190gat), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n973), .B1(new_n972), .B2(G190gat), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n971), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n972), .A2(G190gat), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(KEYINPUT126), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n972), .A2(new_n973), .A3(G190gat), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n978), .A2(KEYINPUT61), .A3(new_n979), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n957), .A2(new_n328), .A3(new_n713), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n976), .A2(new_n980), .A3(new_n981), .ZN(G1351gat));
  NOR2_X1   g781(.A1(new_n933), .A2(new_n682), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n891), .A2(new_n521), .ZN(new_n984));
  AND2_X1   g783(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g784(.A(G197gat), .B1(new_n985), .B2(new_n257), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n930), .A2(new_n934), .ZN(new_n987));
  NOR3_X1   g786(.A1(new_n682), .A2(new_n521), .A3(new_n381), .ZN(new_n988));
  INV_X1    g787(.A(new_n988), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g789(.A1(new_n837), .A2(new_n409), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n986), .B1(new_n990), .B2(new_n991), .ZN(G1352gat));
  XNOR2_X1  g791(.A(KEYINPUT127), .B(G204gat), .ZN(new_n993));
  AND4_X1   g792(.A1(new_n676), .A2(new_n983), .A3(new_n984), .A4(new_n993), .ZN(new_n994));
  XNOR2_X1  g793(.A(new_n994), .B(KEYINPUT62), .ZN(new_n995));
  NOR3_X1   g794(.A1(new_n987), .A2(new_n675), .A3(new_n989), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n995), .B1(new_n996), .B2(new_n993), .ZN(G1353gat));
  NAND3_X1  g796(.A1(new_n985), .A2(new_n416), .A3(new_n711), .ZN(new_n998));
  OAI211_X1 g797(.A(new_n711), .B(new_n988), .C1(new_n930), .C2(new_n934), .ZN(new_n999));
  AND3_X1   g798(.A1(new_n999), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1000));
  AOI21_X1  g799(.A(KEYINPUT63), .B1(new_n999), .B2(G211gat), .ZN(new_n1001));
  OAI21_X1  g800(.A(new_n998), .B1(new_n1000), .B2(new_n1001), .ZN(G1354gat));
  NAND3_X1  g801(.A1(new_n985), .A2(new_n417), .A3(new_n713), .ZN(new_n1003));
  NOR3_X1   g802(.A1(new_n987), .A2(new_n648), .A3(new_n989), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n1003), .B1(new_n1004), .B2(new_n417), .ZN(G1355gat));
endmodule


