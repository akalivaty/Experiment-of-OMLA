//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 0 0 1 1 0 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 0 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n554,
    new_n555, new_n556, new_n557, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n566, new_n568, new_n569, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n599, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n636, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1164, new_n1165, new_n1166,
    new_n1167;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT65), .Z(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  AOI22_X1  g035(.A1(new_n460), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AND3_X1   g038(.A1(KEYINPUT66), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(KEYINPUT3), .B1(KEYINPUT66), .B2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n463), .B1(G137), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  XOR2_X1   g046(.A(new_n471), .B(KEYINPUT67), .Z(new_n472));
  AND2_X1   g047(.A1(new_n468), .A2(new_n472), .ZN(G160));
  NOR2_X1   g048(.A1(new_n464), .A2(new_n465), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(new_n462), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n467), .A2(G136), .ZN(new_n477));
  NOR2_X1   g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(new_n462), .B2(G112), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n476), .B(new_n477), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  NOR2_X1   g056(.A1(KEYINPUT4), .A2(G2105), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n460), .A2(G138), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n483), .B(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  OAI21_X1  g061(.A(KEYINPUT4), .B1(new_n466), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n469), .B1(new_n490), .B2(G2105), .ZN(new_n491));
  AOI22_X1  g066(.A1(new_n475), .A2(G126), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n488), .A2(new_n492), .ZN(G164));
  INV_X1    g068(.A(KEYINPUT72), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G543), .ZN(new_n495));
  INV_X1    g070(.A(G543), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT72), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n495), .A2(new_n497), .A3(KEYINPUT5), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT73), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT73), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT5), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n496), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT74), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT74), .B1(new_n507), .B2(new_n496), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n499), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT69), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT69), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n509), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT71), .B1(new_n511), .B2(KEYINPUT6), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n519), .A2(new_n520), .A3(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT70), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n524), .B1(new_n515), .B2(KEYINPUT6), .ZN(new_n525));
  AOI211_X1 g100(.A(KEYINPUT70), .B(new_n520), .C1(new_n512), .C2(new_n514), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n517), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n516), .A2(new_n528), .ZN(G166));
  INV_X1    g104(.A(KEYINPUT76), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT69), .B(G651), .ZN(new_n532));
  OAI21_X1  g107(.A(KEYINPUT70), .B1(new_n532), .B2(new_n520), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n515), .A2(new_n524), .A3(KEYINPUT6), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n535), .A2(KEYINPUT76), .A3(new_n523), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n531), .A2(G543), .A3(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G51), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n540), .A2(new_n541), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT7), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n522), .B1(new_n533), .B2(new_n534), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n509), .A2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  XNOR2_X1  g124(.A(KEYINPUT77), .B(G89), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n539), .A2(new_n544), .A3(new_n546), .A4(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(G168));
  AND2_X1   g128(.A1(new_n538), .A2(G52), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G90), .ZN(new_n556));
  OAI22_X1  g131(.A1(new_n555), .A2(new_n515), .B1(new_n556), .B2(new_n548), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n554), .A2(new_n557), .ZN(G171));
  NAND2_X1  g133(.A1(new_n538), .A2(G43), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n560));
  OR2_X1    g135(.A1(new_n560), .A2(new_n515), .ZN(new_n561));
  INV_X1    g136(.A(G81), .ZN(new_n562));
  OAI211_X1 g137(.A(new_n559), .B(new_n561), .C1(new_n562), .C2(new_n548), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  AND3_X1   g140(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G36), .ZN(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT8), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n566), .A2(new_n569), .ZN(G188));
  AOI21_X1  g145(.A(KEYINPUT76), .B1(new_n535), .B2(new_n523), .ZN(new_n571));
  AOI211_X1 g146(.A(new_n530), .B(new_n522), .C1(new_n533), .C2(new_n534), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n573), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n531), .A2(G53), .A3(G543), .A4(new_n536), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT9), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n504), .A2(new_n505), .ZN(new_n578));
  NOR3_X1   g153(.A1(new_n507), .A2(KEYINPUT74), .A3(new_n496), .ZN(new_n579));
  OAI211_X1 g154(.A(G65), .B(new_n498), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(G78), .A2(G543), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n511), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AND3_X1   g157(.A1(new_n509), .A2(new_n547), .A3(G91), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n574), .A2(new_n577), .A3(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT78), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n574), .A2(new_n577), .A3(KEYINPUT78), .A4(new_n584), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G299));
  INV_X1    g165(.A(G171), .ZN(G301));
  INV_X1    g166(.A(KEYINPUT79), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n552), .A2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n542), .A2(new_n543), .B1(new_n549), .B2(new_n550), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n594), .A2(KEYINPUT79), .A3(new_n546), .A4(new_n539), .ZN(new_n595));
  AND2_X1   g170(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G286));
  INV_X1    g172(.A(G166), .ZN(G303));
  NAND2_X1  g173(.A1(new_n538), .A2(G49), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n509), .A2(G74), .ZN(new_n600));
  AOI22_X1  g175(.A1(G87), .A2(new_n549), .B1(new_n600), .B2(G651), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n599), .A2(new_n601), .ZN(G288));
  NAND2_X1  g177(.A1(new_n509), .A2(G61), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT80), .ZN(new_n604));
  AND2_X1   g179(.A1(G73), .A2(G543), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n532), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AND2_X1   g181(.A1(new_n509), .A2(G86), .ZN(new_n607));
  AND2_X1   g182(.A1(G48), .A2(G543), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n547), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n606), .A2(new_n609), .ZN(G305));
  AOI22_X1  g185(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n611), .A2(new_n515), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n549), .A2(G85), .ZN(new_n613));
  INV_X1    g188(.A(G47), .ZN(new_n614));
  OAI211_X1 g189(.A(new_n612), .B(new_n613), .C1(new_n614), .C2(new_n537), .ZN(G290));
  NAND2_X1  g190(.A1(G301), .A2(G868), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT81), .ZN(new_n617));
  INV_X1    g192(.A(G66), .ZN(new_n618));
  AOI211_X1 g193(.A(new_n618), .B(new_n499), .C1(new_n506), .C2(new_n508), .ZN(new_n619));
  NAND2_X1  g194(.A1(G79), .A2(G543), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n617), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n509), .A2(G66), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n623), .A2(KEYINPUT81), .A3(new_n620), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n622), .A2(new_n624), .A3(G651), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n573), .A2(G54), .A3(G543), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT10), .ZN(new_n627));
  INV_X1    g202(.A(G92), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n548), .B2(new_n628), .ZN(new_n629));
  NAND4_X1  g204(.A1(new_n509), .A2(new_n547), .A3(KEYINPUT10), .A4(G92), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AND3_X1   g206(.A1(new_n625), .A2(new_n626), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT82), .Z(new_n633));
  OAI21_X1  g208(.A(new_n616), .B1(new_n633), .B2(G868), .ZN(G284));
  OAI21_X1  g209(.A(new_n616), .B1(new_n633), .B2(G868), .ZN(G321));
  NAND2_X1  g210(.A1(G286), .A2(G868), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(G868), .B2(new_n589), .ZN(G297));
  XOR2_X1   g212(.A(G297), .B(KEYINPUT83), .Z(G280));
  INV_X1    g213(.A(G559), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n633), .B1(new_n639), .B2(G860), .ZN(G148));
  NAND2_X1  g215(.A1(new_n633), .A2(new_n639), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(G868), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n642), .A2(KEYINPUT84), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(KEYINPUT84), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n643), .B(new_n644), .C1(G868), .C2(new_n564), .ZN(G323));
  XNOR2_X1  g220(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g221(.A1(new_n460), .A2(new_n470), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT12), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT13), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2100), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n475), .A2(G123), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n467), .A2(G135), .ZN(new_n652));
  NOR2_X1   g227(.A1(G99), .A2(G2105), .ZN(new_n653));
  OAI21_X1  g228(.A(G2104), .B1(new_n462), .B2(G111), .ZN(new_n654));
  OAI211_X1 g229(.A(new_n651), .B(new_n652), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2096), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n650), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT85), .Z(G156));
  XNOR2_X1  g233(.A(G2451), .B(G2454), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2443), .B(G2446), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1341), .B(G1348), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n662), .B(new_n663), .Z(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT15), .B(G2430), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2435), .ZN(new_n666));
  XOR2_X1   g241(.A(G2427), .B(G2438), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(KEYINPUT14), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n664), .B(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(G14), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(G401));
  XOR2_X1   g247(.A(G2072), .B(G2078), .Z(new_n673));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G2067), .B(G2678), .Z(new_n676));
  OR2_X1    g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n673), .B1(new_n677), .B2(KEYINPUT18), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(G2100), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n675), .A2(new_n676), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n677), .A2(new_n680), .A3(KEYINPUT17), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT18), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n679), .B(new_n683), .Z(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT86), .B(G2096), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(G227));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  XOR2_X1   g263(.A(G1956), .B(G2474), .Z(new_n689));
  XOR2_X1   g264(.A(G1961), .B(G1966), .Z(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n688), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n689), .A2(new_n690), .ZN(new_n694));
  AOI22_X1  g269(.A1(new_n692), .A2(KEYINPUT20), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n694), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n696), .A2(new_n688), .A3(new_n691), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n695), .B(new_n697), .C1(KEYINPUT20), .C2(new_n692), .ZN(new_n698));
  XOR2_X1   g273(.A(G1991), .B(G1996), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(G229));
  MUX2_X1   g279(.A(G24), .B(G290), .S(G16), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(G1986), .ZN(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G6), .ZN(new_n708));
  INV_X1    g283(.A(G305), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(new_n707), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT89), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT32), .B(G1981), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G288), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n714), .A2(new_n707), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n707), .B2(G23), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT33), .B(G1976), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT90), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n716), .A2(new_n718), .ZN(new_n720));
  NOR2_X1   g295(.A1(G166), .A2(new_n707), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n707), .B2(G22), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  AOI211_X1 g298(.A(new_n719), .B(new_n720), .C1(G1971), .C2(new_n723), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n713), .B(new_n724), .C1(G1971), .C2(new_n723), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n706), .B1(new_n725), .B2(KEYINPUT34), .ZN(new_n726));
  INV_X1    g301(.A(G29), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G25), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n467), .A2(G131), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT87), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G119), .B2(new_n475), .ZN(new_n731));
  OR2_X1    g306(.A1(G95), .A2(G2105), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n732), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n728), .B1(new_n735), .B2(new_n727), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT88), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT35), .B(G1991), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n726), .B(new_n739), .C1(KEYINPUT34), .C2(new_n725), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT36), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n655), .A2(new_n727), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT96), .Z(new_n743));
  NOR2_X1   g318(.A1(G164), .A2(new_n727), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G27), .B2(new_n727), .ZN(new_n745));
  INV_X1    g320(.A(G2078), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n727), .A2(G33), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n467), .A2(G139), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT93), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n470), .A2(G103), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT25), .Z(new_n751));
  AOI22_X1  g326(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n749), .B(new_n751), .C1(new_n462), .C2(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n747), .B1(new_n753), .B2(G29), .ZN(new_n754));
  INV_X1    g329(.A(G2072), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n745), .A2(new_n746), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT27), .B(G1996), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT95), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n467), .A2(G141), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT94), .ZN(new_n760));
  NAND3_X1  g335(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT26), .Z(new_n762));
  AOI22_X1  g337(.A1(new_n475), .A2(G129), .B1(G105), .B2(new_n470), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n760), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(G29), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G29), .B2(G32), .ZN(new_n767));
  OAI221_X1 g342(.A(new_n756), .B1(new_n746), .B2(new_n745), .C1(new_n758), .C2(new_n767), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT31), .B(G11), .Z(new_n769));
  INV_X1    g344(.A(KEYINPUT30), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n727), .B1(new_n770), .B2(G28), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n770), .B2(G28), .ZN(new_n772));
  AND2_X1   g347(.A1(KEYINPUT24), .A2(G34), .ZN(new_n773));
  NOR2_X1   g348(.A1(KEYINPUT24), .A2(G34), .ZN(new_n774));
  NOR3_X1   g349(.A1(new_n773), .A2(new_n774), .A3(G29), .ZN(new_n775));
  INV_X1    g350(.A(G160), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(G29), .ZN(new_n777));
  INV_X1    g352(.A(G2084), .ZN(new_n778));
  AOI211_X1 g353(.A(new_n769), .B(new_n772), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n767), .A2(new_n758), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n754), .A2(new_n755), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n777), .A2(new_n778), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n779), .A2(new_n780), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n768), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n707), .A2(G19), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n564), .B2(new_n707), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(G1341), .Z(new_n787));
  AND2_X1   g362(.A1(new_n727), .A2(G26), .ZN(new_n788));
  OR2_X1    g363(.A1(G104), .A2(G2105), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT92), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n469), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI221_X1 g366(.A(new_n791), .B1(new_n790), .B2(new_n789), .C1(G116), .C2(new_n462), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n475), .A2(G128), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n467), .A2(G140), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n788), .B1(new_n795), .B2(G29), .ZN(new_n796));
  MUX2_X1   g371(.A(new_n788), .B(new_n796), .S(KEYINPUT28), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G2067), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n727), .A2(G35), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G162), .B2(new_n727), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT29), .B(G2090), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n784), .A2(new_n787), .A3(new_n798), .A4(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(G4), .A2(G16), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(new_n633), .B2(G16), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT91), .B(G1348), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n707), .A2(G20), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT97), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT23), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n589), .B2(new_n707), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(G1956), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n707), .A2(G21), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G168), .B2(new_n707), .ZN(new_n814));
  INV_X1    g389(.A(G1966), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n707), .A2(G5), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G171), .B2(new_n707), .ZN(new_n818));
  INV_X1    g393(.A(G1961), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  NOR4_X1   g396(.A1(new_n803), .A2(new_n807), .A3(new_n812), .A4(new_n821), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n741), .A2(new_n743), .A3(new_n822), .ZN(G150));
  INV_X1    g398(.A(G150), .ZN(G311));
  INV_X1    g399(.A(G55), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n537), .A2(new_n825), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n827));
  INV_X1    g402(.A(G93), .ZN(new_n828));
  OAI22_X1  g403(.A1(new_n827), .A2(new_n515), .B1(new_n828), .B2(new_n548), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(G860), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT37), .Z(new_n833));
  NAND2_X1  g408(.A1(new_n633), .A2(G559), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT38), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n563), .B(new_n830), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT39), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n835), .B(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n833), .B1(new_n838), .B2(G860), .ZN(G145));
  XNOR2_X1  g414(.A(G160), .B(G162), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n655), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n475), .A2(G130), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n467), .A2(G142), .ZN(new_n843));
  NOR2_X1   g418(.A1(G106), .A2(G2105), .ZN(new_n844));
  OAI21_X1  g419(.A(G2104), .B1(new_n462), .B2(G118), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n842), .B(new_n843), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n734), .B(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT100), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n648), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n764), .B(new_n795), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT98), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n485), .A2(new_n851), .A3(new_n487), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n851), .B1(new_n485), .B2(new_n487), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n492), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n850), .B(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n753), .B(KEYINPUT99), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT99), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n856), .B1(new_n859), .B2(new_n753), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n849), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(KEYINPUT101), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n849), .A2(new_n862), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n863), .A2(KEYINPUT101), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n841), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(G37), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n862), .B1(new_n849), .B2(KEYINPUT102), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n870), .B1(new_n865), .B2(KEYINPUT102), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n868), .B(new_n869), .C1(new_n841), .C2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT40), .ZN(G395));
  NAND3_X1  g448(.A1(new_n587), .A2(new_n588), .A3(new_n632), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n587), .A2(KEYINPUT103), .A3(new_n588), .A4(new_n632), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n632), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n589), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT104), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n632), .B1(new_n587), .B2(new_n588), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(KEYINPUT104), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n878), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT41), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n878), .A2(KEYINPUT41), .A3(new_n880), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n641), .B(new_n836), .ZN(new_n891));
  MUX2_X1   g466(.A(new_n881), .B(new_n890), .S(new_n891), .Z(new_n892));
  NAND2_X1  g467(.A1(new_n714), .A2(G303), .ZN(new_n893));
  NAND2_X1  g468(.A1(G288), .A2(G166), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n893), .A2(G305), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(G305), .B1(new_n893), .B2(new_n894), .ZN(new_n896));
  XNOR2_X1  g471(.A(G290), .B(KEYINPUT105), .ZN(new_n897));
  OR3_X1    g472(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n897), .B1(new_n895), .B2(new_n896), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n900), .B(KEYINPUT42), .Z(new_n901));
  AND2_X1   g476(.A1(new_n892), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n892), .A2(new_n901), .ZN(new_n903));
  OAI21_X1  g478(.A(G868), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n904), .B1(G868), .B2(new_n830), .ZN(G295));
  OAI21_X1  g480(.A(new_n904), .B1(G868), .B2(new_n830), .ZN(G331));
  NOR2_X1   g481(.A1(G171), .A2(new_n552), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  OAI211_X1 g483(.A(new_n836), .B(new_n908), .C1(new_n596), .C2(G301), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n563), .B(new_n831), .ZN(new_n910));
  AOI21_X1  g485(.A(G301), .B1(new_n593), .B2(new_n595), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n910), .B1(new_n911), .B2(new_n907), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n884), .A2(KEYINPUT104), .ZN(new_n914));
  AOI211_X1 g489(.A(new_n882), .B(new_n632), .C1(new_n587), .C2(new_n588), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(KEYINPUT41), .B1(new_n916), .B2(new_n878), .ZN(new_n917));
  INV_X1    g492(.A(new_n889), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n913), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n909), .A2(new_n912), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n881), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n919), .A2(new_n900), .A3(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(KEYINPUT109), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n898), .A2(KEYINPUT107), .A3(new_n899), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT107), .B1(new_n898), .B2(new_n899), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n920), .A2(new_n881), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(KEYINPUT110), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n881), .A2(KEYINPUT41), .ZN(new_n930));
  AOI211_X1 g505(.A(new_n920), .B(new_n930), .C1(KEYINPUT41), .C2(new_n886), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n927), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n924), .A2(KEYINPUT43), .A3(new_n932), .A4(new_n869), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n920), .B1(new_n888), .B2(new_n889), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT106), .B1(new_n934), .B2(new_n928), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n919), .A2(new_n936), .A3(new_n921), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n935), .A2(new_n927), .A3(new_n937), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n938), .A2(KEYINPUT108), .A3(new_n869), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT108), .B1(new_n938), .B2(new_n869), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n939), .A2(new_n940), .A3(new_n923), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n933), .B1(new_n941), .B2(KEYINPUT43), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT44), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n924), .A2(new_n944), .A3(new_n932), .A4(new_n869), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n945), .B1(new_n941), .B2(new_n944), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n943), .A2(new_n948), .ZN(G397));
  INV_X1    g524(.A(KEYINPUT49), .ZN(new_n950));
  NOR2_X1   g525(.A1(G305), .A2(G1981), .ZN(new_n951));
  INV_X1    g526(.A(G1981), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n952), .B1(new_n606), .B2(new_n609), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n950), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT115), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT115), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n956), .B(new_n950), .C1(new_n951), .C2(new_n953), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  OR3_X1    g533(.A1(new_n951), .A2(new_n950), .A3(new_n953), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n488), .A2(KEYINPUT98), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n852), .ZN(new_n961));
  AOI21_X1  g536(.A(G1384), .B1(new_n961), .B2(new_n492), .ZN(new_n962));
  XOR2_X1   g537(.A(KEYINPUT111), .B(G40), .Z(new_n963));
  NAND2_X1  g538(.A1(G160), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G8), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n958), .A2(new_n959), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G1976), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n969), .B1(new_n971), .B2(G288), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT52), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT52), .B1(G288), .B2(new_n971), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n969), .B(new_n974), .C1(new_n971), .C2(G288), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n970), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT113), .ZN(new_n978));
  INV_X1    g553(.A(G1384), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n855), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n978), .B1(new_n980), .B2(KEYINPUT50), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT50), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n962), .A2(KEYINPUT113), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G2090), .ZN(new_n985));
  NOR2_X1   g560(.A1(G164), .A2(G1384), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n986), .A2(new_n982), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n984), .A2(new_n985), .A3(new_n965), .A4(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n962), .A2(KEYINPUT45), .ZN(new_n990));
  OR2_X1    g565(.A1(G164), .A2(G1384), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n990), .A2(new_n993), .A3(new_n965), .ZN(new_n994));
  XNOR2_X1  g569(.A(KEYINPUT112), .B(G1971), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n968), .B1(new_n989), .B2(new_n996), .ZN(new_n997));
  NOR2_X1   g572(.A1(G166), .A2(new_n968), .ZN(new_n998));
  XOR2_X1   g573(.A(KEYINPUT114), .B(KEYINPUT55), .Z(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n1001));
  OAI22_X1  g576(.A1(G166), .A2(new_n968), .B1(KEYINPUT114), .B2(new_n1001), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n997), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n986), .A2(new_n982), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1006), .B(new_n965), .C1(new_n962), .C2(new_n982), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n1007), .A2(G2090), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1008), .A2(KEYINPUT118), .A3(new_n996), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(G8), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT118), .B1(new_n1008), .B2(new_n996), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1003), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n984), .A2(new_n778), .A3(new_n965), .A4(new_n988), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n980), .A2(new_n992), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1014), .B(new_n965), .C1(new_n992), .C2(new_n991), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n815), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n968), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n1017), .A2(new_n596), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n977), .A2(new_n1005), .A3(new_n1012), .A4(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT63), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1005), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT63), .B1(new_n997), .B2(new_n1004), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n976), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n1019), .A2(new_n1020), .B1(new_n1023), .B2(new_n1018), .ZN(new_n1024));
  NOR2_X1   g599(.A1(G168), .A2(new_n968), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1025), .B1(new_n1017), .B2(KEYINPUT123), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1017), .A2(KEYINPUT123), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT51), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT51), .B1(new_n1030), .B2(G8), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1025), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT124), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT124), .ZN(new_n1034));
  NOR4_X1   g609(.A1(new_n1017), .A2(new_n1034), .A3(KEYINPUT51), .A4(new_n1025), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n1029), .A2(new_n1036), .B1(new_n1030), .B2(new_n1025), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n984), .A2(new_n965), .A3(new_n988), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n819), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1040), .B1(new_n994), .B2(G2078), .ZN(new_n1041));
  NAND2_X1  g616(.A1(G160), .A2(G40), .ZN(new_n1042));
  OAI211_X1 g617(.A(KEYINPUT53), .B(new_n746), .C1(new_n1042), .C2(KEYINPUT125), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1043), .B1(KEYINPUT125), .B2(new_n1042), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1044), .A2(new_n1014), .A3(new_n990), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1039), .A2(new_n1041), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(G171), .ZN(new_n1047));
  OR3_X1    g622(.A1(new_n1015), .A2(new_n1040), .A3(G2078), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1048), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1047), .B(KEYINPUT54), .C1(G171), .C2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n977), .A2(new_n1050), .A3(new_n1005), .A4(new_n1012), .ZN(new_n1051));
  OR2_X1    g626(.A1(new_n1046), .A2(G171), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1049), .A2(G171), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT54), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NOR3_X1   g629(.A1(new_n1037), .A2(new_n1051), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n806), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1038), .A2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n966), .A2(G2067), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT120), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT120), .ZN(new_n1061));
  AOI211_X1 g636(.A(new_n1061), .B(new_n1058), .C1(new_n1038), .C2(new_n1056), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(G1956), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1007), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT119), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n585), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1071));
  XNOR2_X1  g646(.A(KEYINPUT56), .B(G2072), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n990), .A2(new_n993), .A3(new_n965), .A4(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1065), .A2(new_n1070), .A3(new_n1071), .A4(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1063), .A2(new_n632), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1065), .A2(new_n1073), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1071), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1076), .B1(new_n1069), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n1074), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT61), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n1082));
  INV_X1    g657(.A(G1996), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n990), .A2(new_n993), .A3(new_n1083), .A4(new_n965), .ZN(new_n1084));
  XOR2_X1   g659(.A(KEYINPUT58), .B(G1341), .Z(new_n1085));
  NAND2_X1  g660(.A1(new_n966), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n563), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT121), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1082), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1089), .B1(new_n1088), .B2(new_n1087), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1078), .A2(KEYINPUT61), .A3(new_n1074), .ZN(new_n1091));
  OR3_X1    g666(.A1(new_n1087), .A2(new_n1088), .A3(KEYINPUT59), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1081), .A2(new_n1090), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT122), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1095));
  XNOR2_X1  g670(.A(new_n1089), .B(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT122), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1096), .A2(new_n1097), .A3(new_n1081), .A4(new_n1091), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1094), .A2(new_n1098), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n1060), .A2(new_n1062), .A3(KEYINPUT60), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT60), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n632), .B1(new_n1063), .B2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g677(.A(KEYINPUT60), .B(new_n879), .C1(new_n1060), .C2(new_n1062), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1100), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1075), .B(new_n1078), .C1(new_n1099), .C2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1024), .B1(new_n1055), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n977), .A2(new_n1005), .A3(new_n1012), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT62), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1108), .B1(new_n1037), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1030), .A2(new_n1025), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n1034), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1031), .A2(KEYINPUT124), .A3(new_n1032), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT51), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1028), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1116), .B1(new_n1117), .B2(new_n1026), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1109), .B(new_n1111), .C1(new_n1115), .C2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1053), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(KEYINPUT126), .B1(new_n1110), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1111), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1107), .B1(new_n1123), .B2(KEYINPUT62), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT126), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1124), .A2(new_n1125), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n970), .A2(new_n971), .A3(new_n714), .ZN(new_n1127));
  INV_X1    g702(.A(new_n951), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n969), .B(KEYINPUT116), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n1129), .A2(new_n1130), .B1(new_n977), .B2(new_n1021), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT117), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n1131), .B(new_n1132), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1106), .A2(new_n1122), .A3(new_n1126), .A4(new_n1133), .ZN(new_n1134));
  OR2_X1    g709(.A1(new_n734), .A2(new_n738), .ZN(new_n1135));
  INV_X1    g710(.A(G2067), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n795), .B(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n764), .A2(G1996), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n765), .A2(new_n1083), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1135), .A2(new_n1137), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1140), .B1(new_n738), .B2(new_n734), .ZN(new_n1141));
  OR2_X1    g716(.A1(G290), .A2(G1986), .ZN(new_n1142));
  NAND2_X1  g717(.A1(G290), .A2(G1986), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1014), .A2(new_n964), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1134), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1145), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1148), .B1(new_n765), .B2(new_n1137), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1145), .A2(KEYINPUT46), .A3(new_n1083), .ZN(new_n1150));
  AOI21_X1  g725(.A(KEYINPUT46), .B1(new_n1145), .B2(new_n1083), .ZN(new_n1151));
  NOR3_X1   g726(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  XOR2_X1   g727(.A(new_n1152), .B(KEYINPUT47), .Z(new_n1153));
  NOR2_X1   g728(.A1(new_n1148), .A2(new_n1142), .ZN(new_n1154));
  XOR2_X1   g729(.A(new_n1154), .B(KEYINPUT48), .Z(new_n1155));
  OAI21_X1  g730(.A(new_n1155), .B1(new_n1148), .B2(new_n1141), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1139), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1157));
  OAI22_X1  g732(.A1(new_n1135), .A2(new_n1157), .B1(G2067), .B2(new_n795), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(new_n1145), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1153), .A2(new_n1156), .A3(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(KEYINPUT127), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1147), .A2(new_n1161), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g737(.A(G319), .ZN(new_n1164));
  NOR2_X1   g738(.A1(G229), .A2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g739(.A1(G227), .A2(G401), .ZN(new_n1166));
  AND2_X1   g740(.A1(new_n872), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g741(.A1(new_n946), .A2(new_n1165), .A3(new_n1167), .ZN(G225));
  INV_X1    g742(.A(G225), .ZN(G308));
endmodule


