//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 1 0 1 0 0 1 0 0 0 1 1 1 1 0 0 1 1 1 1 0 1 1 1 1 1 0 1 0 1 0 0 0 1 1 0 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n598, new_n599, new_n600, new_n601,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937;
  INV_X1    g000(.A(G116), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT69), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT69), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G116), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G119), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n187), .A2(G119), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT2), .B(G113), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT70), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n193), .B1(new_n191), .B2(G119), .ZN(new_n199));
  INV_X1    g013(.A(G113), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT2), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT2), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G113), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n198), .B1(new_n199), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G119), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n206), .B1(new_n188), .B2(new_n190), .ZN(new_n207));
  NOR4_X1   g021(.A1(new_n207), .A2(new_n196), .A3(KEYINPUT70), .A4(new_n193), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n197), .B1(new_n205), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT71), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT69), .B(G116), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n204), .B(new_n194), .C1(new_n211), .C2(new_n206), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT70), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n192), .A2(new_n198), .A3(new_n194), .A4(new_n204), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT71), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n216), .A3(new_n197), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n210), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G146), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(KEYINPUT66), .A3(G143), .ZN(new_n220));
  INV_X1    g034(.A(G128), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n223));
  INV_X1    g037(.A(G143), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n223), .B1(new_n224), .B2(G146), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n224), .A2(G146), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n220), .B(new_n222), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT68), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n219), .A2(G143), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n219), .A2(G143), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n229), .B1(new_n230), .B2(new_n223), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n231), .A2(new_n232), .A3(new_n220), .A4(new_n222), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n224), .A2(G146), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n229), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT1), .ZN(new_n236));
  OAI21_X1  g050(.A(G128), .B1(new_n226), .B2(new_n236), .ZN(new_n237));
  AOI22_X1  g051(.A1(new_n228), .A2(new_n233), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G137), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(G134), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G131), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT11), .ZN(new_n243));
  INV_X1    g057(.A(G134), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n243), .B1(new_n244), .B2(G137), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n239), .A2(KEYINPUT11), .A3(G134), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n241), .A2(new_n242), .A3(new_n245), .A4(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n244), .A2(G137), .ZN(new_n248));
  OAI21_X1  g062(.A(G131), .B1(new_n240), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n245), .A2(new_n246), .ZN(new_n251));
  OAI21_X1  g065(.A(G131), .B1(new_n251), .B2(new_n240), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n247), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT0), .ZN(new_n255));
  AOI21_X1  g069(.A(KEYINPUT65), .B1(new_n255), .B2(new_n221), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT65), .ZN(new_n257));
  NOR3_X1   g071(.A1(new_n257), .A2(KEYINPUT0), .A3(G128), .ZN(new_n258));
  OAI221_X1 g072(.A(new_n235), .B1(new_n255), .B2(new_n221), .C1(new_n256), .C2(new_n258), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n231), .A2(KEYINPUT0), .A3(G128), .A4(new_n220), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI22_X1  g075(.A1(new_n238), .A2(new_n250), .B1(new_n254), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n218), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n259), .A2(new_n260), .A3(KEYINPUT67), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(new_n253), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT67), .B1(new_n259), .B2(new_n260), .ZN(new_n266));
  OAI22_X1  g080(.A1(new_n265), .A2(new_n266), .B1(new_n238), .B2(new_n250), .ZN(new_n267));
  XOR2_X1   g081(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n268));
  NAND2_X1  g082(.A1(new_n228), .A2(new_n233), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n237), .A2(new_n235), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n250), .ZN(new_n272));
  INV_X1    g086(.A(new_n261), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n271), .A2(new_n272), .B1(new_n273), .B2(new_n253), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n267), .A2(new_n268), .B1(new_n274), .B2(KEYINPUT30), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n263), .B1(new_n275), .B2(new_n218), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT74), .ZN(new_n277));
  NOR2_X1   g091(.A1(G237), .A2(G953), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G210), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n279), .B(KEYINPUT73), .ZN(new_n280));
  XOR2_X1   g094(.A(KEYINPUT26), .B(G101), .Z(new_n281));
  XNOR2_X1  g095(.A(new_n280), .B(new_n281), .ZN(new_n282));
  XNOR2_X1  g096(.A(KEYINPUT72), .B(KEYINPUT27), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n282), .B(new_n283), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n276), .A2(new_n277), .A3(KEYINPUT31), .A4(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n267), .A2(new_n268), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n274), .A2(KEYINPUT30), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n287), .A3(new_n218), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n215), .A2(new_n216), .A3(new_n197), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n216), .B1(new_n215), .B2(new_n197), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n274), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n288), .A2(new_n277), .A3(new_n292), .A4(new_n284), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT31), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n285), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT28), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n297), .B1(new_n218), .B2(new_n262), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n291), .A2(KEYINPUT28), .A3(new_n274), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n218), .A2(new_n267), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n284), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n296), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT32), .ZN(new_n306));
  NOR2_X1   g120(.A1(G472), .A2(G902), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  AOI22_X1  g122(.A1(new_n285), .A2(new_n295), .B1(new_n302), .B2(new_n303), .ZN(new_n309));
  INV_X1    g123(.A(new_n307), .ZN(new_n310));
  OAI21_X1  g124(.A(KEYINPUT32), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT76), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n313), .B1(new_n218), .B2(new_n262), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n298), .A2(new_n314), .A3(new_n299), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n263), .A2(new_n313), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n303), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(G902), .B1(new_n317), .B2(KEYINPUT29), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT75), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n300), .A2(new_n319), .A3(new_n301), .A4(new_n284), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n288), .A2(new_n292), .ZN(new_n321));
  AOI21_X1  g135(.A(KEYINPUT29), .B1(new_n321), .B2(new_n303), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n298), .A2(new_n299), .A3(new_n284), .A4(new_n301), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT75), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n320), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n318), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g140(.A(KEYINPUT77), .B1(new_n326), .B2(G472), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT77), .ZN(new_n328));
  INV_X1    g142(.A(G472), .ZN(new_n329));
  AOI211_X1 g143(.A(new_n328), .B(new_n329), .C1(new_n318), .C2(new_n325), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n312), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(G214), .B1(G237), .B2(G902), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  XOR2_X1   g147(.A(G110), .B(G122), .Z(new_n334));
  INV_X1    g148(.A(G104), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT3), .B1(new_n335), .B2(G107), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT3), .ZN(new_n337));
  INV_X1    g151(.A(G107), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(new_n338), .A3(G104), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n335), .A2(G107), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n336), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G101), .ZN(new_n342));
  INV_X1    g156(.A(G101), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n336), .A2(new_n339), .A3(new_n343), .A4(new_n340), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n342), .A2(KEYINPUT80), .A3(KEYINPUT4), .A4(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(KEYINPUT80), .A2(KEYINPUT4), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n341), .A2(G101), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n348), .B1(new_n210), .B2(new_n217), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT5), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n193), .A2(new_n350), .ZN(new_n351));
  OAI211_X1 g165(.A(G113), .B(new_n351), .C1(new_n195), .C2(new_n350), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n215), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT81), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n354), .B1(new_n335), .B2(G107), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n338), .A2(KEYINPUT81), .A3(G104), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n355), .A2(new_n340), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G101), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n344), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT82), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT84), .ZN(new_n361));
  AOI21_X1  g175(.A(KEYINPUT82), .B1(new_n357), .B2(G101), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n360), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT82), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n365), .B1(new_n358), .B2(new_n344), .ZN(new_n366));
  OAI21_X1  g180(.A(KEYINPUT84), .B1(new_n366), .B2(new_n362), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n353), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n334), .B1(new_n349), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n348), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n370), .B1(new_n289), .B2(new_n290), .ZN(new_n371));
  INV_X1    g185(.A(new_n334), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n352), .A2(new_n215), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n361), .B1(new_n360), .B2(new_n363), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n366), .A2(KEYINPUT84), .A3(new_n362), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n371), .A2(new_n372), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n369), .A2(KEYINPUT6), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT6), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n379), .B(new_n334), .C1(new_n349), .C2(new_n368), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n271), .A2(G125), .ZN(new_n381));
  INV_X1    g195(.A(G125), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n273), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G224), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(G953), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n386), .B(KEYINPUT85), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n384), .B(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n378), .A2(new_n380), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G902), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n360), .A2(new_n363), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n373), .A2(new_n391), .ZN(new_n392));
  XOR2_X1   g206(.A(new_n334), .B(KEYINPUT8), .Z(new_n393));
  NOR2_X1   g207(.A1(new_n366), .A2(new_n362), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n353), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n392), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT86), .ZN(new_n397));
  OAI22_X1  g211(.A1(new_n381), .A2(new_n383), .B1(KEYINPUT87), .B2(new_n386), .ZN(new_n398));
  OAI21_X1  g212(.A(KEYINPUT7), .B1(new_n385), .B2(G953), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  AOI22_X1  g214(.A1(new_n396), .A2(new_n397), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  OR2_X1    g215(.A1(new_n398), .A2(new_n400), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n392), .A2(KEYINPUT86), .A3(new_n393), .A4(new_n395), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n401), .A2(new_n402), .A3(new_n403), .A4(new_n377), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n389), .A2(new_n390), .A3(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(G210), .B1(G237), .B2(G902), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n389), .A2(new_n404), .A3(new_n390), .A4(new_n406), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n333), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  XOR2_X1   g224(.A(KEYINPUT9), .B(G234), .Z(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(G221), .B1(new_n412), .B2(G902), .ZN(new_n413));
  INV_X1    g227(.A(G469), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n231), .A2(new_n220), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n237), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n269), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(KEYINPUT10), .B1(new_n417), .B2(new_n394), .ZN(new_n418));
  AOI22_X1  g232(.A1(new_n418), .A2(KEYINPUT83), .B1(new_n273), .B2(new_n370), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT83), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n228), .A2(new_n233), .B1(new_n415), .B2(new_n237), .ZN(new_n421));
  NOR3_X1   g235(.A1(new_n421), .A2(new_n366), .A3(new_n362), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n420), .B1(new_n422), .B2(KEYINPUT10), .ZN(new_n423));
  OAI211_X1 g237(.A(KEYINPUT10), .B(new_n271), .C1(new_n374), .C2(new_n375), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n419), .A2(new_n254), .A3(new_n423), .A4(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(G110), .B(G140), .ZN(new_n426));
  INV_X1    g240(.A(G953), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G227), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n426), .B(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n391), .A2(new_n238), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n417), .A2(new_n394), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n254), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT12), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n433), .B(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n430), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n418), .A2(KEYINPUT83), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n370), .A2(new_n273), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n423), .A2(new_n437), .A3(new_n424), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n253), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n429), .B1(new_n440), .B2(new_n425), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n414), .B(new_n390), .C1(new_n436), .C2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(G469), .A2(G902), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n429), .B(KEYINPUT79), .ZN(new_n444));
  INV_X1    g258(.A(new_n425), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n444), .B1(new_n445), .B2(new_n435), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n440), .A2(new_n425), .A3(new_n429), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(G469), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n442), .A2(new_n443), .A3(new_n448), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n410), .A2(new_n413), .A3(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(G125), .B(G140), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT16), .ZN(new_n452));
  OR3_X1    g266(.A1(new_n382), .A2(KEYINPUT16), .A3(G140), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n219), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n452), .A2(G146), .A3(new_n453), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n206), .A2(G128), .ZN(new_n458));
  OR2_X1    g272(.A1(new_n458), .A2(KEYINPUT23), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n206), .A2(G128), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n458), .A2(KEYINPUT23), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(G110), .ZN(new_n463));
  INV_X1    g277(.A(new_n460), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(new_n458), .ZN(new_n465));
  XOR2_X1   g279(.A(KEYINPUT24), .B(G110), .Z(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n457), .A2(new_n463), .A3(new_n467), .ZN(new_n468));
  OAI22_X1  g282(.A1(new_n462), .A2(G110), .B1(new_n465), .B2(new_n466), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n451), .A2(new_n219), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n469), .A2(new_n456), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n427), .A2(G221), .A3(G234), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(G137), .ZN(new_n474));
  XNOR2_X1  g288(.A(KEYINPUT78), .B(KEYINPUT22), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n474), .B(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n472), .B(new_n476), .ZN(new_n477));
  OR3_X1    g291(.A1(new_n477), .A2(KEYINPUT25), .A3(G902), .ZN(new_n478));
  INV_X1    g292(.A(G217), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n479), .B1(G234), .B2(new_n390), .ZN(new_n480));
  OAI21_X1  g294(.A(KEYINPUT25), .B1(new_n477), .B2(G902), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  OR3_X1    g296(.A1(new_n477), .A2(G902), .A3(new_n480), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(G122), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n211), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n187), .A2(G122), .ZN(new_n488));
  OAI21_X1  g302(.A(G107), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n488), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n338), .B(new_n490), .C1(new_n211), .C2(new_n486), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT91), .ZN(new_n493));
  XNOR2_X1  g307(.A(G128), .B(G143), .ZN(new_n494));
  AOI22_X1  g308(.A1(new_n492), .A2(new_n493), .B1(new_n244), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(KEYINPUT13), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n224), .A2(G128), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n496), .B(G134), .C1(KEYINPUT13), .C2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n489), .A2(KEYINPUT91), .A3(new_n491), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n495), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(KEYINPUT92), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT92), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n495), .A2(new_n502), .A3(new_n498), .A4(new_n499), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n494), .B(new_n244), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT14), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n490), .B1(new_n487), .B2(new_n506), .ZN(new_n507));
  OR2_X1    g321(.A1(new_n507), .A2(KEYINPUT93), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n487), .A2(new_n506), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n507), .A2(KEYINPUT93), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n491), .B(new_n505), .C1(new_n511), .C2(new_n338), .ZN(new_n512));
  NOR3_X1   g326(.A1(new_n412), .A2(new_n479), .A3(G953), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n504), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n513), .B1(new_n504), .B2(new_n512), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n390), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT15), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n517), .A3(G478), .ZN(new_n518));
  INV_X1    g332(.A(G478), .ZN(new_n519));
  OAI221_X1 g333(.A(new_n390), .B1(KEYINPUT15), .B2(new_n519), .C1(new_n514), .C2(new_n515), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n457), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n278), .A2(G214), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n523), .A2(KEYINPUT88), .A3(G143), .ZN(new_n524));
  OR2_X1    g338(.A1(KEYINPUT88), .A2(G143), .ZN(new_n525));
  NAND2_X1  g339(.A1(KEYINPUT88), .A2(G143), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n525), .A2(G214), .A3(new_n278), .A4(new_n526), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n524), .A2(new_n527), .A3(KEYINPUT17), .A4(G131), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n524), .A2(new_n527), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(new_n242), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n522), .B(new_n528), .C1(new_n530), .C2(KEYINPUT17), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT90), .ZN(new_n532));
  NAND2_X1  g346(.A1(KEYINPUT18), .A2(G131), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT89), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n529), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n524), .A2(new_n535), .A3(new_n527), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n451), .B(new_n219), .ZN(new_n539));
  NAND3_X1  g353(.A1(KEYINPUT90), .A2(KEYINPUT18), .A3(G131), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n537), .A2(new_n538), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n531), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g356(.A(G113), .B(G122), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(new_n335), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n542), .B(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(G475), .B1(new_n545), .B2(G902), .ZN(new_n546));
  XOR2_X1   g360(.A(new_n451), .B(KEYINPUT19), .Z(new_n547));
  OAI211_X1 g361(.A(new_n530), .B(new_n456), .C1(G146), .C2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n541), .ZN(new_n549));
  INV_X1    g363(.A(new_n544), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n531), .A2(new_n544), .A3(new_n541), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(G475), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n553), .A2(new_n554), .A3(new_n390), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT20), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n553), .A2(KEYINPUT20), .A3(new_n554), .A4(new_n390), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n546), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(G234), .A2(G237), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n560), .A2(G902), .A3(G953), .ZN(new_n561));
  XOR2_X1   g375(.A(new_n561), .B(KEYINPUT94), .Z(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT21), .B(G898), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n427), .A2(G952), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n565), .B1(G234), .B2(G237), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NOR3_X1   g381(.A1(new_n521), .A2(new_n559), .A3(new_n567), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n331), .A2(new_n450), .A3(new_n485), .A4(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(G101), .ZN(G3));
  AOI211_X1 g384(.A(new_n333), .B(new_n567), .C1(new_n408), .C2(new_n409), .ZN(new_n571));
  OAI21_X1  g385(.A(KEYINPUT33), .B1(new_n514), .B2(new_n515), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n504), .A2(new_n512), .ZN(new_n573));
  INV_X1    g387(.A(new_n513), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT33), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n504), .A2(new_n512), .A3(new_n513), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n572), .A2(new_n578), .A3(G478), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n519), .A2(new_n390), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n519), .B(new_n390), .C1(new_n514), .C2(new_n515), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n579), .A2(new_n559), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  AND3_X1   g398(.A1(new_n571), .A2(new_n584), .A3(KEYINPUT95), .ZN(new_n585));
  AOI21_X1  g399(.A(KEYINPUT95), .B1(new_n571), .B2(new_n584), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n449), .A2(new_n413), .ZN(new_n589));
  OAI21_X1  g403(.A(G472), .B1(new_n309), .B2(G902), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n305), .A2(new_n307), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n589), .A2(new_n592), .A3(new_n484), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(new_n335), .ZN(new_n595));
  XOR2_X1   g409(.A(KEYINPUT96), .B(KEYINPUT34), .Z(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(G6));
  AOI21_X1  g411(.A(new_n559), .B1(new_n518), .B2(new_n520), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n593), .A2(new_n571), .A3(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(new_n338), .ZN(new_n600));
  XNOR2_X1  g414(.A(KEYINPUT97), .B(KEYINPUT35), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(G9));
  NOR2_X1   g416(.A1(new_n476), .A2(KEYINPUT36), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n472), .B(new_n603), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n604), .B(new_n390), .C1(new_n479), .C2(G234), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n482), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n590), .A2(new_n591), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT98), .ZN(new_n608));
  OR2_X1    g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n607), .A2(new_n608), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n609), .A2(new_n450), .A3(new_n568), .A4(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT37), .B(G110), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G12));
  INV_X1    g427(.A(new_n559), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n521), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(G900), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n566), .B1(new_n562), .B2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(KEYINPUT99), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n331), .A2(new_n450), .A3(new_n606), .A4(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT100), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G128), .ZN(G30));
  AND2_X1   g437(.A1(new_n449), .A2(new_n413), .ZN(new_n624));
  XOR2_X1   g438(.A(new_n618), .B(KEYINPUT39), .Z(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(new_n626), .B(KEYINPUT40), .Z(new_n627));
  INV_X1    g441(.A(new_n606), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n408), .A2(new_n409), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n312), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n316), .A2(new_n303), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n314), .A2(new_n292), .ZN(new_n634));
  OAI22_X1  g448(.A1(new_n633), .A2(new_n634), .B1(new_n321), .B2(new_n303), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n329), .B1(new_n635), .B2(new_n390), .ZN(new_n636));
  XOR2_X1   g450(.A(new_n636), .B(KEYINPUT102), .Z(new_n637));
  NOR2_X1   g451(.A1(new_n632), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n614), .B1(new_n518), .B2(new_n520), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n638), .A2(new_n333), .A3(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n627), .A2(new_n628), .A3(new_n631), .A4(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G143), .ZN(G45));
  AND2_X1   g457(.A1(new_n331), .A2(new_n606), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n583), .A2(new_n618), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n644), .A2(new_n450), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G146), .ZN(G48));
  NOR2_X1   g461(.A1(new_n436), .A2(new_n441), .ZN(new_n648));
  OAI21_X1  g462(.A(G469), .B1(new_n648), .B2(G902), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n649), .A2(new_n413), .A3(new_n442), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n331), .A2(new_n485), .A3(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n588), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT41), .B(G113), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G15));
  NAND3_X1  g470(.A1(new_n653), .A2(new_n571), .A3(new_n598), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G116), .ZN(G18));
  AND2_X1   g472(.A1(new_n408), .A2(new_n409), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n650), .A2(new_n659), .A3(new_n333), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n660), .A2(new_n331), .A3(new_n568), .A4(new_n606), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G119), .ZN(G21));
  NOR2_X1   g476(.A1(new_n640), .A2(new_n650), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n329), .B1(new_n305), .B2(new_n390), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n315), .A2(new_n303), .A3(new_n316), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n310), .B1(new_n296), .B2(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(KEYINPUT103), .B1(new_n667), .B2(new_n485), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT103), .ZN(new_n669));
  NOR4_X1   g483(.A1(new_n664), .A2(new_n666), .A3(new_n484), .A4(new_n669), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n663), .B(new_n571), .C1(new_n668), .C2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G122), .ZN(G24));
  NOR3_X1   g486(.A1(new_n664), .A2(new_n628), .A3(new_n666), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n660), .A2(new_n645), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G125), .ZN(G27));
  NAND2_X1  g489(.A1(new_n659), .A2(new_n332), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n676), .A2(new_n589), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n677), .A2(new_n485), .A3(new_n331), .A4(new_n645), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT42), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G131), .ZN(G33));
  AND2_X1   g495(.A1(new_n331), .A2(new_n485), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n682), .A2(new_n619), .A3(new_n677), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G134), .ZN(G36));
  AND2_X1   g498(.A1(new_n579), .A2(new_n582), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n614), .A3(new_n581), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(KEYINPUT43), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(KEYINPUT106), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n688), .A2(new_n693), .A3(new_n690), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n692), .A2(new_n592), .A3(new_n606), .A4(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n697), .A2(new_n676), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n446), .A2(new_n447), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT45), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n446), .A2(KEYINPUT45), .A3(new_n447), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n701), .A2(G469), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(KEYINPUT104), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n443), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT46), .ZN(new_n706));
  OAI21_X1  g520(.A(KEYINPUT105), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n705), .A2(new_n706), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT105), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n704), .A2(new_n709), .A3(KEYINPUT46), .A4(new_n443), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n707), .A2(new_n708), .A3(new_n442), .A4(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n413), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n695), .A2(new_n696), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n698), .A2(new_n625), .A3(new_n713), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(KEYINPUT107), .B(G137), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G39));
  NOR2_X1   g531(.A1(new_n629), .A2(new_n333), .ZN(new_n718));
  OR4_X1    g532(.A1(new_n485), .A2(new_n331), .A3(new_n583), .A4(new_n618), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n711), .A2(KEYINPUT47), .A3(new_n413), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(KEYINPUT47), .B1(new_n711), .B2(new_n413), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n718), .B(new_n720), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT108), .B(G140), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G42));
  INV_X1    g540(.A(KEYINPUT49), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n649), .A2(new_n442), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n687), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n729), .B1(new_n727), .B2(new_n728), .ZN(new_n730));
  INV_X1    g544(.A(new_n638), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(new_n484), .ZN(new_n732));
  INV_X1    g546(.A(new_n413), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n631), .A2(new_n333), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n730), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT53), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n598), .B1(new_n583), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n738), .B1(new_n737), .B2(new_n583), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(new_n571), .A3(new_n593), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n569), .A3(new_n611), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT110), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT110), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n740), .A2(new_n611), .A3(new_n743), .A4(new_n569), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n659), .A2(new_n332), .A3(new_n614), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n521), .A2(new_n618), .ZN(new_n747));
  OAI21_X1  g561(.A(KEYINPUT111), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n521), .A2(new_n618), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT111), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n718), .A2(new_n749), .A3(new_n750), .A4(new_n614), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n624), .A3(new_n644), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n677), .A2(new_n645), .A3(new_n673), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(new_n683), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(KEYINPUT112), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT112), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n753), .A2(new_n757), .A3(new_n683), .A4(new_n754), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n745), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n671), .B(new_n661), .C1(new_n587), .C2(new_n652), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n653), .A2(new_n571), .A3(new_n598), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n680), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n620), .A2(new_n621), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n620), .A2(new_n621), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n674), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(KEYINPUT113), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n640), .A2(new_n333), .A3(new_n659), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n589), .A2(new_n606), .A3(new_n618), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n731), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n771), .A2(KEYINPUT52), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n773), .B(new_n674), .C1(new_n765), .C2(new_n766), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n768), .A2(new_n646), .A3(new_n772), .A4(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n622), .A2(new_n646), .A3(new_n674), .A4(new_n771), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n775), .A2(new_n776), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n776), .B1(new_n775), .B2(new_n779), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n736), .B(new_n764), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n772), .A2(new_n622), .A3(new_n646), .A4(new_n674), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n764), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(KEYINPUT53), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n782), .A2(KEYINPUT54), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT115), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n760), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n790), .A2(new_n791), .A3(new_n680), .A4(new_n657), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(KEYINPUT53), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n791), .B1(new_n762), .B2(new_n680), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n793), .A2(new_n759), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n795), .B1(new_n780), .B2(new_n781), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n785), .A2(new_n736), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n788), .B1(new_n787), .B2(new_n799), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n651), .A2(new_n566), .A3(new_n718), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n732), .A2(new_n584), .A3(new_n801), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n691), .A2(new_n801), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n682), .ZN(new_n804));
  XOR2_X1   g618(.A(new_n804), .B(KEYINPUT48), .Z(new_n805));
  OR2_X1    g619(.A1(new_n668), .A2(new_n670), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n806), .A2(new_n566), .A3(new_n691), .ZN(new_n807));
  AOI211_X1 g621(.A(new_n565), .B(new_n805), .C1(new_n660), .C2(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n631), .A2(new_n650), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n807), .A2(new_n333), .A3(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT118), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT50), .ZN(new_n812));
  OAI21_X1  g626(.A(KEYINPUT117), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n815));
  AOI22_X1  g629(.A1(new_n803), .A2(new_n673), .B1(KEYINPUT119), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n685), .A2(new_n581), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n732), .A2(new_n614), .A3(new_n817), .A4(new_n801), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n814), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n820));
  OAI21_X1  g634(.A(KEYINPUT118), .B1(new_n810), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n819), .B1(new_n812), .B2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n723), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n728), .A2(new_n733), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(new_n721), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n825), .A2(new_n718), .A3(new_n807), .ZN(new_n826));
  OR2_X1    g640(.A1(new_n815), .A2(KEYINPUT119), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n822), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n827), .B1(new_n822), .B2(new_n826), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n808), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NOR4_X1   g644(.A1(new_n789), .A2(new_n800), .A3(new_n802), .A4(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(G952), .A2(G953), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n735), .B1(new_n831), .B2(new_n832), .ZN(G75));
  INV_X1    g647(.A(new_n759), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n763), .A2(KEYINPUT116), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n834), .A2(new_n835), .A3(KEYINPUT53), .A4(new_n792), .ZN(new_n836));
  INV_X1    g650(.A(new_n781), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n775), .A2(new_n776), .A3(new_n779), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT53), .B1(new_n764), .B2(new_n784), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n390), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT56), .B1(new_n842), .B2(G210), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n378), .A2(new_n380), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(new_n388), .ZN(new_n845));
  XNOR2_X1  g659(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n846));
  XOR2_X1   g660(.A(new_n845), .B(new_n846), .Z(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n843), .A2(new_n848), .ZN(new_n849));
  AOI211_X1 g663(.A(KEYINPUT56), .B(new_n847), .C1(new_n842), .C2(G210), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n427), .A2(G952), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(G51));
  INV_X1    g666(.A(KEYINPUT122), .ZN(new_n853));
  AOI211_X1 g667(.A(new_n390), .B(new_n704), .C1(new_n796), .C2(new_n798), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n443), .B(KEYINPUT121), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(KEYINPUT57), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n797), .B1(new_n796), .B2(new_n798), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n648), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n854), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n853), .B1(new_n861), .B2(new_n851), .ZN(new_n862));
  INV_X1    g676(.A(new_n851), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT54), .B1(new_n839), .B2(new_n840), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(new_n799), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n648), .B1(new_n865), .B2(new_n856), .ZN(new_n866));
  OAI211_X1 g680(.A(KEYINPUT122), .B(new_n863), .C1(new_n866), .C2(new_n854), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n862), .A2(new_n867), .ZN(G54));
  NAND3_X1  g682(.A1(new_n842), .A2(KEYINPUT58), .A3(G475), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n869), .A2(new_n552), .A3(new_n551), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n842), .A2(KEYINPUT58), .A3(G475), .A4(new_n553), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n870), .A2(new_n863), .A3(new_n871), .ZN(G60));
  AND2_X1   g686(.A1(new_n572), .A2(new_n578), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n580), .B(KEYINPUT59), .ZN(new_n874));
  AOI211_X1 g688(.A(new_n873), .B(new_n874), .C1(new_n864), .C2(new_n799), .ZN(new_n875));
  INV_X1    g689(.A(new_n874), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n876), .B1(new_n789), .B2(new_n800), .ZN(new_n877));
  AOI211_X1 g691(.A(new_n851), .B(new_n875), .C1(new_n877), .C2(new_n873), .ZN(G63));
  NAND2_X1  g692(.A1(G217), .A2(G902), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT60), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n477), .B1(new_n841), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n880), .B1(new_n796), .B2(new_n798), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n851), .B1(new_n882), .B2(new_n604), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT123), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT61), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n884), .B(new_n885), .ZN(G66));
  OAI21_X1  g700(.A(G953), .B1(new_n563), .B2(new_n385), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n745), .A2(new_n762), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n887), .B1(new_n889), .B2(G953), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n844), .B1(G898), .B2(new_n427), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n890), .B(new_n891), .ZN(G69));
  XNOR2_X1  g706(.A(new_n275), .B(KEYINPUT124), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(new_n547), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n739), .B(KEYINPUT125), .Z(new_n895));
  AND4_X1   g709(.A1(new_n682), .A2(new_n895), .A3(new_n625), .A4(new_n677), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n768), .A2(new_n774), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n897), .A2(new_n646), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n898), .A2(KEYINPUT62), .A3(new_n642), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n897), .A2(new_n642), .A3(new_n646), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT62), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n896), .B1(new_n899), .B2(new_n902), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n715), .A2(new_n724), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n894), .B1(new_n905), .B2(G953), .ZN(new_n906));
  INV_X1    g720(.A(G227), .ZN(new_n907));
  OAI21_X1  g721(.A(G953), .B1(new_n907), .B2(new_n616), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(KEYINPUT126), .ZN(new_n909));
  OR2_X1    g723(.A1(new_n908), .A2(KEYINPUT126), .ZN(new_n910));
  INV_X1    g724(.A(new_n894), .ZN(new_n911));
  NAND2_X1  g725(.A1(G900), .A2(G953), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n711), .A2(new_n682), .A3(new_n413), .A4(new_n625), .ZN(new_n913));
  INV_X1    g727(.A(new_n769), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n680), .B(new_n683), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n904), .A2(new_n898), .A3(new_n916), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n911), .B(new_n912), .C1(new_n917), .C2(G953), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n906), .A2(new_n909), .A3(new_n910), .A4(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n903), .A2(new_n904), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n911), .B1(new_n920), .B2(new_n427), .ZN(new_n921));
  INV_X1    g735(.A(new_n918), .ZN(new_n922));
  OAI211_X1 g736(.A(KEYINPUT126), .B(new_n908), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n919), .A2(new_n923), .ZN(G72));
  NAND2_X1  g738(.A1(G472), .A2(G902), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT63), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n927), .B1(new_n917), .B2(new_n888), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n928), .A2(new_n303), .A3(new_n276), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n321), .B(new_n303), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n782), .A2(new_n786), .A3(new_n927), .A4(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n929), .A2(new_n863), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n926), .B1(new_n905), .B2(new_n889), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT127), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n303), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n927), .B1(new_n920), .B2(new_n888), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n276), .B1(new_n936), .B2(KEYINPUT127), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n932), .B1(new_n935), .B2(new_n937), .ZN(G57));
endmodule


