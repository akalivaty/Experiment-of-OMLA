//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 1 1 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 1 1 0 0 0 0 1 1 0 0 0 1 1 1 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n559, new_n560, new_n562, new_n563, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n580, new_n581, new_n582,
    new_n583, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1140, new_n1141, new_n1142;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n452));
  XOR2_X1   g027(.A(new_n451), .B(new_n452), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(G325));
  XOR2_X1   g031(.A(new_n455), .B(KEYINPUT66), .Z(G261));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  AOI22_X1  g034(.A1(new_n458), .A2(G2106), .B1(G567), .B2(new_n459), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n464), .A2(new_n466), .A3(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n464), .A2(new_n466), .A3(G137), .A4(new_n462), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n469), .A2(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n464), .A2(new_n466), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G136), .ZN(new_n476));
  OAI21_X1  g051(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n462), .A2(G112), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n474), .A2(new_n462), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n479), .B1(G124), .B2(new_n480), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT68), .ZN(G162));
  NAND4_X1  g057(.A1(new_n464), .A2(new_n466), .A3(G126), .A4(G2105), .ZN(new_n483));
  OR2_X1    g058(.A1(G102), .A2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G114), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n484), .A2(new_n486), .A3(G2104), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n462), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  XNOR2_X1  g065(.A(KEYINPUT3), .B(G2104), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n491), .A2(new_n492), .A3(G138), .A4(new_n462), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n488), .B1(new_n490), .B2(new_n493), .ZN(G164));
  INV_X1    g069(.A(KEYINPUT6), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G651), .ZN(new_n496));
  INV_X1    g071(.A(G651), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(KEYINPUT6), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n499), .A2(G50), .A3(G543), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT69), .ZN(new_n501));
  XNOR2_X1  g076(.A(new_n500), .B(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT70), .B1(new_n503), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT5), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n503), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n499), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G88), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n504), .A2(new_n507), .B1(new_n503), .B2(G543), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  OAI211_X1 g090(.A(new_n502), .B(new_n513), .C1(new_n497), .C2(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  NAND3_X1  g092(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n518));
  OAI21_X1  g093(.A(KEYINPUT71), .B1(new_n496), .B2(new_n498), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n497), .A2(KEYINPUT6), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n495), .A2(G651), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT71), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n519), .A2(G543), .A3(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G51), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT72), .B(KEYINPUT7), .ZN(new_n527));
  AND3_X1   g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n527), .B(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n514), .A2(G89), .A3(new_n499), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n531), .A2(KEYINPUT73), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(KEYINPUT73), .ZN(new_n533));
  OAI211_X1 g108(.A(new_n518), .B(new_n526), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(G168));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n514), .A2(new_n499), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n536), .A2(new_n524), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n497), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT74), .ZN(new_n542));
  OR3_X1    g117(.A1(new_n539), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n539), .B2(new_n541), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(G171));
  INV_X1    g120(.A(G43), .ZN(new_n546));
  INV_X1    g121(.A(G81), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n546), .A2(new_n524), .B1(new_n537), .B2(new_n547), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT76), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n514), .A2(G56), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT75), .ZN(new_n551));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  AND3_X1   g127(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n551), .B1(new_n550), .B2(new_n552), .ZN(new_n554));
  NOR3_X1   g129(.A1(new_n553), .A2(new_n554), .A3(new_n497), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n549), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT77), .ZN(G153));
  AND3_X1   g133(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G36), .ZN(new_n560));
  XOR2_X1   g135(.A(new_n560), .B(KEYINPUT78), .Z(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n559), .A2(new_n563), .ZN(G188));
  AND3_X1   g139(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n522), .B1(new_n520), .B2(new_n521), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n567), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n519), .A2(G53), .A3(G543), .A4(new_n523), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  XOR2_X1   g147(.A(KEYINPUT79), .B(G65), .Z(new_n573));
  AOI22_X1  g148(.A1(new_n514), .A2(new_n573), .B1(G78), .B2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G91), .ZN(new_n575));
  OAI22_X1  g150(.A1(new_n574), .A2(new_n497), .B1(new_n575), .B2(new_n537), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(G299));
  INV_X1    g153(.A(G171), .ZN(G301));
  INV_X1    g154(.A(KEYINPUT80), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n534), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n531), .B(KEYINPUT73), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n582), .A2(KEYINPUT80), .A3(new_n518), .A4(new_n526), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(G286));
  NAND2_X1  g159(.A1(new_n525), .A2(G49), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n512), .A2(G87), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n588), .B(KEYINPUT81), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G288));
  AOI22_X1  g165(.A1(new_n514), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(new_n497), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n514), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n593), .A2(new_n511), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G305));
  INV_X1    g171(.A(G47), .ZN(new_n597));
  INV_X1    g172(.A(G85), .ZN(new_n598));
  OAI22_X1  g173(.A1(new_n597), .A2(new_n524), .B1(new_n537), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(new_n497), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(new_n512), .A2(G92), .ZN(new_n604));
  OR2_X1    g179(.A1(new_n604), .A2(KEYINPUT10), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n514), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n606), .A2(new_n497), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n525), .A2(G54), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n604), .A2(KEYINPUT10), .ZN(new_n609));
  NAND4_X1  g184(.A1(new_n605), .A2(new_n607), .A3(new_n608), .A4(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G171), .B2(new_n611), .ZN(G284));
  OAI21_X1  g188(.A(new_n612), .B1(G171), .B2(new_n611), .ZN(G321));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT82), .Z(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n577), .ZN(G297));
  OAI21_X1  g192(.A(new_n616), .B1(G868), .B2(new_n577), .ZN(G280));
  INV_X1    g193(.A(new_n610), .ZN(new_n619));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G860), .ZN(G148));
  NOR2_X1   g196(.A1(new_n610), .A2(G559), .ZN(new_n622));
  OR3_X1    g197(.A1(new_n622), .A2(KEYINPUT83), .A3(new_n611), .ZN(new_n623));
  OAI21_X1  g198(.A(KEYINPUT83), .B1(new_n622), .B2(new_n611), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n623), .B(new_n624), .C1(G868), .C2(new_n556), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g201(.A1(new_n480), .A2(G123), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n475), .A2(G135), .ZN(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n462), .A2(G111), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n627), .B(new_n628), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(G2096), .Z(new_n632));
  NAND3_X1  g207(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT12), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT13), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2100), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n632), .A2(new_n636), .ZN(G156));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT15), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n642), .A2(G2435), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(G2435), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(KEYINPUT14), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT84), .B(KEYINPUT16), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n647), .A2(new_n650), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n639), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n655), .A2(new_n651), .A3(new_n638), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n654), .A2(new_n656), .A3(G14), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(KEYINPUT85), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT85), .ZN(new_n659));
  NAND4_X1  g234(.A1(new_n654), .A2(new_n656), .A3(new_n659), .A4(G14), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT86), .ZN(G401));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  XNOR2_X1  g238(.A(G2072), .B(G2078), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2067), .B(G2678), .Z(new_n666));
  AOI21_X1  g241(.A(new_n663), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n664), .B(KEYINPUT17), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n667), .B1(new_n669), .B2(new_n666), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT87), .Z(new_n671));
  INV_X1    g246(.A(new_n666), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n672), .A2(new_n664), .A3(new_n663), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT18), .Z(new_n674));
  NAND3_X1  g249(.A1(new_n669), .A2(new_n663), .A3(new_n666), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n671), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT88), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2096), .B(G2100), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G227));
  XNOR2_X1  g254(.A(G1956), .B(G2474), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT89), .ZN(new_n681));
  XOR2_X1   g256(.A(G1961), .B(G1966), .Z(new_n682));
  AND2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G1971), .B(G1976), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT19), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT20), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n681), .A2(new_n682), .ZN(new_n688));
  AOI22_X1  g263(.A1(new_n686), .A2(new_n687), .B1(new_n685), .B2(new_n688), .ZN(new_n689));
  OR3_X1    g264(.A1(new_n683), .A2(new_n688), .A3(new_n685), .ZN(new_n690));
  OAI211_X1 g265(.A(new_n689), .B(new_n690), .C1(new_n687), .C2(new_n686), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1991), .B(G1996), .ZN(new_n694));
  INV_X1    g269(.A(G1981), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G1986), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n693), .B(new_n697), .ZN(G229));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G22), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G166), .B2(new_n699), .ZN(new_n701));
  INV_X1    g276(.A(G1971), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n699), .A2(G6), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(new_n595), .B2(new_n699), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT32), .B(G1981), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT90), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n705), .B(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n699), .A2(G23), .ZN(new_n709));
  INV_X1    g284(.A(new_n588), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(new_n699), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT33), .B(G1976), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT91), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n711), .B(new_n713), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n703), .A2(new_n708), .A3(new_n714), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n715), .A2(KEYINPUT34), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n480), .A2(G119), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n475), .A2(G131), .ZN(new_n718));
  OAI21_X1  g293(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n462), .A2(G107), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n717), .B(new_n718), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  MUX2_X1   g296(.A(G25), .B(new_n721), .S(G29), .Z(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT35), .B(G1991), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n722), .B(new_n723), .Z(new_n724));
  NAND2_X1  g299(.A1(new_n715), .A2(KEYINPUT34), .ZN(new_n725));
  NAND4_X1  g300(.A1(new_n716), .A2(KEYINPUT92), .A3(new_n724), .A4(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT36), .ZN(new_n727));
  NOR2_X1   g302(.A1(G16), .A2(G24), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n602), .B2(G16), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G1986), .ZN(new_n730));
  OR3_X1    g305(.A1(new_n726), .A2(new_n727), .A3(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G29), .ZN(new_n732));
  AND2_X1   g307(.A1(new_n732), .A2(G26), .ZN(new_n733));
  OR2_X1    g308(.A1(G104), .A2(G2105), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n734), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT93), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n480), .A2(G128), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n475), .A2(G140), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT94), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n733), .B1(new_n740), .B2(G29), .ZN(new_n741));
  MUX2_X1   g316(.A(new_n733), .B(new_n741), .S(KEYINPUT28), .Z(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G2067), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n699), .A2(KEYINPUT23), .A3(G20), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT23), .ZN(new_n745));
  INV_X1    g320(.A(G20), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n745), .B1(new_n746), .B2(G16), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n744), .B(new_n747), .C1(new_n577), .C2(new_n699), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G1956), .ZN(new_n749));
  NOR2_X1   g324(.A1(G29), .A2(G35), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G162), .B2(G29), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT29), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n749), .B1(new_n752), .B2(G2090), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT24), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n754), .A2(G34), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(G34), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n755), .A2(new_n756), .A3(new_n732), .ZN(new_n757));
  INV_X1    g332(.A(G160), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n757), .B1(new_n758), .B2(new_n732), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(G2084), .Z(new_n760));
  NAND2_X1  g335(.A1(new_n475), .A2(G141), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n480), .A2(G129), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n763));
  NAND3_X1  g338(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT26), .Z(new_n765));
  NAND4_X1  g340(.A1(new_n761), .A2(new_n762), .A3(new_n763), .A4(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(G29), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G29), .B2(G32), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT27), .B(G1996), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n760), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n699), .A2(G4), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n619), .B2(new_n699), .ZN(new_n773));
  INV_X1    g348(.A(G1348), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n743), .A2(new_n753), .A3(new_n771), .A4(new_n775), .ZN(new_n776));
  OR2_X1    g351(.A1(G29), .A2(G33), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT25), .Z(new_n779));
  NAND2_X1  g354(.A1(new_n475), .A2(G139), .ZN(new_n780));
  AND3_X1   g355(.A1(new_n779), .A2(new_n780), .A3(KEYINPUT95), .ZN(new_n781));
  AOI21_X1  g356(.A(KEYINPUT95), .B1(new_n779), .B2(new_n780), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n491), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n783));
  OAI22_X1  g358(.A1(new_n781), .A2(new_n782), .B1(new_n462), .B2(new_n783), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT96), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n777), .B1(new_n785), .B2(new_n732), .ZN(new_n786));
  INV_X1    g361(.A(G2072), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n752), .B2(G2090), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n699), .A2(G19), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n556), .B2(new_n699), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(G1341), .Z(new_n792));
  NOR2_X1   g367(.A1(G5), .A2(G16), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G171), .B2(G16), .ZN(new_n794));
  INV_X1    g369(.A(G1961), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n792), .B(new_n796), .C1(new_n787), .C2(new_n786), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n699), .A2(G21), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G168), .B2(new_n699), .ZN(new_n799));
  INV_X1    g374(.A(G1966), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(G164), .A2(G29), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G27), .B2(G29), .ZN(new_n803));
  INV_X1    g378(.A(G2078), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT97), .B(KEYINPUT30), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G28), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n803), .A2(new_n804), .B1(new_n732), .B2(new_n806), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n801), .B(new_n807), .C1(new_n804), .C2(new_n803), .ZN(new_n808));
  NOR4_X1   g383(.A1(new_n776), .A2(new_n789), .A3(new_n797), .A4(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT31), .B(G11), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n727), .B1(new_n726), .B2(new_n730), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n731), .A2(new_n809), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n769), .A2(new_n770), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n631), .A2(new_n732), .ZN(new_n815));
  NOR3_X1   g390(.A1(new_n812), .A2(new_n814), .A3(new_n815), .ZN(G311));
  INV_X1    g391(.A(G311), .ZN(G150));
  INV_X1    g392(.A(G55), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT98), .B(G93), .ZN(new_n819));
  OAI22_X1  g394(.A1(new_n818), .A2(new_n524), .B1(new_n537), .B2(new_n819), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n821), .A2(new_n497), .ZN(new_n822));
  OAI21_X1  g397(.A(G860), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT37), .Z(new_n824));
  NOR2_X1   g399(.A1(new_n610), .A2(new_n620), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT39), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n825), .B(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT76), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n548), .B(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n555), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n830), .B(new_n831), .C1(new_n822), .C2(new_n820), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n820), .A2(new_n822), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(new_n549), .B2(new_n555), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n828), .B(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n824), .B1(new_n837), .B2(G860), .ZN(G145));
  NAND2_X1  g413(.A1(new_n490), .A2(new_n493), .ZN(new_n839));
  INV_X1    g414(.A(new_n488), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n766), .B(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n740), .B(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n785), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n475), .A2(G142), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT100), .Z(new_n846));
  NAND2_X1  g421(.A1(new_n480), .A2(G130), .ZN(new_n847));
  OAI21_X1  g422(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n462), .A2(G118), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n846), .B(new_n847), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n721), .B(new_n634), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT101), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n844), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(new_n844), .B2(new_n852), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n631), .B(new_n758), .ZN(new_n856));
  XNOR2_X1  g431(.A(G162), .B(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(G37), .ZN(new_n859));
  INV_X1    g434(.A(new_n857), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n844), .A2(new_n853), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n860), .B1(new_n861), .B2(new_n854), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n858), .A2(new_n859), .A3(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g439(.A(new_n611), .B1(new_n820), .B2(new_n822), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n835), .B(new_n622), .Z(new_n866));
  AND2_X1   g441(.A1(new_n610), .A2(G299), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n610), .A2(G299), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(KEYINPUT41), .B1(new_n867), .B2(new_n868), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n619), .A2(new_n577), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT41), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n610), .A2(G299), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n871), .A2(new_n875), .A3(KEYINPUT102), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT102), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n869), .A2(new_n877), .A3(new_n873), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n870), .B1(new_n866), .B2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n595), .B(new_n588), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n881), .A2(G303), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(G303), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n602), .B(KEYINPUT103), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n882), .A2(new_n885), .A3(new_n883), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT42), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n880), .B(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n865), .B1(new_n891), .B2(new_n611), .ZN(G295));
  OAI21_X1  g467(.A(new_n865), .B1(new_n891), .B2(new_n611), .ZN(G331));
  NAND2_X1  g468(.A1(G301), .A2(new_n534), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n581), .A2(G171), .A3(new_n583), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(new_n836), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n835), .A2(new_n894), .A3(new_n895), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(new_n869), .A3(new_n898), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n835), .A2(new_n894), .A3(new_n895), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n835), .B1(new_n895), .B2(new_n894), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n899), .B1(new_n902), .B2(new_n879), .ZN(new_n903));
  INV_X1    g478(.A(new_n889), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI211_X1 g480(.A(new_n889), .B(new_n899), .C1(new_n902), .C2(new_n879), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n905), .A2(new_n859), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT43), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT104), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n871), .A2(new_n875), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n869), .A2(KEYINPUT104), .A3(new_n873), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n910), .B(new_n911), .C1(new_n900), .C2(new_n901), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n889), .B1(new_n912), .B2(new_n899), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(G37), .B1(new_n913), .B2(new_n914), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(new_n916), .A3(new_n906), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n908), .B1(new_n917), .B2(KEYINPUT43), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n907), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n912), .A2(new_n899), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n924), .A2(new_n914), .A3(new_n904), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n859), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n906), .B1(new_n913), .B2(new_n914), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n923), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n915), .A2(new_n916), .A3(KEYINPUT106), .A4(new_n906), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n922), .B1(new_n930), .B2(KEYINPUT43), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n920), .B1(new_n931), .B2(new_n919), .ZN(G397));
  NAND2_X1  g507(.A1(new_n595), .A2(new_n695), .ZN(new_n933));
  OAI21_X1  g508(.A(G1981), .B1(new_n592), .B2(new_n594), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT110), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n933), .B(new_n934), .C1(new_n935), .C2(KEYINPUT49), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(KEYINPUT49), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(G40), .ZN(new_n939));
  NOR3_X1   g514(.A1(new_n469), .A2(new_n472), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(G1384), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(new_n841), .A3(new_n941), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n933), .A2(new_n935), .A3(KEYINPUT49), .A4(new_n934), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n938), .A2(G8), .A3(new_n942), .A4(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(G8), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n945), .B1(G1976), .B2(new_n710), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT52), .ZN(new_n947));
  OR2_X1    g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n946), .B(new_n947), .C1(new_n589), .C2(G1976), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n944), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(G303), .A2(G8), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n951), .B(KEYINPUT55), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT45), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n953), .B1(G164), .B2(G1384), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n841), .A2(KEYINPUT45), .A3(new_n941), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n954), .A2(new_n955), .A3(new_n940), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n702), .ZN(new_n957));
  OAI21_X1  g532(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT50), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n841), .A2(new_n959), .A3(new_n941), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n958), .A2(new_n960), .A3(new_n940), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n957), .B1(G2090), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(G8), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n952), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n952), .A2(new_n963), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n950), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  NOR2_X1   g541(.A1(KEYINPUT112), .A2(KEYINPUT63), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n956), .A2(new_n800), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n968), .B1(G2084), .B2(new_n961), .ZN(new_n969));
  AND4_X1   g544(.A1(G8), .A2(new_n969), .A3(new_n581), .A4(new_n583), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n966), .A2(new_n967), .A3(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n964), .A2(new_n965), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n944), .A2(new_n948), .A3(new_n949), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(new_n973), .A3(new_n970), .ZN(new_n974));
  XOR2_X1   g549(.A(KEYINPUT112), .B(KEYINPUT63), .Z(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G1976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n944), .A2(new_n977), .A3(new_n589), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n933), .ZN(new_n979));
  XOR2_X1   g554(.A(new_n945), .B(KEYINPUT111), .Z(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n973), .A2(new_n965), .ZN(new_n982));
  AND4_X1   g557(.A1(new_n971), .A2(new_n976), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G1956), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n961), .A2(new_n984), .ZN(new_n985));
  XNOR2_X1  g560(.A(KEYINPUT56), .B(G2072), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n954), .A2(new_n955), .A3(new_n940), .A4(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n569), .B(KEYINPUT9), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n514), .A2(new_n573), .ZN(new_n990));
  NAND2_X1  g565(.A1(G78), .A2(G543), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AOI22_X1  g567(.A1(new_n992), .A2(G651), .B1(new_n512), .B2(G91), .ZN(new_n993));
  OR2_X1    g568(.A1(KEYINPUT113), .A2(KEYINPUT57), .ZN(new_n994));
  NAND2_X1  g569(.A1(KEYINPUT113), .A2(KEYINPUT57), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n989), .A2(new_n993), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  OAI211_X1 g571(.A(KEYINPUT113), .B(KEYINPUT57), .C1(new_n572), .C2(new_n576), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n988), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G2067), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n467), .A2(new_n468), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(G2105), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n470), .A2(new_n471), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1002), .A2(new_n1003), .A3(G40), .ZN(new_n1004));
  NOR3_X1   g579(.A1(new_n1004), .A2(G164), .A3(G1384), .ZN(new_n1005));
  AOI22_X1  g580(.A1(new_n961), .A2(new_n774), .B1(new_n1000), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n999), .B1(new_n610), .B2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n985), .A2(new_n987), .A3(new_n996), .A4(new_n997), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT114), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n996), .A2(new_n997), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1010), .A2(new_n1011), .A3(new_n985), .A4(new_n987), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1007), .A2(new_n1009), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g589(.A(KEYINPUT58), .B(G1341), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT115), .B1(new_n1005), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G1996), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n954), .A2(new_n955), .A3(new_n1017), .A4(new_n940), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT115), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1015), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n942), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1016), .A2(new_n1018), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(new_n556), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT116), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT117), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1022), .A2(new_n1026), .A3(new_n556), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1024), .A2(new_n1025), .A3(KEYINPUT59), .A4(new_n1027), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n1022), .A2(new_n1026), .A3(new_n556), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1026), .B1(new_n1022), .B2(new_n556), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT59), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1025), .B1(new_n1023), .B2(KEYINPUT59), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  OAI211_X1 g609(.A(KEYINPUT118), .B(new_n1028), .C1(new_n1032), .C2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1024), .A2(KEYINPUT59), .A3(new_n1027), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n1033), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT118), .B1(new_n1038), .B2(new_n1028), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n999), .A2(KEYINPUT61), .A3(new_n1008), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n1009), .A2(new_n999), .A3(new_n1012), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1041), .B1(new_n1042), .B2(KEYINPUT61), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1006), .A2(KEYINPUT60), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT60), .ZN(new_n1045));
  AOI221_X4 g620(.A(new_n1045), .B1(new_n1005), .B2(new_n1000), .C1(new_n961), .C2(new_n774), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n619), .B1(new_n1046), .B2(KEYINPUT119), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1006), .A2(KEYINPUT60), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT119), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1048), .A2(new_n1049), .A3(new_n610), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1047), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1046), .A2(KEYINPUT119), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1044), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1043), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1014), .B1(new_n1040), .B2(new_n1054), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n954), .A2(new_n955), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1056), .A2(new_n804), .A3(new_n940), .ZN(new_n1057));
  XOR2_X1   g632(.A(KEYINPUT121), .B(KEYINPUT53), .Z(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n961), .A2(new_n795), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1060), .B1(new_n1057), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT120), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1059), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  XOR2_X1   g641(.A(G171), .B(KEYINPUT54), .Z(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(G8), .B1(new_n969), .B2(new_n534), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT51), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1070), .B1(new_n969), .B2(new_n534), .ZN(new_n1071));
  OR2_X1    g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1069), .A2(KEYINPUT51), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT122), .ZN(new_n1075));
  OAI21_X1  g650(.A(KEYINPUT53), .B1(new_n1004), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1076), .B1(new_n1075), .B2(new_n1004), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1077), .A2(new_n804), .A3(new_n1056), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1079));
  OR3_X1    g654(.A1(new_n1067), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n966), .A2(new_n1068), .A3(new_n1074), .A4(new_n1080), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n983), .B(KEYINPUT123), .C1(new_n1055), .C2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT123), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1028), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1054), .A2(new_n1086), .A3(new_n1035), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1081), .B1(new_n1087), .B2(new_n1013), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n976), .A2(new_n971), .A3(new_n981), .A4(new_n982), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1083), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT124), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1074), .A2(KEYINPUT62), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT62), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1072), .A2(new_n1093), .A3(new_n1073), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1092), .A2(G171), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n966), .A2(new_n1066), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1091), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1096), .ZN(new_n1098));
  AOI21_X1  g673(.A(G301), .B1(new_n1074), .B2(KEYINPUT62), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1098), .A2(new_n1099), .A3(KEYINPUT124), .A4(new_n1094), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1082), .A2(new_n1090), .A3(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n740), .B(new_n1000), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1103), .B1(new_n1017), .B2(new_n767), .ZN(new_n1104));
  INV_X1    g679(.A(new_n954), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n940), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1106), .A2(G1996), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1108), .B(KEYINPUT108), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1104), .A2(new_n1107), .B1(new_n767), .B2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n721), .A2(new_n723), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n721), .A2(new_n723), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1107), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1114));
  OR2_X1    g689(.A1(G290), .A2(G1986), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(KEYINPUT107), .ZN(new_n1116));
  NAND2_X1  g691(.A1(G290), .A2(G1986), .ZN(new_n1117));
  XOR2_X1   g692(.A(new_n1116), .B(new_n1117), .Z(new_n1118));
  OAI21_X1  g693(.A(new_n1114), .B1(new_n1106), .B2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n1119), .B(KEYINPUT109), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1102), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1106), .B1(new_n1103), .B2(new_n767), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT125), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1122), .B1(new_n1123), .B2(KEYINPUT46), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1109), .B1(new_n1123), .B2(KEYINPUT46), .ZN(new_n1125));
  OR3_X1    g700(.A1(new_n1109), .A2(new_n1123), .A3(KEYINPUT46), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1127), .B(KEYINPUT47), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1115), .A2(new_n1106), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n1129), .B(KEYINPUT126), .ZN(new_n1130));
  XOR2_X1   g705(.A(new_n1130), .B(KEYINPUT48), .Z(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n1114), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n740), .A2(G2067), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1107), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1128), .A2(new_n1132), .A3(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1136), .B(KEYINPUT127), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1121), .A2(new_n1137), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g713(.A(G227), .B1(new_n658), .B2(new_n660), .ZN(new_n1140));
  AND2_X1   g714(.A1(new_n1140), .A2(new_n863), .ZN(new_n1141));
  INV_X1    g715(.A(G229), .ZN(new_n1142));
  NAND4_X1  g716(.A1(new_n1141), .A2(new_n460), .A3(new_n918), .A4(new_n1142), .ZN(G225));
  INV_X1    g717(.A(G225), .ZN(G308));
endmodule


