//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 1 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 0 0 0 1 0 0 1 1 0 0 0 1 1 1 0 1 0 0 0 1 1 1 1 0 0 0 1 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n819, new_n820, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G140), .ZN(new_n189));
  INV_X1    g003(.A(G227), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G953), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n189), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G143), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT1), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n199), .B1(G143), .B2(new_n194), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n198), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n204));
  AND3_X1   g018(.A1(new_n196), .A2(KEYINPUT64), .A3(G146), .ZN(new_n205));
  AOI21_X1  g019(.A(KEYINPUT64), .B1(new_n196), .B2(G146), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n195), .B(new_n204), .C1(new_n205), .C2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n210), .B1(new_n194), .B2(G143), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n196), .A2(KEYINPUT64), .A3(G146), .ZN(new_n212));
  AOI22_X1  g026(.A1(new_n211), .A2(new_n212), .B1(G143), .B2(new_n194), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(KEYINPUT65), .A3(new_n204), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n203), .B1(new_n209), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT10), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n218));
  INV_X1    g032(.A(G107), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n219), .A3(G104), .ZN(new_n220));
  INV_X1    g034(.A(G104), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G107), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G101), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT3), .B1(new_n221), .B2(G107), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n223), .A2(KEYINPUT78), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n225), .A2(new_n220), .A3(new_n224), .A4(new_n222), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT78), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n219), .A2(G104), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(new_n222), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G101), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT80), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n231), .A2(KEYINPUT80), .A3(G101), .ZN(new_n235));
  AOI22_X1  g049(.A1(new_n226), .A2(new_n229), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n225), .A2(new_n220), .A3(new_n222), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G101), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n227), .A2(new_n228), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n227), .A2(new_n228), .ZN(new_n240));
  OAI211_X1 g054(.A(KEYINPUT4), .B(new_n238), .C1(new_n239), .C2(new_n240), .ZN(new_n241));
  AND2_X1   g055(.A1(KEYINPUT0), .A2(G128), .ZN(new_n242));
  NOR2_X1   g056(.A1(KEYINPUT0), .A2(G128), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n213), .A2(new_n242), .B1(new_n244), .B2(new_n198), .ZN(new_n245));
  XOR2_X1   g059(.A(KEYINPUT79), .B(KEYINPUT4), .Z(new_n246));
  NAND3_X1  g060(.A1(new_n237), .A2(G101), .A3(new_n246), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n217), .A2(new_n236), .B1(new_n241), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT82), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n195), .B1(new_n205), .B2(new_n206), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT81), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n195), .A2(new_n252), .A3(KEYINPUT1), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G128), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n200), .A2(new_n252), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n251), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n207), .A2(new_n208), .ZN(new_n257));
  AOI21_X1  g071(.A(KEYINPUT65), .B1(new_n213), .B2(new_n204), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n236), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n250), .B1(new_n260), .B2(new_n216), .ZN(new_n261));
  AOI211_X1 g075(.A(KEYINPUT82), .B(KEYINPUT10), .C1(new_n259), .C2(new_n236), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n249), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT83), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT11), .ZN(new_n266));
  INV_X1    g080(.A(G134), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n266), .B1(new_n267), .B2(G137), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(G137), .ZN(new_n269));
  INV_X1    g083(.A(G137), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(KEYINPUT11), .A3(G134), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n268), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G131), .ZN(new_n273));
  INV_X1    g087(.A(G131), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n268), .A2(new_n271), .A3(new_n274), .A4(new_n269), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  OAI211_X1 g090(.A(KEYINPUT83), .B(new_n249), .C1(new_n261), .C2(new_n262), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n265), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n276), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n279), .B(new_n249), .C1(new_n261), .C2(new_n262), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n193), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n226), .A2(new_n229), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n234), .A2(new_n235), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n215), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n279), .B1(new_n285), .B2(new_n260), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n286), .A2(KEYINPUT12), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n286), .A2(KEYINPUT12), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n280), .A2(new_n193), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n187), .B(new_n188), .C1(new_n281), .C2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n187), .A2(new_n188), .ZN(new_n293));
  INV_X1    g107(.A(new_n290), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n280), .B1(new_n287), .B2(new_n288), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n278), .A2(new_n294), .B1(new_n192), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n293), .B1(new_n296), .B2(G469), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G125), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT73), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT73), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G125), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n245), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n304), .B1(new_n215), .B2(new_n303), .ZN(new_n305));
  INV_X1    g119(.A(G224), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n306), .A2(G953), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n307), .B(KEYINPUT86), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n305), .B(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT2), .ZN(new_n311));
  INV_X1    g125(.A(G113), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(new_n312), .A3(KEYINPUT66), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT66), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n314), .B1(KEYINPUT2), .B2(G113), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(KEYINPUT2), .A2(G113), .ZN(new_n317));
  XNOR2_X1  g131(.A(G116), .B(G119), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT67), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI22_X1  g135(.A1(new_n313), .A2(new_n315), .B1(KEYINPUT2), .B2(G113), .ZN(new_n322));
  AOI21_X1  g136(.A(KEYINPUT67), .B1(new_n322), .B2(new_n318), .ZN(new_n323));
  OAI22_X1  g137(.A1(new_n321), .A2(new_n323), .B1(new_n322), .B2(new_n318), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n324), .A2(new_n241), .A3(new_n247), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n319), .A2(new_n320), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n322), .A2(KEYINPUT67), .A3(new_n318), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G116), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n329), .A2(G119), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT5), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n312), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT84), .ZN(new_n333));
  INV_X1    g147(.A(G119), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G116), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n329), .A2(G119), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n335), .A2(new_n336), .A3(KEYINPUT5), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n332), .A2(new_n333), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n333), .B1(new_n332), .B2(new_n337), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n236), .A2(new_n328), .A3(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(G110), .B(G122), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n325), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  AND2_X1   g157(.A1(KEYINPUT85), .A2(KEYINPUT6), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n342), .B1(new_n325), .B2(new_n341), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n344), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n310), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n342), .B(KEYINPUT8), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n340), .A2(new_n328), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n284), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n332), .A2(new_n337), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n328), .A2(new_n355), .ZN(new_n356));
  AOI22_X1  g170(.A1(new_n354), .A2(KEYINPUT87), .B1(new_n356), .B2(new_n236), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n340), .A2(new_n328), .B1(new_n282), .B2(new_n283), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT87), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n352), .B1(new_n357), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(KEYINPUT7), .B1(new_n306), .B2(G953), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n304), .B(new_n362), .C1(new_n215), .C2(new_n303), .ZN(new_n363));
  INV_X1    g177(.A(new_n362), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n305), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n343), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n188), .B1(new_n361), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(G210), .B1(G237), .B2(G902), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NOR3_X1   g183(.A1(new_n350), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n346), .B1(new_n344), .B2(new_n343), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n346), .A2(new_n344), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n309), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AND3_X1   g187(.A1(new_n343), .A2(new_n363), .A3(new_n365), .ZN(new_n374));
  INV_X1    g188(.A(new_n360), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n236), .A2(new_n328), .A3(new_n355), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n376), .B1(new_n358), .B2(new_n359), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n351), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(G902), .B1(new_n374), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n368), .B1(new_n373), .B2(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n370), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(G214), .B1(G237), .B2(G902), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT9), .B(G234), .ZN(new_n385));
  OAI21_X1  g199(.A(G221), .B1(new_n385), .B2(G902), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n298), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G953), .ZN(new_n388));
  AND2_X1   g202(.A1(new_n388), .A2(G952), .ZN(new_n389));
  NAND2_X1  g203(.A1(G234), .A2(G237), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(G902), .A3(G953), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(KEYINPUT21), .B(G898), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n392), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  AND2_X1   g211(.A1(new_n387), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT91), .ZN(new_n399));
  XNOR2_X1  g213(.A(G113), .B(G122), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n400), .B(new_n221), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  OR2_X1    g216(.A1(new_n196), .A2(KEYINPUT88), .ZN(new_n403));
  INV_X1    g217(.A(G237), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(new_n388), .A3(G214), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT88), .B(G143), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n406), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(KEYINPUT18), .A2(G131), .ZN(new_n409));
  OR3_X1    g223(.A1(new_n408), .A2(KEYINPUT89), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT18), .ZN(new_n411));
  OAI22_X1  g225(.A1(new_n408), .A2(KEYINPUT89), .B1(new_n411), .B2(new_n274), .ZN(new_n412));
  XOR2_X1   g226(.A(G125), .B(G140), .Z(new_n413));
  NOR2_X1   g227(.A1(new_n413), .A2(G146), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G140), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n416), .B1(new_n300), .B2(new_n302), .ZN(new_n417));
  NOR2_X1   g231(.A1(G125), .A2(G140), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G146), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n410), .A2(new_n412), .B1(new_n415), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n408), .A2(G131), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT17), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n406), .B(new_n274), .C1(new_n405), .C2(new_n407), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT16), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n301), .A2(G125), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n299), .A2(KEYINPUT73), .ZN(new_n428));
  OAI21_X1  g242(.A(G140), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n418), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n426), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n303), .A2(new_n426), .A3(new_n416), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n194), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(KEYINPUT16), .B1(new_n417), .B2(new_n418), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(G146), .A3(new_n432), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n408), .A2(KEYINPUT17), .A3(G131), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n434), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n425), .B1(new_n438), .B2(KEYINPUT90), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT90), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n434), .A2(new_n440), .A3(new_n436), .A4(new_n437), .ZN(new_n441));
  AOI211_X1 g255(.A(new_n402), .B(new_n421), .C1(new_n439), .C2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n421), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n413), .A2(KEYINPUT19), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n444), .B1(KEYINPUT19), .B2(new_n419), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n194), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n422), .A2(new_n424), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n436), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n401), .B1(new_n443), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n399), .B1(new_n442), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(G475), .A2(G902), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n439), .A2(new_n441), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(new_n401), .A3(new_n443), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n443), .A2(new_n448), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n402), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n453), .A2(KEYINPUT91), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n450), .A2(new_n451), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(KEYINPUT20), .ZN(new_n458));
  NOR3_X1   g272(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n459), .B1(new_n442), .B2(new_n449), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G217), .ZN(new_n462));
  NOR3_X1   g276(.A1(new_n385), .A2(new_n462), .A3(G953), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT93), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n201), .A2(G143), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n196), .A2(G128), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT13), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n201), .A2(G143), .ZN(new_n470));
  OAI21_X1  g284(.A(KEYINPUT92), .B1(new_n470), .B2(KEYINPUT13), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT92), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n467), .A2(new_n472), .A3(new_n468), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n469), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(new_n267), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n467), .A2(new_n466), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n267), .ZN(new_n478));
  INV_X1    g292(.A(G122), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G116), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n329), .A2(G122), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(new_n481), .A3(new_n219), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n219), .B1(new_n480), .B2(new_n481), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n478), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n465), .B1(new_n475), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n484), .ZN(new_n487));
  AOI22_X1  g301(.A1(new_n487), .A2(new_n482), .B1(new_n477), .B2(new_n267), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n488), .B(KEYINPUT93), .C1(new_n267), .C2(new_n474), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n476), .A2(G134), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n483), .B1(new_n478), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT14), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n494), .B1(new_n329), .B2(G122), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT94), .ZN(new_n496));
  OR2_X1    g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n495), .A2(new_n496), .B1(G116), .B2(new_n479), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT95), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n494), .A2(new_n329), .A3(G122), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n497), .A2(new_n498), .A3(KEYINPUT95), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n493), .B1(new_n504), .B2(G107), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n464), .B1(new_n490), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n503), .A2(new_n502), .ZN(new_n507));
  AOI21_X1  g321(.A(KEYINPUT95), .B1(new_n497), .B2(new_n498), .ZN(new_n508));
  OAI21_X1  g322(.A(G107), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n492), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n486), .A2(new_n489), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n511), .A3(new_n463), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n506), .A2(KEYINPUT96), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT96), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n514), .B(new_n464), .C1(new_n490), .C2(new_n505), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n513), .A2(new_n188), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(G478), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n517), .A2(KEYINPUT15), .ZN(new_n518));
  XOR2_X1   g332(.A(new_n516), .B(new_n518), .Z(new_n519));
  INV_X1    g333(.A(G475), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n401), .B1(new_n452), .B2(new_n443), .ZN(new_n521));
  OR2_X1    g335(.A1(new_n521), .A2(new_n442), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n520), .B1(new_n522), .B2(new_n188), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n461), .A2(new_n519), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT23), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n527), .B1(new_n334), .B2(G128), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n334), .A2(G128), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n201), .A2(KEYINPUT23), .A3(G119), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(G110), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT72), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n534), .B1(new_n334), .B2(G128), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n201), .A2(KEYINPUT72), .A3(G119), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n535), .A2(new_n536), .A3(new_n529), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT24), .B(G110), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n414), .B1(new_n533), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n436), .ZN(new_n541));
  XNOR2_X1  g355(.A(KEYINPUT22), .B(G137), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n388), .A2(G221), .A3(G234), .ZN(new_n543));
  XOR2_X1   g357(.A(new_n542), .B(new_n543), .Z(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n434), .A2(new_n436), .ZN(new_n546));
  OAI22_X1  g360(.A1(new_n531), .A2(new_n532), .B1(new_n538), .B2(new_n537), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT74), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT74), .ZN(new_n550));
  AOI211_X1 g364(.A(new_n550), .B(new_n547), .C1(new_n434), .C2(new_n436), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n541), .B(new_n545), .C1(new_n549), .C2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n541), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n435), .A2(G146), .A3(new_n432), .ZN(new_n554));
  AOI21_X1  g368(.A(G146), .B1(new_n435), .B2(new_n432), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n548), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n550), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n546), .A2(KEYINPUT74), .A3(new_n548), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n553), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n544), .B(KEYINPUT75), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n552), .B(new_n188), .C1(new_n559), .C2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT25), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT76), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n557), .A2(new_n558), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n561), .B1(new_n566), .B2(new_n541), .ZN(new_n567));
  AOI211_X1 g381(.A(new_n553), .B(new_n544), .C1(new_n557), .C2(new_n558), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n569), .A2(KEYINPUT77), .A3(KEYINPUT25), .A4(new_n188), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT77), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n571), .B1(new_n562), .B2(new_n563), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT76), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n562), .A2(new_n573), .A3(new_n563), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n565), .A2(new_n570), .A3(new_n572), .A4(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n462), .B1(G234), .B2(new_n188), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n576), .A2(G902), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n569), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT31), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n322), .A2(new_n318), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n582), .B1(new_n326), .B2(new_n327), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n245), .A2(new_n276), .ZN(new_n584));
  INV_X1    g398(.A(new_n269), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n267), .A2(G137), .ZN(new_n586));
  OAI21_X1  g400(.A(G131), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n275), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n583), .B(new_n584), .C1(new_n215), .C2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n584), .B1(new_n215), .B2(new_n588), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT30), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT30), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n584), .B(new_n593), .C1(new_n215), .C2(new_n588), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n590), .B1(new_n595), .B2(new_n324), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n404), .A2(new_n388), .A3(G210), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(KEYINPUT27), .ZN(new_n598));
  XNOR2_X1  g412(.A(KEYINPUT26), .B(G101), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n598), .B(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n581), .B1(new_n596), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n583), .B1(new_n592), .B2(new_n594), .ZN(new_n602));
  INV_X1    g416(.A(new_n600), .ZN(new_n603));
  NOR4_X1   g417(.A1(new_n602), .A2(KEYINPUT31), .A3(new_n590), .A4(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT28), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n589), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n202), .B1(new_n257), .B2(new_n258), .ZN(new_n607));
  INV_X1    g421(.A(new_n588), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n609), .A2(KEYINPUT28), .A3(new_n583), .A4(new_n584), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n591), .A2(new_n324), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n606), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n603), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n601), .A2(new_n604), .A3(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(G472), .A2(G902), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(KEYINPUT68), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT32), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n593), .B1(new_n609), .B2(new_n584), .ZN(new_n620));
  INV_X1    g434(.A(new_n594), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n324), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n622), .A2(new_n589), .A3(new_n600), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT31), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n596), .A2(new_n581), .A3(new_n600), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n624), .A2(new_n613), .A3(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT68), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n626), .A2(new_n627), .A3(new_n616), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n618), .A2(new_n619), .A3(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n626), .A2(KEYINPUT32), .A3(new_n616), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT69), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n611), .A2(new_n632), .A3(new_n589), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n591), .A2(KEYINPUT69), .A3(new_n324), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n633), .A2(KEYINPUT28), .A3(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT29), .ZN(new_n636));
  AOI211_X1 g450(.A(new_n636), .B(new_n603), .C1(new_n589), .C2(new_n605), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n188), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT70), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n638), .A2(KEYINPUT70), .A3(new_n188), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n622), .A2(new_n589), .A3(new_n603), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n612), .A2(new_n600), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n636), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n641), .A2(new_n642), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(G472), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(KEYINPUT71), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT71), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n647), .A2(new_n650), .A3(G472), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n580), .B1(new_n631), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n398), .A2(new_n526), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G101), .ZN(G3));
  NAND2_X1  g469(.A1(new_n298), .A2(new_n386), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n626), .A2(new_n188), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(G472), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n658), .A2(new_n618), .A3(new_n628), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n656), .A2(new_n580), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT97), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT33), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n513), .A2(new_n662), .A3(new_n515), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n506), .A2(KEYINPUT33), .A3(new_n512), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n517), .A2(G902), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT99), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n516), .A2(new_n517), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n667), .B1(new_n666), .B2(new_n668), .ZN(new_n670));
  INV_X1    g484(.A(new_n460), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n671), .B1(new_n457), .B2(KEYINPUT20), .ZN(new_n672));
  OAI22_X1  g486(.A1(new_n669), .A2(new_n670), .B1(new_n672), .B2(new_n523), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n383), .B1(new_n380), .B2(KEYINPUT98), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n369), .B1(new_n350), .B2(new_n367), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT98), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n373), .A2(new_n379), .A3(new_n368), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n674), .A2(new_n678), .A3(new_n397), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n661), .A2(new_n673), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G104), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G6));
  NAND2_X1  g498(.A1(new_n458), .A2(KEYINPUT101), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT101), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n457), .A2(new_n686), .A3(KEYINPUT20), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n450), .A2(new_n456), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n459), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n685), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n516), .B(new_n518), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n690), .A2(new_n524), .A3(new_n691), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n661), .A2(new_n680), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(KEYINPUT35), .B(G107), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G9));
  NOR2_X1   g509(.A1(new_n560), .A2(KEYINPUT36), .ZN(new_n696));
  XOR2_X1   g510(.A(new_n559), .B(new_n696), .Z(new_n697));
  AND2_X1   g511(.A1(new_n697), .A2(new_n578), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n698), .B1(new_n575), .B2(new_n576), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n525), .A2(new_n699), .A3(new_n396), .ZN(new_n700));
  INV_X1    g514(.A(new_n659), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n700), .A2(new_n387), .A3(new_n701), .ZN(new_n702));
  XOR2_X1   g516(.A(KEYINPUT37), .B(G110), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G12));
  INV_X1    g518(.A(new_n386), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n705), .B1(new_n292), .B2(new_n297), .ZN(new_n706));
  INV_X1    g520(.A(new_n698), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n577), .A2(new_n707), .ZN(new_n708));
  AND2_X1   g522(.A1(new_n674), .A2(new_n678), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n706), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n388), .A2(G900), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n711), .A2(G902), .A3(new_n390), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n712), .A2(KEYINPUT102), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(KEYINPUT102), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n713), .A2(new_n391), .A3(new_n714), .ZN(new_n715));
  AND4_X1   g529(.A1(new_n524), .A2(new_n690), .A3(new_n691), .A4(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(G472), .ZN(new_n717));
  AOI22_X1  g531(.A1(new_n639), .A2(new_n640), .B1(new_n645), .B2(new_n636), .ZN(new_n718));
  AOI211_X1 g532(.A(KEYINPUT71), .B(new_n717), .C1(new_n718), .C2(new_n642), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n650), .B1(new_n647), .B2(G472), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n629), .B(new_n630), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n710), .A2(new_n716), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G128), .ZN(G30));
  XOR2_X1   g537(.A(new_n715), .B(KEYINPUT39), .Z(new_n724));
  NOR2_X1   g538(.A1(new_n656), .A2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT40), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT104), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n708), .A2(new_n383), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n691), .B1(new_n672), .B2(new_n523), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n381), .A2(KEYINPUT38), .ZN(new_n732));
  OR2_X1    g546(.A1(new_n381), .A2(KEYINPUT38), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n729), .A2(new_n731), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n633), .A2(new_n634), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n623), .B1(new_n735), .B2(new_n600), .ZN(new_n736));
  AOI21_X1  g550(.A(G902), .B1(new_n736), .B2(KEYINPUT103), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n737), .B1(KEYINPUT103), .B2(new_n736), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(G472), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n629), .A2(new_n739), .A3(new_n630), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n728), .B1(new_n734), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n733), .A2(new_n732), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n743), .A2(new_n383), .A3(new_n708), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n744), .A2(KEYINPUT104), .A3(new_n740), .A4(new_n731), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n727), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  XOR2_X1   g560(.A(KEYINPUT105), .B(G143), .Z(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G45));
  INV_X1    g562(.A(new_n715), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n673), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n710), .A2(new_n721), .A3(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G146), .ZN(G48));
  NOR2_X1   g566(.A1(new_n680), .A2(new_n673), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n607), .A2(new_n236), .A3(KEYINPUT10), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n241), .A2(new_n248), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n195), .A2(KEYINPUT1), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT81), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(G128), .A3(new_n253), .ZN(new_n759));
  AOI22_X1  g573(.A1(new_n209), .A2(new_n214), .B1(new_n759), .B2(new_n251), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n216), .B1(new_n284), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(KEYINPUT82), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n260), .A2(new_n250), .A3(new_n216), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n756), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n276), .B1(new_n764), .B2(KEYINPUT83), .ZN(new_n765));
  INV_X1    g579(.A(new_n277), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n280), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n291), .B1(new_n767), .B2(new_n192), .ZN(new_n768));
  OAI21_X1  g582(.A(G469), .B1(new_n768), .B2(G902), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n769), .A2(new_n386), .A3(new_n292), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n653), .A2(new_n753), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(KEYINPUT41), .B(G113), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n771), .B(new_n772), .ZN(G15));
  NOR2_X1   g587(.A1(new_n692), .A2(new_n680), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n653), .A2(new_n774), .A3(new_n770), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G116), .ZN(G18));
  NAND2_X1  g590(.A1(new_n769), .A2(new_n292), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n674), .A2(new_n678), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n777), .A2(new_n705), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(new_n700), .A3(new_n721), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G119), .ZN(G21));
  AND2_X1   g595(.A1(new_n635), .A2(new_n606), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n624), .B(new_n625), .C1(new_n782), .C2(new_n600), .ZN(new_n783));
  AOI22_X1  g597(.A1(new_n657), .A2(G472), .B1(new_n783), .B2(new_n616), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n580), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n730), .A2(new_n778), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n786), .A2(new_n397), .A3(new_n770), .A4(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(KEYINPUT106), .B(G122), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n788), .B(new_n789), .ZN(G24));
  NAND4_X1  g604(.A1(new_n709), .A2(new_n386), .A3(new_n292), .A4(new_n769), .ZN(new_n791));
  INV_X1    g605(.A(new_n576), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n570), .A2(new_n572), .ZN(new_n793));
  INV_X1    g607(.A(new_n574), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n573), .B1(new_n562), .B2(new_n563), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n792), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n784), .B1(new_n797), .B2(new_n698), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n666), .A2(new_n668), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(KEYINPUT99), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n461), .A2(new_n524), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n803), .A3(new_n715), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n791), .A2(new_n798), .A3(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(new_n299), .ZN(G27));
  INV_X1    g620(.A(new_n580), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n675), .A2(new_n382), .A3(new_n677), .ZN(new_n808));
  AOI211_X1 g622(.A(new_n705), .B(new_n808), .C1(new_n292), .C2(new_n297), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n721), .A2(new_n807), .A3(new_n750), .A4(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT42), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n619), .B1(new_n615), .B2(new_n617), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n652), .A2(new_n630), .A3(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n804), .A2(new_n811), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n814), .A2(new_n815), .A3(new_n807), .A4(new_n809), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G131), .ZN(G33));
  NAND2_X1  g632(.A1(new_n716), .A2(KEYINPUT107), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT107), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n820), .B1(new_n692), .B2(new_n749), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n819), .A2(new_n653), .A3(new_n809), .A4(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(G134), .ZN(G36));
  INV_X1    g637(.A(new_n293), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT45), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n278), .A2(new_n294), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n295), .A2(new_n192), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n296), .A2(KEYINPUT45), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(G469), .A3(new_n829), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n830), .A2(KEYINPUT108), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n830), .A2(KEYINPUT108), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n824), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT46), .ZN(new_n834));
  OAI21_X1  g648(.A(KEYINPUT109), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n833), .A2(new_n834), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n830), .B(KEYINPUT108), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT109), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n837), .A2(new_n838), .A3(KEYINPUT46), .A4(new_n824), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n835), .A2(new_n836), .A3(new_n292), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(new_n386), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n724), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT110), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n672), .A2(new_n523), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n802), .A2(new_n844), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n845), .A2(KEYINPUT43), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(KEYINPUT43), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n701), .A2(new_n699), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT44), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n843), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n846), .A2(KEYINPUT44), .A3(new_n847), .A4(new_n848), .ZN(new_n852));
  INV_X1    g666(.A(new_n808), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n849), .A2(new_n843), .A3(new_n850), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n842), .A2(new_n858), .ZN(new_n859));
  XOR2_X1   g673(.A(KEYINPUT111), .B(G137), .Z(new_n860));
  XNOR2_X1  g674(.A(new_n859), .B(new_n860), .ZN(G39));
  NOR4_X1   g675(.A1(new_n721), .A2(new_n804), .A3(new_n807), .A4(new_n808), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n840), .A2(KEYINPUT47), .A3(new_n386), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT47), .B1(new_n840), .B2(new_n386), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(G140), .ZN(G42));
  NAND4_X1  g680(.A1(new_n846), .A2(new_n392), .A3(new_n786), .A4(new_n847), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n743), .A2(new_n770), .A3(new_n383), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(KEYINPUT50), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n777), .A2(new_n705), .A3(new_n808), .ZN(new_n871));
  AND4_X1   g685(.A1(new_n392), .A2(new_n871), .A3(new_n807), .A4(new_n741), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n872), .A2(new_n844), .A3(new_n801), .A4(new_n800), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n846), .A2(new_n871), .A3(new_n392), .A4(new_n847), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n874), .A2(KEYINPUT116), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(KEYINPUT116), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n870), .B(new_n873), .C1(new_n798), .C2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n777), .A2(new_n386), .ZN(new_n879));
  OR3_X1    g693(.A1(new_n863), .A2(new_n864), .A3(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n867), .A2(new_n808), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n878), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n882), .A2(KEYINPUT51), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(KEYINPUT51), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n814), .A2(new_n807), .ZN(new_n885));
  AOI211_X1 g699(.A(new_n885), .B(new_n877), .C1(KEYINPUT118), .C2(KEYINPUT48), .ZN(new_n886));
  NOR2_X1   g700(.A1(KEYINPUT118), .A2(KEYINPUT48), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n886), .B(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n872), .A2(new_n803), .A3(new_n802), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n889), .B(new_n389), .C1(new_n791), .C2(new_n867), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT117), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n883), .A2(new_n884), .A3(new_n888), .A4(new_n891), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n780), .A2(new_n702), .A3(new_n788), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT112), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n673), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n802), .A2(new_n803), .A3(KEYINPUT112), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n844), .A2(new_n691), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n398), .A2(new_n807), .A3(new_n701), .A4(new_n898), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n653), .B(new_n770), .C1(new_n753), .C2(new_n774), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n893), .A2(new_n654), .A3(new_n899), .A4(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n690), .A2(new_n524), .A3(new_n519), .A4(new_n715), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n902), .B1(new_n631), .B2(new_n652), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n804), .A2(new_n785), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n708), .B(new_n809), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n817), .A2(new_n822), .A3(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n901), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT52), .ZN(new_n908));
  AOI211_X1 g722(.A(new_n698), .B(new_n749), .C1(new_n575), .C2(new_n576), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n740), .A2(new_n787), .A3(new_n706), .A4(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT113), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n910), .B(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n785), .A2(new_n699), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n779), .A2(new_n750), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n722), .A2(new_n751), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n908), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n699), .A2(new_n778), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n721), .A2(new_n706), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n805), .B1(new_n918), .B2(new_n716), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n909), .A2(new_n706), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n920), .A2(new_n911), .A3(new_n740), .A4(new_n787), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n910), .A2(KEYINPUT113), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n919), .A2(new_n923), .A3(KEYINPUT52), .A4(new_n751), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n916), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n907), .A2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT53), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT54), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n907), .A2(new_n925), .A3(KEYINPUT53), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT115), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n907), .A2(KEYINPUT53), .A3(new_n925), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT53), .B1(new_n907), .B2(new_n925), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n936), .A2(KEYINPUT115), .A3(new_n929), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n935), .A2(KEYINPUT114), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n928), .A2(new_n930), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n938), .B1(new_n939), .B2(KEYINPUT114), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n933), .B(new_n937), .C1(new_n940), .C2(new_n929), .ZN(new_n941));
  OAI22_X1  g755(.A1(new_n892), .A2(new_n941), .B1(G952), .B2(G953), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n777), .B(KEYINPUT49), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n743), .A2(new_n807), .A3(new_n386), .A4(new_n382), .ZN(new_n944));
  OR4_X1    g758(.A1(new_n740), .A2(new_n943), .A3(new_n944), .A4(new_n845), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n942), .A2(new_n945), .ZN(G75));
  NOR2_X1   g760(.A1(new_n388), .A2(G952), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n371), .A2(new_n372), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(new_n309), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT55), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n939), .A2(G210), .A3(G902), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT56), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(G902), .B1(new_n934), .B2(new_n935), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(KEYINPUT119), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT119), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n956), .B(G902), .C1(new_n934), .C2(new_n935), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n955), .A2(new_n369), .A3(new_n957), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n950), .A2(new_n952), .ZN(new_n959));
  AOI211_X1 g773(.A(new_n947), .B(new_n953), .C1(new_n958), .C2(new_n959), .ZN(G51));
  INV_X1    g774(.A(new_n947), .ZN(new_n961));
  INV_X1    g775(.A(new_n837), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n955), .A2(new_n962), .A3(new_n957), .ZN(new_n963));
  OAI21_X1  g777(.A(KEYINPUT54), .B1(new_n934), .B2(new_n935), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n931), .ZN(new_n965));
  XNOR2_X1  g779(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(new_n293), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n768), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n961), .B1(new_n963), .B2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT121), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI211_X1 g785(.A(KEYINPUT121), .B(new_n961), .C1(new_n963), .C2(new_n968), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(G54));
  NAND4_X1  g787(.A1(new_n955), .A2(KEYINPUT58), .A3(G475), .A4(new_n957), .ZN(new_n974));
  INV_X1    g788(.A(new_n688), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n974), .A2(new_n975), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n976), .A2(new_n977), .A3(new_n947), .ZN(G60));
  XOR2_X1   g792(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n979));
  NOR2_X1   g793(.A1(new_n517), .A2(new_n188), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n979), .B(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  AOI22_X1  g796(.A1(new_n941), .A2(new_n982), .B1(new_n663), .B2(new_n664), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n663), .A2(new_n664), .A3(new_n982), .ZN(new_n984));
  AND3_X1   g798(.A1(new_n965), .A2(KEYINPUT123), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(KEYINPUT123), .B1(new_n965), .B2(new_n984), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n961), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n983), .A2(new_n987), .ZN(G63));
  NAND2_X1  g802(.A1(G217), .A2(G902), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n989), .B(KEYINPUT60), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n936), .A2(new_n990), .ZN(new_n991));
  OR2_X1    g805(.A1(new_n991), .A2(new_n569), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n697), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n992), .A2(new_n961), .A3(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT61), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n992), .A2(KEYINPUT61), .A3(new_n961), .A4(new_n993), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(G66));
  OAI21_X1  g812(.A(G953), .B1(new_n395), .B2(new_n306), .ZN(new_n999));
  INV_X1    g813(.A(new_n901), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n999), .B1(new_n1000), .B2(G953), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n948), .B1(G898), .B2(new_n388), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1001), .B(new_n1002), .ZN(G69));
  AOI21_X1  g817(.A(new_n711), .B1(new_n190), .B2(G953), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n595), .B(new_n445), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n817), .A2(new_n919), .A3(new_n751), .A4(new_n822), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n814), .A2(new_n807), .A3(new_n787), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n857), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1006), .B1(new_n1008), .B2(new_n842), .ZN(new_n1009));
  AOI21_X1  g823(.A(G953), .B1(new_n1009), .B2(new_n865), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1005), .B1(new_n1010), .B2(new_n711), .ZN(new_n1011));
  OAI21_X1  g825(.A(KEYINPUT62), .B1(new_n746), .B2(new_n915), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(KEYINPUT124), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT124), .ZN(new_n1014));
  OAI211_X1 g828(.A(new_n1014), .B(KEYINPUT62), .C1(new_n746), .C2(new_n915), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  NOR3_X1   g830(.A1(new_n746), .A2(KEYINPUT62), .A3(new_n915), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n653), .A2(new_n809), .ZN(new_n1018));
  INV_X1    g832(.A(new_n898), .ZN(new_n1019));
  NOR3_X1   g833(.A1(new_n1018), .A2(new_n724), .A3(new_n1019), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g835(.A1(new_n1016), .A2(new_n859), .A3(new_n865), .A4(new_n1021), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1005), .B1(new_n1022), .B2(new_n388), .ZN(new_n1023));
  INV_X1    g837(.A(KEYINPUT125), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1011), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  AOI211_X1 g839(.A(KEYINPUT125), .B(new_n1005), .C1(new_n1022), .C2(new_n388), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1004), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AND3_X1   g841(.A1(new_n859), .A2(new_n1021), .A3(new_n865), .ZN(new_n1028));
  AOI21_X1  g842(.A(G953), .B1(new_n1028), .B2(new_n1016), .ZN(new_n1029));
  OAI21_X1  g843(.A(KEYINPUT125), .B1(new_n1029), .B2(new_n1005), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1031));
  INV_X1    g845(.A(new_n1004), .ZN(new_n1032));
  NAND4_X1  g846(.A1(new_n1030), .A2(new_n1031), .A3(new_n1011), .A4(new_n1032), .ZN(new_n1033));
  AND2_X1   g847(.A1(new_n1027), .A2(new_n1033), .ZN(G72));
  NAND3_X1  g848(.A1(new_n1028), .A2(new_n1000), .A3(new_n1016), .ZN(new_n1035));
  XNOR2_X1  g849(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1036));
  NOR2_X1   g850(.A1(new_n717), .A2(new_n188), .ZN(new_n1037));
  XOR2_X1   g851(.A(new_n1036), .B(new_n1037), .Z(new_n1038));
  AND2_X1   g852(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n600), .B1(new_n602), .B2(new_n590), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n643), .A2(new_n1040), .A3(new_n1038), .ZN(new_n1041));
  OAI22_X1  g855(.A1(new_n1039), .A2(new_n1040), .B1(new_n940), .B2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n1009), .A2(new_n865), .A3(new_n1000), .ZN(new_n1043));
  AOI21_X1  g857(.A(new_n643), .B1(new_n1043), .B2(new_n1038), .ZN(new_n1044));
  NOR2_X1   g858(.A1(new_n1044), .A2(new_n947), .ZN(new_n1045));
  OR2_X1    g859(.A1(new_n1045), .A2(KEYINPUT127), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1045), .A2(KEYINPUT127), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n1042), .B1(new_n1046), .B2(new_n1047), .ZN(G57));
endmodule


