//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 1 1 1 0 0 0 1 1 1 1 1 1 0 0 1 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n558,
    new_n560, new_n561, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n625,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G137), .ZN(new_n467));
  INV_X1    g042(.A(G101), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n469), .B1(G2104), .B2(new_n470), .ZN(new_n471));
  NOR3_X1   g046(.A1(new_n463), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n467), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  XNOR2_X1  g050(.A(new_n475), .B(KEYINPUT66), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n477), .B1(new_n464), .B2(new_n465), .ZN(new_n478));
  OAI21_X1  g053(.A(G2105), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI211_X1 g056(.A(KEYINPUT67), .B(G2105), .C1(new_n476), .C2(new_n478), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n474), .B1(new_n481), .B2(new_n482), .ZN(G160));
  AOI21_X1  g058(.A(new_n470), .B1(new_n464), .B2(new_n465), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n488), .B1(G136), .B2(new_n466), .ZN(G162));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n466), .A2(new_n490), .A3(G138), .ZN(new_n491));
  INV_X1    g066(.A(new_n465), .ZN(new_n492));
  NOR2_X1   g067(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n493));
  OAI211_X1 g068(.A(G138), .B(new_n470), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n470), .A2(G114), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n499), .B1(new_n484), .B2(G126), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT69), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n496), .A2(new_n503), .A3(new_n500), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(G164));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(G651), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(KEYINPUT70), .A3(KEYINPUT6), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n509), .A2(KEYINPUT6), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n511), .A2(G543), .A3(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G50), .ZN(new_n516));
  OR2_X1    g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n511), .A2(new_n513), .A3(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G88), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n519), .A2(G62), .ZN(new_n523));
  NAND2_X1  g098(.A1(G75), .A2(G543), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT71), .ZN(new_n525));
  OAI21_X1  g100(.A(G651), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n516), .A2(new_n522), .A3(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  NAND4_X1  g103(.A1(new_n511), .A2(G89), .A3(new_n519), .A4(new_n513), .ZN(new_n529));
  NAND4_X1  g104(.A1(new_n511), .A2(G51), .A3(G543), .A4(new_n513), .ZN(new_n530));
  AND2_X1   g105(.A1(G63), .A2(G651), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT7), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n534), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n519), .A2(new_n531), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  AND3_X1   g111(.A1(new_n529), .A2(new_n530), .A3(new_n536), .ZN(G168));
  AOI21_X1  g112(.A(new_n512), .B1(new_n508), .B2(new_n510), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n538), .A2(G90), .A3(new_n519), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n538), .A2(G52), .A3(G543), .ZN(new_n540));
  INV_X1    g115(.A(G64), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n541), .B1(new_n517), .B2(new_n518), .ZN(new_n542));
  AND2_X1   g117(.A1(G77), .A2(G543), .ZN(new_n543));
  OAI21_X1  g118(.A(G651), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n539), .A2(new_n540), .A3(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  INV_X1    g121(.A(G56), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n547), .B1(new_n517), .B2(new_n518), .ZN(new_n548));
  AND2_X1   g123(.A1(G68), .A2(G543), .ZN(new_n549));
  OAI21_X1  g124(.A(G651), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  XNOR2_X1  g125(.A(KEYINPUT72), .B(G43), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n511), .A2(G543), .A3(new_n513), .A4(new_n551), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n511), .A2(G81), .A3(new_n519), .A4(new_n513), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n550), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(G860), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT73), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT74), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  NAND4_X1  g137(.A1(new_n511), .A2(G91), .A3(new_n519), .A4(new_n513), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT75), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n538), .A2(KEYINPUT75), .A3(G91), .A4(new_n519), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AND2_X1   g142(.A1(G53), .A2(G543), .ZN(new_n568));
  AND4_X1   g143(.A1(KEYINPUT9), .A2(new_n511), .A3(new_n513), .A4(new_n568), .ZN(new_n569));
  AOI21_X1  g144(.A(KEYINPUT9), .B1(new_n538), .B2(new_n568), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n573));
  INV_X1    g148(.A(new_n518), .ZN(new_n574));
  NOR2_X1   g149(.A1(KEYINPUT5), .A2(G543), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n517), .A2(KEYINPUT76), .A3(new_n518), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n572), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n567), .A2(new_n571), .A3(new_n581), .ZN(G299));
  INV_X1    g157(.A(G168), .ZN(G286));
  OAI21_X1  g158(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n584));
  INV_X1    g159(.A(G49), .ZN(new_n585));
  INV_X1    g160(.A(G87), .ZN(new_n586));
  OAI221_X1 g161(.A(new_n584), .B1(new_n514), .B2(new_n585), .C1(new_n586), .C2(new_n520), .ZN(G288));
  NAND2_X1  g162(.A1(new_n515), .A2(G48), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n519), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n589), .A2(new_n509), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n521), .A2(G86), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(G305));
  NAND2_X1  g167(.A1(new_n521), .A2(G85), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n594), .A2(new_n509), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n515), .A2(G47), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n593), .A2(new_n595), .A3(new_n596), .ZN(G290));
  INV_X1    g172(.A(G868), .ZN(new_n598));
  NOR2_X1   g173(.A1(G301), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g174(.A(KEYINPUT77), .B(G66), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  NOR3_X1   g176(.A1(new_n574), .A2(new_n575), .A3(new_n573), .ZN(new_n602));
  AOI21_X1  g177(.A(KEYINPUT76), .B1(new_n517), .B2(new_n518), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT78), .ZN(new_n605));
  NAND2_X1  g180(.A1(G79), .A2(G543), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n600), .B1(new_n576), .B2(new_n577), .ZN(new_n608));
  INV_X1    g183(.A(new_n606), .ZN(new_n609));
  OAI21_X1  g184(.A(KEYINPUT78), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n607), .A2(new_n610), .A3(G651), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  INV_X1    g187(.A(G92), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n520), .B2(new_n613), .ZN(new_n614));
  NAND4_X1  g189(.A1(new_n538), .A2(KEYINPUT10), .A3(G92), .A4(new_n519), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n614), .A2(new_n615), .B1(new_n515), .B2(G54), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT79), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n599), .B1(new_n618), .B2(new_n598), .ZN(G284));
  XOR2_X1   g194(.A(G284), .B(KEYINPUT80), .Z(G321));
  NOR2_X1   g195(.A1(G286), .A2(new_n598), .ZN(new_n621));
  XOR2_X1   g196(.A(G299), .B(KEYINPUT81), .Z(new_n622));
  AOI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(new_n598), .ZN(G297));
  AOI21_X1  g198(.A(new_n621), .B1(new_n622), .B2(new_n598), .ZN(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n618), .B1(new_n625), .B2(G860), .ZN(G148));
  NAND2_X1  g201(.A1(new_n554), .A2(new_n598), .ZN(new_n627));
  AND2_X1   g202(.A1(new_n618), .A2(new_n625), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(new_n598), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g205(.A1(new_n464), .A2(new_n465), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(new_n471), .B2(new_n472), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT12), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT13), .Z(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(G2100), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT82), .ZN(new_n636));
  AOI22_X1  g211(.A1(G123), .A2(new_n484), .B1(new_n466), .B2(G135), .ZN(new_n637));
  OAI21_X1  g212(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n638));
  INV_X1    g213(.A(KEYINPUT83), .ZN(new_n639));
  INV_X1    g214(.A(G111), .ZN(new_n640));
  AOI22_X1  g215(.A1(new_n638), .A2(new_n639), .B1(new_n640), .B2(G2105), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(new_n639), .B2(new_n638), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(G2096), .Z(new_n644));
  OAI211_X1 g219(.A(new_n636), .B(new_n644), .C1(G2100), .C2(new_n634), .ZN(G156));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT84), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2427), .B(G2430), .Z(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(KEYINPUT14), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT85), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n653), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1341), .B(G1348), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n660), .A2(new_n661), .A3(G14), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(G401));
  XOR2_X1   g238(.A(G2072), .B(G2078), .Z(new_n664));
  INV_X1    g239(.A(KEYINPUT87), .ZN(new_n665));
  AND2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  NOR3_X1   g243(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n669), .B1(new_n665), .B2(new_n664), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n664), .A2(KEYINPUT17), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n664), .A2(KEYINPUT17), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n671), .B(new_n672), .C1(new_n667), .C2(new_n668), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n667), .A2(new_n668), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n670), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n674), .A2(new_n664), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT86), .B(KEYINPUT18), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G2096), .B(G2100), .Z(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT88), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n679), .B(new_n681), .ZN(G227));
  XNOR2_X1  g257(.A(G1956), .B(G2474), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT89), .ZN(new_n684));
  XOR2_X1   g259(.A(G1961), .B(G1966), .Z(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT20), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n684), .A2(new_n685), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n692), .A2(new_n688), .A3(new_n686), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n691), .B(new_n693), .C1(new_n688), .C2(new_n692), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1991), .B(G1996), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1981), .B(G1986), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(G229));
  NOR2_X1   g275(.A1(G6), .A2(G16), .ZN(new_n701));
  INV_X1    g276(.A(G305), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n701), .B1(new_n702), .B2(G16), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT32), .B(G1981), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G16), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G22), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G166), .B2(new_n706), .ZN(new_n708));
  INV_X1    g283(.A(G1971), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n705), .A2(new_n710), .ZN(new_n711));
  OR2_X1    g286(.A1(G16), .A2(G23), .ZN(new_n712));
  NAND2_X1  g287(.A1(G288), .A2(KEYINPUT93), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n515), .A2(G49), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n521), .A2(G87), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT93), .ZN(new_n716));
  NAND4_X1  g291(.A1(new_n714), .A2(new_n715), .A3(new_n716), .A4(new_n584), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n712), .B1(new_n718), .B2(new_n706), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT33), .B(G1976), .Z(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n719), .A2(new_n721), .ZN(new_n723));
  NOR3_X1   g298(.A1(new_n711), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT92), .B(KEYINPUT34), .Z(new_n725));
  OR2_X1    g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  INV_X1    g302(.A(G290), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G16), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G16), .B2(G24), .ZN(new_n730));
  INV_X1    g305(.A(G1986), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  INV_X1    g308(.A(G29), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n734), .A2(KEYINPUT90), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(KEYINPUT90), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n737), .A2(G25), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n466), .A2(G131), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n484), .A2(G119), .ZN(new_n740));
  OR2_X1    g315(.A1(G95), .A2(G2105), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n741), .B(G2104), .C1(G107), .C2(new_n470), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n739), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n738), .B1(new_n744), .B2(new_n737), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT35), .B(G1991), .Z(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT91), .Z(new_n747));
  XNOR2_X1  g322(.A(new_n745), .B(new_n747), .ZN(new_n748));
  NOR3_X1   g323(.A1(new_n732), .A2(new_n733), .A3(new_n748), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n726), .A2(new_n727), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT36), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n706), .A2(G5), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G171), .B2(new_n706), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n753), .A2(G1961), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n734), .A2(G33), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n631), .A2(G127), .ZN(new_n756));
  NAND2_X1  g331(.A1(G115), .A2(G2104), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n470), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n466), .A2(G139), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT25), .ZN(new_n762));
  NOR3_X1   g337(.A1(new_n758), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n755), .B1(new_n763), .B2(new_n734), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(G2072), .Z(new_n765));
  NAND3_X1  g340(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT97), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT26), .Z(new_n768));
  AOI22_X1  g343(.A1(G129), .A2(new_n484), .B1(new_n466), .B2(G141), .ZN(new_n769));
  INV_X1    g344(.A(G105), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n769), .B1(new_n770), .B2(new_n473), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n772), .A2(new_n734), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n734), .B2(G32), .ZN(new_n774));
  XOR2_X1   g349(.A(KEYINPUT27), .B(G1996), .Z(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT98), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n765), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  AOI211_X1 g352(.A(new_n754), .B(new_n777), .C1(new_n776), .C2(new_n774), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n737), .A2(G27), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G164), .B2(new_n737), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(G2078), .Z(new_n781));
  INV_X1    g356(.A(KEYINPUT24), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n782), .A2(G34), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n782), .A2(G34), .ZN(new_n784));
  NOR3_X1   g359(.A1(new_n737), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G160), .B2(G29), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n786), .A2(G2084), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT101), .Z(new_n788));
  NAND3_X1  g363(.A1(new_n778), .A2(new_n781), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n706), .A2(G21), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G168), .B2(new_n706), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT99), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n792), .A2(G1966), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(G1966), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT31), .B(G11), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT30), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n796), .A2(G28), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n734), .B1(new_n796), .B2(G28), .ZN(new_n798));
  INV_X1    g373(.A(new_n737), .ZN(new_n799));
  OAI221_X1 g374(.A(new_n795), .B1(new_n797), .B2(new_n798), .C1(new_n643), .C2(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n753), .B2(G1961), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n793), .A2(new_n794), .A3(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n802), .A2(KEYINPUT100), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n802), .A2(KEYINPUT100), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n737), .A2(G35), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G162), .B2(new_n737), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT29), .ZN(new_n807));
  INV_X1    g382(.A(G2090), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n786), .A2(G2084), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n810), .A2(KEYINPUT96), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n810), .A2(KEYINPUT96), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n809), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n706), .A2(G20), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT23), .Z(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(G299), .B2(G16), .ZN(new_n816));
  INV_X1    g391(.A(G1956), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n813), .A2(new_n818), .ZN(new_n819));
  NOR4_X1   g394(.A1(new_n789), .A2(new_n803), .A3(new_n804), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n706), .A2(G4), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n618), .B2(new_n706), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n822), .A2(G1348), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(G1348), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n706), .A2(G19), .ZN(new_n825));
  AND3_X1   g400(.A1(new_n550), .A2(new_n552), .A3(new_n553), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(new_n706), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(G1341), .Z(new_n828));
  NAND2_X1  g403(.A1(new_n799), .A2(G26), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT28), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n466), .A2(G140), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT94), .ZN(new_n832));
  OAI21_X1  g407(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n833));
  INV_X1    g408(.A(G116), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n833), .B1(new_n834), .B2(G2105), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(G128), .B2(new_n484), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n832), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n830), .B1(new_n837), .B2(new_n734), .ZN(new_n838));
  INV_X1    g413(.A(G2067), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n823), .A2(new_n824), .A3(new_n828), .A4(new_n840), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n841), .A2(KEYINPUT95), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(KEYINPUT95), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n751), .A2(new_n820), .A3(new_n842), .A4(new_n843), .ZN(G150));
  INV_X1    g419(.A(G150), .ZN(G311));
  INV_X1    g420(.A(KEYINPUT103), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n554), .A2(KEYINPUT102), .A3(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n846), .B1(new_n554), .B2(KEYINPUT102), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n538), .A2(G93), .A3(new_n519), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n538), .A2(G55), .A3(G543), .ZN(new_n851));
  INV_X1    g426(.A(G67), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n852), .B1(new_n517), .B2(new_n518), .ZN(new_n853));
  AND2_X1   g428(.A1(G80), .A2(G543), .ZN(new_n854));
  OAI21_X1  g429(.A(G651), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n850), .A2(new_n851), .A3(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n554), .A2(KEYINPUT102), .ZN(new_n857));
  OAI22_X1  g432(.A1(new_n848), .A2(new_n849), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT102), .ZN(new_n859));
  OAI21_X1  g434(.A(KEYINPUT103), .B1(new_n826), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n856), .B1(new_n826), .B2(new_n859), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n860), .A2(new_n861), .A3(new_n847), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n858), .A2(new_n862), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(KEYINPUT38), .Z(new_n864));
  NAND2_X1  g439(.A1(new_n618), .A2(G559), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n866), .A2(KEYINPUT39), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(KEYINPUT39), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n867), .A2(new_n555), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n856), .A2(G860), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(KEYINPUT37), .Z(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(G145));
  AND3_X1   g447(.A1(new_n491), .A2(new_n495), .A3(KEYINPUT104), .ZN(new_n873));
  AOI21_X1  g448(.A(KEYINPUT104), .B1(new_n491), .B2(new_n495), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n500), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n837), .B(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(new_n743), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n772), .B(new_n763), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n484), .A2(G130), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n470), .A2(G118), .ZN(new_n880));
  OAI21_X1  g455(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n882), .B1(G142), .B2(new_n466), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n883), .B(new_n633), .Z(new_n884));
  XNOR2_X1  g459(.A(new_n878), .B(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n877), .B(new_n885), .ZN(new_n886));
  XOR2_X1   g461(.A(G160), .B(G162), .Z(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n643), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  XOR2_X1   g464(.A(KEYINPUT105), .B(G37), .Z(new_n890));
  NAND2_X1  g465(.A1(new_n886), .A2(new_n888), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT106), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(KEYINPUT106), .B1(new_n886), .B2(new_n888), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n889), .B(new_n890), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g471(.A(KEYINPUT107), .ZN(new_n897));
  NAND2_X1  g472(.A1(G299), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n567), .A2(new_n571), .A3(KEYINPUT107), .A4(new_n581), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n898), .A2(new_n611), .A3(new_n616), .A4(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n617), .A2(new_n897), .A3(G299), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n618), .A2(new_n625), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(new_n863), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n618), .A2(new_n625), .A3(new_n862), .A4(new_n858), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n902), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n906), .A2(KEYINPUT108), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT109), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n899), .A2(new_n611), .A3(new_n616), .ZN(new_n910));
  OAI21_X1  g485(.A(G65), .B1(new_n602), .B2(new_n603), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(new_n579), .ZN(new_n912));
  AOI22_X1  g487(.A1(new_n912), .A2(G651), .B1(new_n565), .B2(new_n566), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT107), .B1(new_n913), .B2(new_n571), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n617), .A2(new_n897), .A3(G299), .ZN(new_n916));
  OAI21_X1  g491(.A(KEYINPUT41), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT41), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n900), .A2(new_n918), .A3(new_n901), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n909), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n900), .A2(new_n918), .A3(new_n901), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n909), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n905), .B(new_n904), .C1(new_n920), .C2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n904), .A2(new_n905), .ZN(new_n925));
  INV_X1    g500(.A(new_n902), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n925), .A2(KEYINPUT108), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n908), .A2(new_n924), .A3(new_n927), .ZN(new_n928));
  XOR2_X1   g503(.A(G290), .B(G303), .Z(new_n929));
  AOI21_X1  g504(.A(G305), .B1(new_n713), .B2(new_n717), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n713), .A2(new_n717), .A3(G305), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n929), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n930), .ZN(new_n934));
  XNOR2_X1  g509(.A(G290), .B(G303), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n934), .A2(new_n935), .A3(new_n931), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT42), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n928), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n927), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n941), .A2(new_n907), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n942), .A2(new_n924), .A3(new_n938), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n598), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n856), .A2(new_n598), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT110), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n938), .B1(new_n942), .B2(new_n924), .ZN(new_n948));
  AND4_X1   g523(.A1(new_n924), .A2(new_n908), .A3(new_n927), .A4(new_n938), .ZN(new_n949));
  OAI21_X1  g524(.A(G868), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT110), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(new_n951), .A3(new_n945), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n947), .A2(new_n952), .ZN(G295));
  NAND2_X1  g528(.A1(new_n950), .A2(new_n945), .ZN(G331));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n933), .A2(KEYINPUT112), .A3(new_n936), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT112), .B1(new_n933), .B2(new_n936), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(G168), .B(G301), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n858), .A2(new_n862), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n959), .B1(new_n858), .B2(new_n862), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n900), .A2(new_n918), .A3(new_n901), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n918), .B1(new_n900), .B2(new_n901), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT109), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n963), .B1(new_n966), .B2(new_n922), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT111), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n962), .A2(new_n968), .ZN(new_n969));
  AOI211_X1 g544(.A(KEYINPUT111), .B(new_n959), .C1(new_n858), .C2(new_n862), .ZN(new_n970));
  NOR4_X1   g545(.A1(new_n969), .A2(new_n970), .A3(new_n961), .A4(new_n902), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n958), .B1(new_n967), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n963), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n973), .B1(new_n920), .B2(new_n923), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n969), .A2(new_n970), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n961), .A2(new_n902), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n974), .A2(new_n937), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT43), .ZN(new_n979));
  INV_X1    g554(.A(G37), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n972), .A2(new_n978), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT114), .ZN(new_n982));
  INV_X1    g557(.A(new_n962), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n976), .A2(new_n983), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n969), .A2(new_n970), .A3(new_n961), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n964), .A2(new_n965), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n984), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n958), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n988), .A2(new_n978), .A3(new_n890), .ZN(new_n989));
  AOI22_X1  g564(.A1(new_n981), .A2(new_n982), .B1(new_n989), .B2(KEYINPUT43), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n978), .A2(new_n980), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n991), .A2(KEYINPUT114), .A3(new_n979), .A4(new_n972), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n955), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n972), .A2(new_n980), .A3(new_n978), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT113), .B1(new_n994), .B2(KEYINPUT43), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(KEYINPUT43), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n988), .A2(new_n978), .A3(new_n979), .A4(new_n890), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n995), .B1(new_n998), .B2(KEYINPUT113), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n993), .B1(new_n955), .B2(new_n999), .ZN(G397));
  INV_X1    g575(.A(G1384), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n875), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n1003));
  INV_X1    g578(.A(G40), .ZN(new_n1004));
  AOI211_X1 g579(.A(new_n1004), .B(new_n474), .C1(new_n481), .C2(new_n482), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  XOR2_X1   g581(.A(new_n1006), .B(KEYINPUT115), .Z(new_n1007));
  XNOR2_X1  g582(.A(new_n837), .B(G2067), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n772), .B(G1996), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n744), .A2(new_n746), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n744), .A2(new_n746), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(G290), .B(G1986), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1007), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  XOR2_X1   g589(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n1015));
  AOI21_X1  g590(.A(new_n1015), .B1(G303), .B2(G8), .ZN(new_n1016));
  INV_X1    g591(.A(G8), .ZN(new_n1017));
  NOR2_X1   g592(.A1(G166), .A2(new_n1017), .ZN(new_n1018));
  OR2_X1    g593(.A1(KEYINPUT116), .A2(KEYINPUT55), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1016), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n500), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT104), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n496), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n491), .A2(new_n495), .A3(KEYINPUT104), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1021), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT50), .B1(new_n1025), .B2(G1384), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n502), .A2(new_n1027), .A3(new_n1001), .A4(new_n504), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1026), .A2(new_n1005), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT118), .ZN(new_n1030));
  AOI21_X1  g605(.A(G2090), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1026), .A2(KEYINPUT118), .A3(new_n1005), .A4(new_n1028), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n502), .A2(new_n1001), .A3(new_n504), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n1003), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n875), .A2(KEYINPUT45), .A3(new_n1001), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1034), .A2(new_n1005), .A3(new_n1035), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n1031), .A2(new_n1032), .B1(new_n709), .B2(new_n1036), .ZN(new_n1037));
  OAI211_X1 g612(.A(KEYINPUT119), .B(new_n1020), .C1(new_n1037), .C2(new_n1017), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT119), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1028), .A2(new_n1005), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1027), .B1(new_n875), .B2(new_n1001), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1030), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1042), .A2(new_n808), .A3(new_n1032), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1036), .A2(new_n709), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1017), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1020), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1039), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(G160), .A2(G40), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1049));
  AOI21_X1  g624(.A(G1384), .B1(new_n1049), .B2(new_n500), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1048), .B1(new_n1050), .B2(new_n1027), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1033), .A2(KEYINPUT50), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1051), .A2(new_n808), .A3(new_n1052), .ZN(new_n1053));
  AOI211_X1 g628(.A(new_n1017), .B(new_n1020), .C1(new_n1044), .C2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1050), .A2(new_n1005), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n713), .A2(new_n717), .A3(G1976), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1055), .A2(G8), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT52), .ZN(new_n1058));
  INV_X1    g633(.A(G1976), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT52), .B1(G288), .B2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1055), .A2(G8), .A3(new_n1056), .A4(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(G305), .A2(G1981), .ZN(new_n1062));
  XNOR2_X1  g637(.A(KEYINPUT117), .B(G1981), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n588), .A2(new_n590), .A3(new_n591), .A4(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT49), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1062), .A2(KEYINPUT49), .A3(new_n1064), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1067), .A2(G8), .A3(new_n1055), .A4(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1058), .A2(new_n1061), .A3(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1054), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1072), .B1(new_n1036), .B2(G2078), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1048), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n502), .A2(KEYINPUT45), .A3(new_n1001), .A4(new_n504), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1072), .A2(G2078), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n875), .A2(new_n1027), .A3(new_n1001), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1052), .A2(new_n1005), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G1961), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1073), .A2(new_n1077), .A3(new_n1081), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n1082), .A2(G171), .ZN(new_n1083));
  AND4_X1   g658(.A1(new_n1038), .A2(new_n1047), .A3(new_n1071), .A4(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G2084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1051), .A2(new_n1085), .A3(new_n1052), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1005), .B(new_n1075), .C1(new_n1050), .C2(KEYINPUT45), .ZN(new_n1087));
  INV_X1    g662(.A(G1966), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(G8), .ZN(new_n1091));
  NOR2_X1   g666(.A1(G168), .A2(new_n1017), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT51), .B1(new_n1092), .B2(KEYINPUT125), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1091), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1094), .ZN(new_n1096));
  OAI211_X1 g671(.A(G8), .B(new_n1096), .C1(new_n1090), .C2(G286), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1099));
  AOI21_X1  g674(.A(KEYINPUT62), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT62), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1099), .ZN(new_n1102));
  AOI211_X1 g677(.A(new_n1101), .B(new_n1102), .C1(new_n1095), .C2(new_n1097), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1084), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(G1348), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1079), .A2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1002), .A2(new_n1048), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n839), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n617), .B(KEYINPUT124), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1106), .A2(KEYINPUT60), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT60), .ZN(new_n1111));
  AOI21_X1  g686(.A(G1348), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1108), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  AOI221_X4 g689(.A(new_n1111), .B1(new_n1107), .B2(new_n839), .C1(new_n1079), .C2(new_n1105), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT124), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n617), .A2(new_n1116), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1110), .B(new_n1114), .C1(new_n1115), .C2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT61), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n817), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1120));
  XNOR2_X1  g695(.A(KEYINPUT56), .B(G2072), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1121), .B(KEYINPUT123), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1034), .A2(new_n1005), .A3(new_n1035), .A4(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT57), .B1(new_n913), .B2(KEYINPUT122), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(G299), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n913), .B(new_n571), .C1(KEYINPUT122), .C2(KEYINPUT57), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1120), .A2(new_n1123), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1127), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1119), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(G1996), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1034), .A2(new_n1132), .A3(new_n1005), .A4(new_n1035), .ZN(new_n1133));
  XOR2_X1   g708(.A(KEYINPUT58), .B(G1341), .Z(new_n1134));
  NAND2_X1  g709(.A1(new_n1055), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT59), .B1(new_n1136), .B2(new_n826), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT59), .ZN(new_n1138));
  AOI211_X1 g713(.A(new_n1138), .B(new_n554), .C1(new_n1133), .C2(new_n1135), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1130), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1141), .A2(new_n1128), .A3(KEYINPUT61), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1118), .A2(new_n1131), .A3(new_n1140), .A4(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n617), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1130), .B1(new_n1144), .B2(new_n1128), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(G301), .B(KEYINPUT54), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1082), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT126), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1081), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n474), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1151), .A2(G40), .A3(new_n479), .A4(new_n1076), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1152), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1147), .B1(new_n1153), .B2(new_n1035), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1079), .A2(KEYINPUT126), .A3(new_n1080), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1150), .A2(new_n1073), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1148), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1157), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1047), .A2(new_n1038), .A3(new_n1071), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1146), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(G288), .A2(G1976), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1069), .A2(new_n1161), .ZN(new_n1162));
  AOI211_X1 g737(.A(new_n1017), .B(new_n1107), .C1(new_n1162), .C2(new_n1064), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1070), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1163), .B1(new_n1054), .B2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1104), .A2(new_n1160), .A3(new_n1165), .ZN(new_n1166));
  AOI211_X1 g741(.A(new_n1017), .B(G286), .C1(new_n1086), .C2(new_n1089), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1017), .B1(new_n1044), .B2(new_n1053), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1168), .ZN(new_n1169));
  OAI211_X1 g744(.A(new_n1167), .B(new_n1164), .C1(new_n1169), .C2(new_n1020), .ZN(new_n1170));
  OAI21_X1  g745(.A(KEYINPUT63), .B1(new_n1168), .B2(new_n1046), .ZN(new_n1171));
  OAI21_X1  g746(.A(KEYINPUT121), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1079), .A2(G2084), .ZN(new_n1173));
  AOI21_X1  g748(.A(G1966), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1174));
  OAI211_X1 g749(.A(G8), .B(G168), .C1(new_n1173), .C2(new_n1174), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n1054), .A2(new_n1175), .A3(new_n1070), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT121), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1171), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1172), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1176), .A2(new_n1038), .A3(new_n1047), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT120), .ZN(new_n1182));
  AOI21_X1  g757(.A(KEYINPUT63), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1176), .A2(new_n1038), .A3(new_n1047), .A4(KEYINPUT120), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1180), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1014), .B1(new_n1166), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n837), .A2(new_n839), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1187), .B1(new_n1188), .B2(new_n1010), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1189), .A2(new_n1007), .ZN(new_n1190));
  XOR2_X1   g765(.A(new_n1190), .B(KEYINPUT127), .Z(new_n1191));
  NAND3_X1  g766(.A1(new_n1007), .A2(new_n731), .A3(new_n728), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT48), .ZN(new_n1193));
  OR2_X1    g768(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1007), .A2(new_n1012), .ZN(new_n1196));
  AND3_X1   g771(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1007), .A2(new_n1132), .ZN(new_n1198));
  XNOR2_X1  g773(.A(new_n1198), .B(KEYINPUT46), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1008), .A2(new_n772), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1007), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  OR2_X1    g777(.A1(new_n1202), .A2(KEYINPUT47), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1202), .A2(KEYINPUT47), .ZN(new_n1204));
  AOI211_X1 g779(.A(new_n1191), .B(new_n1197), .C1(new_n1203), .C2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1186), .A2(new_n1205), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g781(.A1(G227), .A2(new_n460), .ZN(new_n1208));
  NAND2_X1  g782(.A1(new_n662), .A2(new_n1208), .ZN(new_n1209));
  NOR2_X1   g783(.A1(G229), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g784(.A(KEYINPUT113), .ZN(new_n1211));
  AOI21_X1  g785(.A(new_n1211), .B1(new_n996), .B2(new_n997), .ZN(new_n1212));
  OAI211_X1 g786(.A(new_n1210), .B(new_n895), .C1(new_n1212), .C2(new_n995), .ZN(G225));
  INV_X1    g787(.A(G225), .ZN(G308));
endmodule


