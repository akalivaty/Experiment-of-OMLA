//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 1 0 1 0 1 1 1 1 0 1 0 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n557, new_n558, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n630,
    new_n631, new_n634, new_n636, new_n637, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1185;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT65), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n456), .A2(KEYINPUT67), .ZN(new_n457));
  AOI21_X1  g032(.A(new_n457), .B1(G567), .B2(new_n453), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(KEYINPUT67), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT68), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(G137), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n469));
  XNOR2_X1  g044(.A(new_n469), .B(KEYINPUT69), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n467), .A2(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n466), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n471), .A2(new_n474), .ZN(G160));
  AND2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n466), .A2(G112), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT70), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n466), .A2(new_n478), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(G124), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n484), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n485), .A2(KEYINPUT70), .A3(G124), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n483), .B1(new_n488), .B2(new_n489), .ZN(G162));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(G2105), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n466), .A2(G138), .A3(new_n467), .ZN(new_n494));
  NAND2_X1  g069(.A1(KEYINPUT71), .A2(KEYINPUT4), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(G126), .A2(G2105), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n463), .A2(new_n465), .ZN(new_n498));
  NAND3_X1  g073(.A1(KEYINPUT71), .A2(KEYINPUT4), .A3(G138), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(new_n467), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  INV_X1    g078(.A(KEYINPUT6), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT72), .B1(new_n504), .B2(G651), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT72), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n506), .A2(new_n507), .A3(KEYINPUT6), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  OR2_X1    g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n504), .A2(G651), .ZN(new_n513));
  NAND4_X1  g088(.A1(new_n509), .A2(G88), .A3(new_n512), .A4(new_n513), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n509), .A2(G50), .A3(G543), .A4(new_n513), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT73), .ZN(new_n516));
  AND3_X1   g091(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n516), .B1(new_n514), .B2(new_n515), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n517), .A2(new_n518), .B1(new_n507), .B2(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  AOI22_X1  g096(.A1(new_n505), .A2(new_n508), .B1(new_n504), .B2(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n522), .A2(G51), .A3(G543), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT74), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n510), .A2(new_n524), .A3(new_n511), .ZN(new_n525));
  AND2_X1   g100(.A1(KEYINPUT5), .A2(G543), .ZN(new_n526));
  NOR2_X1   g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  OAI21_X1  g102(.A(KEYINPUT74), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n525), .A2(new_n528), .A3(G63), .A4(G651), .ZN(new_n529));
  NAND4_X1  g104(.A1(new_n509), .A2(G89), .A3(new_n512), .A4(new_n513), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  AND4_X1   g107(.A1(new_n523), .A2(new_n529), .A3(new_n530), .A4(new_n532), .ZN(G168));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n525), .A2(new_n528), .ZN(new_n535));
  INV_X1    g110(.A(G64), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G651), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n509), .A2(G52), .A3(G543), .A4(new_n513), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n509), .A2(G90), .A3(new_n512), .A4(new_n513), .ZN(new_n540));
  AND3_X1   g115(.A1(new_n539), .A2(new_n540), .A3(KEYINPUT75), .ZN(new_n541));
  AOI21_X1  g116(.A(KEYINPUT75), .B1(new_n539), .B2(new_n540), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n538), .B1(new_n541), .B2(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  NAND4_X1  g119(.A1(new_n509), .A2(G43), .A3(G543), .A4(new_n513), .ZN(new_n545));
  NAND4_X1  g120(.A1(new_n509), .A2(G81), .A3(new_n512), .A4(new_n513), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n525), .A2(new_n528), .A3(G56), .ZN(new_n548));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n507), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT76), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n547), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AND2_X1   g127(.A1(new_n550), .A2(new_n551), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  NAND4_X1  g134(.A1(new_n509), .A2(G53), .A3(G543), .A4(new_n513), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(KEYINPUT9), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n522), .A2(new_n562), .A3(G53), .A4(G543), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT77), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n566), .B1(new_n510), .B2(new_n511), .ZN(new_n567));
  AND2_X1   g142(.A1(G78), .A2(G543), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n509), .A2(G91), .A3(new_n512), .A4(new_n513), .ZN(new_n570));
  AND2_X1   g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AND3_X1   g146(.A1(new_n564), .A2(new_n565), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n565), .B1(new_n564), .B2(new_n571), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n572), .A2(new_n573), .ZN(G299));
  INV_X1    g149(.A(G168), .ZN(G286));
  INV_X1    g150(.A(KEYINPUT78), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n509), .A2(new_n512), .A3(new_n513), .ZN(new_n577));
  INV_X1    g152(.A(G87), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n522), .A2(KEYINPUT78), .A3(G87), .A4(new_n512), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n522), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n579), .A2(new_n580), .B1(new_n582), .B2(G49), .ZN(new_n583));
  INV_X1    g158(.A(G74), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n535), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT79), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n585), .A2(new_n586), .A3(G651), .ZN(new_n587));
  AOI21_X1  g162(.A(G74), .B1(new_n525), .B2(new_n528), .ZN(new_n588));
  OAI21_X1  g163(.A(KEYINPUT79), .B1(new_n588), .B2(new_n507), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n583), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT80), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n583), .A2(new_n590), .A3(KEYINPUT80), .ZN(new_n594));
  AND2_X1   g169(.A1(new_n593), .A2(new_n594), .ZN(G288));
  INV_X1    g170(.A(G61), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n596), .B1(new_n510), .B2(new_n511), .ZN(new_n597));
  AND2_X1   g172(.A1(G73), .A2(G543), .ZN(new_n598));
  OAI21_X1  g173(.A(G651), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND4_X1  g174(.A1(new_n509), .A2(G48), .A3(G543), .A4(new_n513), .ZN(new_n600));
  AND2_X1   g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n509), .A2(G86), .A3(new_n512), .A4(new_n513), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(G305));
  NAND2_X1  g178(.A1(G72), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G60), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n535), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(G651), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n522), .A2(G47), .A3(G543), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n522), .A2(G85), .A3(new_n512), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT81), .ZN(new_n610));
  AND3_X1   g185(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n610), .B1(new_n608), .B2(new_n609), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n607), .B1(new_n611), .B2(new_n612), .ZN(G290));
  NAND2_X1  g188(.A1(G301), .A2(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(G79), .A2(G543), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n526), .A2(new_n527), .ZN(new_n616));
  INV_X1    g191(.A(G66), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G651), .ZN(new_n619));
  INV_X1    g194(.A(G54), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(new_n581), .ZN(new_n621));
  NAND4_X1  g196(.A1(new_n509), .A2(G92), .A3(new_n512), .A4(new_n513), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT10), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n621), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n614), .B1(G868), .B2(new_n626), .ZN(G284));
  OAI21_X1  g202(.A(new_n614), .B1(G868), .B2(new_n626), .ZN(G321));
  INV_X1    g203(.A(G868), .ZN(new_n629));
  NOR2_X1   g204(.A1(G286), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(G299), .B(KEYINPUT82), .Z(new_n631));
  AOI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(new_n629), .ZN(G297));
  AOI21_X1  g207(.A(new_n630), .B1(new_n631), .B2(new_n629), .ZN(G280));
  INV_X1    g208(.A(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n626), .B1(new_n634), .B2(G860), .ZN(G148));
  NAND2_X1  g210(.A1(new_n626), .A2(new_n634), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G868), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g213(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g214(.A1(new_n462), .A2(G2104), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n478), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT83), .B(KEYINPUT12), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(KEYINPUT84), .B(KEYINPUT13), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(G2100), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  AOI22_X1  g223(.A1(new_n485), .A2(G123), .B1(new_n479), .B2(G135), .ZN(new_n649));
  INV_X1    g224(.A(G111), .ZN(new_n650));
  INV_X1    g225(.A(KEYINPUT85), .ZN(new_n651));
  OAI21_X1  g226(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n652));
  AOI22_X1  g227(.A1(new_n498), .A2(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(new_n651), .B2(new_n652), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n649), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(G2096), .Z(new_n656));
  NAND3_X1  g231(.A1(new_n647), .A2(new_n648), .A3(new_n656), .ZN(G156));
  XOR2_X1   g232(.A(G1341), .B(G1348), .Z(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT86), .Z(new_n659));
  XOR2_X1   g234(.A(G2451), .B(G2454), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n659), .B(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT14), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2427), .B(G2438), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2430), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT15), .B(G2435), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n663), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n667), .B1(new_n666), .B2(new_n665), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n662), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2443), .B(G2446), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n670), .ZN(new_n672));
  AND3_X1   g247(.A1(new_n671), .A2(G14), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT87), .ZN(G401));
  XOR2_X1   g249(.A(KEYINPUT88), .B(KEYINPUT18), .Z(new_n675));
  XOR2_X1   g250(.A(G2084), .B(G2090), .Z(new_n676));
  XNOR2_X1  g251(.A(G2067), .B(G2678), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(KEYINPUT17), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n676), .A2(new_n677), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n675), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G2072), .B(G2078), .Z(new_n682));
  INV_X1    g257(.A(new_n675), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n682), .B1(new_n678), .B2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n681), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G2096), .B(G2100), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G227));
  XOR2_X1   g262(.A(G1971), .B(G1976), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT19), .ZN(new_n689));
  XOR2_X1   g264(.A(G1956), .B(G2474), .Z(new_n690));
  XOR2_X1   g265(.A(G1961), .B(G1966), .Z(new_n691));
  AND2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT20), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n690), .A2(new_n691), .ZN(new_n695));
  NOR3_X1   g270(.A1(new_n689), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n689), .B2(new_n695), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1991), .B(G1996), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1981), .B(G1986), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(G229));
  NAND3_X1  g279(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT93), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT25), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n479), .A2(G139), .ZN(new_n708));
  AOI22_X1  g283(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT94), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n466), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n710), .B2(new_n709), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n707), .A2(new_n708), .A3(new_n712), .ZN(new_n713));
  MUX2_X1   g288(.A(G33), .B(new_n713), .S(G29), .Z(new_n714));
  OR2_X1    g289(.A1(new_n714), .A2(G2072), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(G2072), .ZN(new_n716));
  NAND2_X1  g291(.A1(G160), .A2(G29), .ZN(new_n717));
  INV_X1    g292(.A(G34), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n718), .A2(KEYINPUT24), .ZN(new_n719));
  AOI21_X1  g294(.A(G29), .B1(new_n718), .B2(KEYINPUT24), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(KEYINPUT95), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(KEYINPUT95), .B2(new_n720), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n717), .A2(G2084), .A3(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G32), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT96), .B(KEYINPUT26), .Z(new_n726));
  NAND3_X1  g301(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n485), .A2(G129), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n479), .A2(G141), .ZN(new_n731));
  AND4_X1   g306(.A1(new_n728), .A2(new_n729), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n725), .B1(new_n732), .B2(new_n724), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT27), .B(G1996), .Z(new_n734));
  NOR2_X1   g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT97), .Z(new_n736));
  NAND4_X1  g311(.A1(new_n715), .A2(new_n716), .A3(new_n723), .A4(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT98), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G16), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G20), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT23), .Z(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G299), .B2(G16), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G1956), .ZN(new_n744));
  NOR2_X1   g319(.A1(G171), .A2(new_n740), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G5), .B2(new_n740), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G1961), .ZN(new_n748));
  INV_X1    g323(.A(G28), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n749), .A2(KEYINPUT30), .ZN(new_n750));
  AOI21_X1  g325(.A(G29), .B1(new_n749), .B2(KEYINPUT30), .ZN(new_n751));
  OR2_X1    g326(.A1(KEYINPUT31), .A2(G11), .ZN(new_n752));
  NAND2_X1  g327(.A1(KEYINPUT31), .A2(G11), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n750), .A2(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n655), .B2(new_n724), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n740), .A2(G21), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G168), .B2(new_n740), .ZN(new_n757));
  AND2_X1   g332(.A1(new_n757), .A2(G1966), .ZN(new_n758));
  NOR2_X1   g333(.A1(G164), .A2(new_n724), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G27), .B2(new_n724), .ZN(new_n760));
  INV_X1    g335(.A(G2078), .ZN(new_n761));
  AOI211_X1 g336(.A(new_n755), .B(new_n758), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n748), .B(new_n762), .C1(G1966), .C2(new_n757), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n724), .A2(G26), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT28), .Z(new_n765));
  NAND2_X1  g340(.A1(new_n479), .A2(G140), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT92), .ZN(new_n767));
  OAI221_X1 g342(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n466), .C2(G116), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n485), .A2(G128), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n765), .B1(new_n770), .B2(G29), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G2067), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n724), .A2(G35), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G162), .B2(new_n724), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT29), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n775), .A2(G2090), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n772), .B(new_n776), .C1(new_n761), .C2(new_n760), .ZN(new_n777));
  NOR2_X1   g352(.A1(G4), .A2(G16), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT91), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n625), .A2(new_n624), .ZN(new_n780));
  INV_X1    g355(.A(new_n621), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n779), .B1(new_n782), .B2(new_n740), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1348), .ZN(new_n784));
  NOR2_X1   g359(.A1(G16), .A2(G19), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n554), .B2(G16), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n786), .A2(G1341), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(G1341), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n784), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n775), .A2(G2090), .ZN(new_n790));
  NOR4_X1   g365(.A1(new_n763), .A2(new_n777), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(G2084), .B1(new_n717), .B2(new_n722), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n733), .B2(new_n734), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n747), .B2(G1961), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT99), .Z(new_n795));
  NAND4_X1  g370(.A1(new_n739), .A2(new_n744), .A3(new_n791), .A4(new_n795), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n724), .A2(G25), .ZN(new_n797));
  OAI221_X1 g372(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n466), .C2(G107), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT89), .Z(new_n799));
  AOI22_X1  g374(.A1(new_n485), .A2(G119), .B1(new_n479), .B2(G131), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n797), .B1(new_n801), .B2(G29), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT35), .B(G1991), .Z(new_n803));
  XOR2_X1   g378(.A(new_n802), .B(new_n803), .Z(new_n804));
  INV_X1    g379(.A(G1986), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n740), .A2(G24), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G290), .B2(G16), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n804), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n805), .B2(new_n807), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n740), .A2(G6), .ZN(new_n810));
  INV_X1    g385(.A(G305), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(new_n740), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT32), .B(G1981), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n740), .A2(G23), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n591), .B2(G16), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT33), .B(G1976), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(G166), .A2(G16), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G16), .B2(G22), .ZN(new_n821));
  INV_X1    g396(.A(G1971), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n821), .A2(new_n822), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n816), .A2(new_n817), .ZN(new_n825));
  NOR4_X1   g400(.A1(new_n819), .A2(new_n823), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT90), .B(KEYINPUT34), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n827), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n809), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n830), .A2(KEYINPUT36), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(KEYINPUT36), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n796), .B1(new_n831), .B2(new_n832), .ZN(G311));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  INV_X1    g409(.A(new_n796), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(G150));
  NAND2_X1  g411(.A1(new_n626), .A2(G559), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT38), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n509), .A2(G55), .A3(G543), .A4(new_n513), .ZN(new_n839));
  INV_X1    g414(.A(G93), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(new_n577), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n525), .A2(new_n528), .A3(G67), .ZN(new_n842));
  NAND2_X1  g417(.A1(G80), .A2(G543), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n507), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(new_n552), .B2(new_n553), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n548), .A2(new_n549), .ZN(new_n847));
  OAI21_X1  g422(.A(KEYINPUT76), .B1(new_n847), .B2(new_n507), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n841), .A2(new_n844), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n550), .A2(new_n551), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n848), .A2(new_n849), .A3(new_n850), .A4(new_n547), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n846), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n838), .B(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT39), .ZN(new_n854));
  AOI21_X1  g429(.A(G860), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(new_n854), .B2(new_n853), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT100), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n845), .A2(G860), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT37), .Z(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(G145));
  XNOR2_X1  g435(.A(new_n655), .B(G160), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(G162), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n713), .B(new_n732), .ZN(new_n863));
  AOI22_X1  g438(.A1(new_n485), .A2(G130), .B1(new_n479), .B2(G142), .ZN(new_n864));
  OAI221_X1 g439(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n466), .C2(G118), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n801), .B(new_n866), .Z(new_n867));
  OR2_X1    g442(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n770), .B(new_n502), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n643), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n863), .A2(new_n867), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n868), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n870), .B1(new_n868), .B2(new_n871), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n862), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(G37), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n863), .B(new_n867), .ZN(new_n877));
  INV_X1    g452(.A(new_n870), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n862), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(new_n880), .A3(new_n872), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n875), .A2(new_n876), .A3(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n884), .B1(new_n849), .B2(G868), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n852), .B(new_n636), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n782), .B1(new_n572), .B2(new_n573), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n564), .A2(new_n571), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(KEYINPUT77), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n564), .A2(new_n565), .A3(new_n571), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(new_n890), .A3(new_n626), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n886), .A2(new_n892), .ZN(new_n893));
  AND3_X1   g468(.A1(new_n887), .A2(new_n891), .A3(KEYINPUT41), .ZN(new_n894));
  AOI21_X1  g469(.A(KEYINPUT41), .B1(new_n887), .B2(new_n891), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n893), .B1(new_n886), .B2(new_n896), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n897), .A2(KEYINPUT42), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(KEYINPUT42), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(G166), .A2(new_n591), .ZN(new_n901));
  NAND3_X1  g476(.A1(G303), .A2(new_n590), .A3(new_n583), .ZN(new_n902));
  NAND2_X1  g477(.A1(G290), .A2(new_n811), .ZN(new_n903));
  OAI211_X1 g478(.A(G305), .B(new_n607), .C1(new_n611), .C2(new_n612), .ZN(new_n904));
  AOI22_X1  g479(.A1(new_n901), .A2(new_n902), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n901), .A2(new_n903), .A3(new_n904), .A4(new_n902), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n629), .B1(new_n900), .B2(new_n908), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n898), .A2(new_n907), .A3(new_n906), .A4(new_n899), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n885), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n909), .A2(new_n910), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n911), .B1(KEYINPUT101), .B2(new_n912), .ZN(G295));
  AOI21_X1  g488(.A(new_n911), .B1(KEYINPUT101), .B2(new_n912), .ZN(G331));
  INV_X1    g489(.A(KEYINPUT108), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n846), .A2(new_n851), .ZN(new_n916));
  NAND2_X1  g491(.A1(G301), .A2(G286), .ZN(new_n917));
  OAI211_X1 g492(.A(G168), .B(new_n538), .C1(new_n542), .C2(new_n541), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n916), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n846), .A2(new_n917), .A3(new_n851), .A4(new_n918), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(KEYINPUT105), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n917), .A2(new_n918), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n852), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT104), .ZN(new_n927));
  AOI22_X1  g502(.A1(new_n846), .A2(new_n851), .B1(new_n917), .B2(new_n918), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT104), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n924), .A2(new_n892), .A3(new_n927), .A4(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n852), .A2(new_n925), .ZN(new_n932));
  OAI22_X1  g507(.A1(new_n894), .A2(new_n895), .B1(new_n932), .B2(new_n928), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT103), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n926), .A2(new_n922), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n936), .B(KEYINPUT103), .C1(new_n894), .C2(new_n895), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n931), .A2(new_n935), .A3(new_n908), .A4(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(new_n876), .ZN(new_n939));
  OR2_X1    g514(.A1(new_n894), .A2(new_n895), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n920), .B1(new_n916), .B2(new_n919), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n922), .A2(KEYINPUT105), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n927), .A2(new_n930), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n940), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n926), .A2(new_n892), .A3(new_n922), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT106), .ZN(new_n949));
  INV_X1    g524(.A(new_n907), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n949), .B1(new_n950), .B2(new_n905), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n906), .A2(KEYINPUT106), .A3(new_n907), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n947), .A2(new_n948), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n946), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n927), .B(new_n930), .C1(new_n941), .C2(new_n942), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n956), .B1(new_n957), .B2(new_n940), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT107), .B1(new_n958), .B2(new_n953), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n939), .B1(new_n955), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT43), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n915), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n938), .A2(new_n876), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n948), .B1(new_n947), .B2(new_n954), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n958), .A2(KEYINPUT107), .A3(new_n953), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n966), .A2(KEYINPUT108), .A3(KEYINPUT43), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n931), .A2(new_n935), .A3(new_n937), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n969), .A2(new_n954), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n970), .A2(new_n939), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n968), .B1(new_n971), .B2(new_n961), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n962), .A2(new_n967), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT43), .B1(new_n970), .B2(new_n939), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n974), .B1(new_n966), .B2(KEYINPUT43), .ZN(new_n975));
  XOR2_X1   g550(.A(KEYINPUT102), .B(KEYINPUT44), .Z(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n973), .A2(new_n977), .ZN(G397));
  INV_X1    g553(.A(G1976), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n593), .A2(new_n979), .A3(new_n594), .ZN(new_n980));
  XOR2_X1   g555(.A(KEYINPUT113), .B(G8), .Z(new_n981));
  AOI21_X1  g556(.A(G1384), .B1(new_n496), .B2(new_n501), .ZN(new_n982));
  INV_X1    g557(.A(G40), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n471), .A2(new_n474), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n981), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n583), .A2(new_n590), .A3(G1976), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n980), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n987), .B1(new_n985), .B2(new_n986), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT114), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AOI211_X1 g567(.A(KEYINPUT114), .B(new_n987), .C1(new_n985), .C2(new_n986), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n989), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G1981), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n599), .A2(new_n602), .A3(new_n600), .A4(new_n995), .ZN(new_n996));
  OR2_X1    g571(.A1(new_n996), .A2(KEYINPUT115), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(KEYINPUT115), .ZN(new_n998));
  XOR2_X1   g573(.A(KEYINPUT116), .B(G86), .Z(new_n999));
  OAI21_X1  g574(.A(new_n601), .B1(new_n577), .B2(new_n999), .ZN(new_n1000));
  AOI22_X1  g575(.A1(new_n997), .A2(new_n998), .B1(new_n1000), .B2(G1981), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT49), .B1(new_n1001), .B2(KEYINPUT117), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT117), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT49), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n1000), .A2(G1981), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT115), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n996), .B(new_n1006), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1003), .B(new_n1004), .C1(new_n1005), .C2(new_n1007), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n1002), .A2(new_n985), .A3(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n994), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(G303), .A2(G8), .ZN(new_n1012));
  XNOR2_X1  g587(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n1013));
  OR2_X1    g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT55), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1012), .B1(KEYINPUT112), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G1384), .ZN(new_n1018));
  INV_X1    g593(.A(new_n501), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n463), .B(new_n465), .C1(new_n476), .C2(new_n477), .ZN(new_n1020));
  INV_X1    g595(.A(G138), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n495), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n493), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1018), .B1(new_n1019), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT50), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n982), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G2090), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1026), .A2(new_n1028), .A3(new_n1029), .A4(new_n984), .ZN(new_n1030));
  INV_X1    g605(.A(new_n474), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1031), .A2(G40), .A3(new_n470), .A4(new_n468), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT45), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1032), .B1(new_n1025), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n982), .A2(KEYINPUT45), .ZN(new_n1035));
  AOI21_X1  g610(.A(G1971), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1030), .B1(new_n1036), .B2(KEYINPUT111), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n984), .B1(new_n982), .B2(KEYINPUT45), .ZN(new_n1038));
  AOI211_X1 g613(.A(new_n1033), .B(G1384), .C1(new_n496), .C2(new_n501), .ZN(new_n1039));
  OAI211_X1 g614(.A(KEYINPUT111), .B(new_n822), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  OAI211_X1 g616(.A(G8), .B(new_n1017), .C1(new_n1037), .C2(new_n1041), .ZN(new_n1042));
  XOR2_X1   g617(.A(new_n1007), .B(KEYINPUT119), .Z(new_n1043));
  NAND3_X1  g618(.A1(new_n1002), .A2(new_n985), .A3(new_n1008), .ZN(new_n1044));
  NOR2_X1   g619(.A1(G288), .A2(G1976), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g621(.A(new_n985), .B(KEYINPUT118), .Z(new_n1047));
  OAI22_X1  g622(.A1(new_n1011), .A2(new_n1042), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g623(.A(KEYINPUT124), .B(KEYINPUT54), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1025), .A2(new_n1033), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1050), .A2(new_n1035), .A3(new_n761), .A4(new_n984), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1026), .A2(new_n1028), .A3(new_n984), .ZN(new_n1053));
  XNOR2_X1  g628(.A(KEYINPUT125), .B(G1961), .ZN(new_n1054));
  AOI22_X1  g629(.A1(new_n1051), .A2(new_n1052), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NOR3_X1   g630(.A1(new_n1032), .A2(new_n1052), .A3(G2078), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1056), .A2(new_n1050), .A3(new_n1035), .ZN(new_n1057));
  AOI21_X1  g632(.A(G301), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n982), .A2(KEYINPUT109), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1033), .B1(new_n982), .B2(KEYINPUT109), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1035), .B(new_n1056), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1063));
  AND4_X1   g638(.A1(G301), .A2(new_n1059), .A3(new_n1060), .A4(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1049), .B1(new_n1058), .B2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1059), .A2(new_n1063), .A3(new_n1060), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(G171), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1055), .A2(G301), .A3(new_n1057), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1067), .A2(new_n1068), .A3(KEYINPUT54), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1065), .A2(new_n1069), .ZN(new_n1070));
  AND2_X1   g645(.A1(new_n985), .A2(new_n986), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT114), .B1(new_n1071), .B2(new_n987), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n990), .A2(new_n991), .ZN(new_n1073));
  AOI22_X1  g648(.A1(new_n1072), .A2(new_n1073), .B1(new_n980), .B2(new_n988), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1075));
  INV_X1    g650(.A(new_n981), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1030), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1076), .B1(new_n1077), .B2(new_n1036), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1042), .A2(new_n1074), .A3(new_n1079), .A4(new_n1044), .ZN(new_n1080));
  INV_X1    g655(.A(G1966), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1082));
  XOR2_X1   g657(.A(KEYINPUT120), .B(G2084), .Z(new_n1083));
  NAND4_X1  g658(.A1(new_n1026), .A2(new_n1028), .A3(new_n984), .A4(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n1076), .ZN(new_n1086));
  NOR2_X1   g661(.A1(G168), .A2(new_n981), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1087), .A2(KEYINPUT51), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G8), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1090), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT51), .B1(new_n1091), .B2(new_n1087), .ZN(new_n1092));
  AOI211_X1 g667(.A(G168), .B(new_n981), .C1(new_n1082), .C2(new_n1084), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1089), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1070), .A2(new_n1080), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(G1956), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1053), .A2(new_n1096), .ZN(new_n1097));
  XOR2_X1   g672(.A(new_n888), .B(KEYINPUT57), .Z(new_n1098));
  XNOR2_X1  g673(.A(KEYINPUT56), .B(G2072), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1034), .A2(new_n1035), .A3(new_n1099), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n1097), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(G1348), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1053), .A2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1025), .A2(new_n1032), .ZN(new_n1104));
  INV_X1    g679(.A(G2067), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n1101), .A2(new_n1107), .A3(new_n782), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1109));
  OR2_X1    g684(.A1(new_n1109), .A2(KEYINPUT122), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1098), .B1(new_n1109), .B2(KEYINPUT122), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1108), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1038), .A2(G1996), .A3(new_n1039), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT58), .B(G1341), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1104), .A2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n554), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n1117));
  OR3_X1    g692(.A1(new_n1116), .A2(KEYINPUT123), .A3(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1116), .B1(KEYINPUT123), .B2(new_n1117), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT61), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1118), .B(new_n1119), .C1(new_n1120), .C2(new_n1101), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT60), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n782), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(new_n1123), .B2(new_n1122), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1098), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1120), .B1(new_n1101), .B2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1107), .A2(KEYINPUT60), .A3(new_n782), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1125), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1112), .B1(new_n1121), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1048), .B1(new_n1095), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT63), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1085), .A2(G168), .A3(new_n1076), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1132), .B1(new_n1080), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT121), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1136), .B(new_n1132), .C1(new_n1080), .C2(new_n1133), .ZN(new_n1137));
  OAI21_X1  g712(.A(G8), .B1(new_n1037), .B2(new_n1041), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n1075), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1133), .A2(new_n1132), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1139), .A2(new_n1010), .A3(new_n1042), .A4(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1135), .A2(new_n1137), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1080), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1094), .A2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1143), .A2(new_n1145), .A3(KEYINPUT126), .A4(new_n1058), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT126), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1010), .A2(new_n1042), .A3(new_n1079), .A4(new_n1058), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1085), .A2(G286), .A3(new_n1076), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1149), .B(KEYINPUT51), .C1(new_n1087), .C2(new_n1091), .ZN(new_n1150));
  AOI21_X1  g725(.A(KEYINPUT62), .B1(new_n1150), .B2(new_n1089), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1147), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1150), .A2(KEYINPUT62), .A3(new_n1089), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1146), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1131), .A2(new_n1142), .A3(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(new_n984), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n770), .B(new_n1105), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n732), .B(G1996), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1157), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(KEYINPUT110), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n801), .B(new_n803), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1161), .B1(new_n1157), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1157), .ZN(new_n1164));
  XNOR2_X1  g739(.A(G290), .B(G1986), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1163), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1155), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1157), .B1(new_n1158), .B2(new_n732), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1168), .B(KEYINPUT127), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1157), .A2(G1996), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1170), .B(KEYINPUT46), .ZN(new_n1171));
  OR3_X1    g746(.A1(new_n1169), .A2(KEYINPUT47), .A3(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(KEYINPUT47), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1157), .A2(G1986), .A3(G290), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n1175), .B(KEYINPUT48), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1174), .B1(new_n1163), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1161), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n799), .A2(new_n803), .A3(new_n800), .ZN(new_n1179));
  OAI22_X1  g754(.A1(new_n1178), .A2(new_n1179), .B1(G2067), .B2(new_n770), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n1180), .A2(new_n1164), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1177), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1167), .A2(new_n1182), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g758(.A1(G229), .A2(new_n460), .A3(new_n673), .A4(G227), .ZN(new_n1185));
  NAND3_X1  g759(.A1(new_n975), .A2(new_n1185), .A3(new_n882), .ZN(G225));
  INV_X1    g760(.A(G225), .ZN(G308));
endmodule


