//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 0 0 0 1 1 1 0 0 0 1 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n789, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n873, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(KEYINPUT93), .A2(G8gat), .ZN(new_n205));
  OAI211_X1 g004(.A(new_n204), .B(new_n205), .C1(G1gat), .C2(new_n202), .ZN(new_n206));
  NOR2_X1   g005(.A1(KEYINPUT93), .A2(G8gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT92), .ZN(new_n210));
  INV_X1    g009(.A(G43gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n210), .B1(new_n211), .B2(G50gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT15), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT14), .ZN(new_n215));
  INV_X1    g014(.A(G29gat), .ZN(new_n216));
  INV_X1    g015(.A(G36gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(G29gat), .A2(G36gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT91), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(KEYINPUT91), .A2(G29gat), .A3(G36gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n214), .A2(new_n220), .A3(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G43gat), .B(G50gat), .ZN(new_n227));
  AOI22_X1  g026(.A1(new_n219), .A2(new_n218), .B1(new_n223), .B2(new_n224), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n226), .B(new_n227), .C1(KEYINPUT15), .C2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n227), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n230), .A3(new_n214), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n209), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G229gat), .A2(G233gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT17), .ZN(new_n235));
  AND3_X1   g034(.A1(new_n229), .A2(new_n235), .A3(new_n231), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n235), .B1(new_n229), .B2(new_n231), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n208), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n233), .A2(new_n234), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT18), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n232), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT94), .B1(new_n208), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n233), .A2(new_n243), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n234), .B(KEYINPUT13), .Z(new_n245));
  NAND3_X1  g044(.A1(new_n209), .A2(KEYINPUT94), .A3(new_n232), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n233), .A2(KEYINPUT18), .A3(new_n234), .A4(new_n238), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n241), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G113gat), .B(G141gat), .ZN(new_n250));
  INV_X1    g049(.A(G197gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT11), .B(G169gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g053(.A(KEYINPUT90), .B(KEYINPUT12), .Z(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n249), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n241), .A2(new_n247), .A3(new_n256), .A4(new_n248), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT27), .B(G183gat), .ZN(new_n263));
  INV_X1    g062(.A(G190gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(KEYINPUT28), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n266));
  AND2_X1   g065(.A1(new_n266), .A2(KEYINPUT27), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n264), .B1(new_n266), .B2(KEYINPUT27), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n265), .B1(new_n269), .B2(KEYINPUT28), .ZN(new_n270));
  INV_X1    g069(.A(G169gat), .ZN(new_n271));
  INV_X1    g070(.A(G176gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT26), .ZN(new_n274));
  NAND2_X1  g073(.A1(G169gat), .A2(G176gat), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n273), .A2(new_n274), .ZN(new_n277));
  INV_X1    g076(.A(G183gat), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n278), .A2(new_n264), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n270), .A2(new_n276), .A3(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n271), .A2(new_n272), .A3(KEYINPUT23), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT23), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n283), .B1(G169gat), .B2(G176gat), .ZN(new_n284));
  AND4_X1   g083(.A1(KEYINPUT25), .A2(new_n282), .A3(new_n284), .A4(new_n275), .ZN(new_n285));
  NAND3_X1  g084(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT24), .B1(new_n286), .B2(KEYINPUT66), .ZN(new_n287));
  NAND2_X1  g086(.A1(KEYINPUT66), .A2(KEYINPUT24), .ZN(new_n288));
  AOI22_X1  g087(.A1(new_n288), .A2(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(G183gat), .A2(G190gat), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n285), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  XOR2_X1   g091(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n293));
  INV_X1    g092(.A(KEYINPUT24), .ZN(new_n294));
  NOR3_X1   g093(.A1(new_n279), .A2(new_n294), .A3(new_n291), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(G183gat), .A3(G190gat), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n282), .A2(new_n284), .A3(new_n296), .A4(new_n275), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n293), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n281), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(G113gat), .B(G120gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT68), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT1), .ZN(new_n303));
  XNOR2_X1  g102(.A(G127gat), .B(G134gat), .ZN(new_n304));
  INV_X1    g103(.A(G113gat), .ZN(new_n305));
  OR3_X1    g104(.A1(new_n305), .A2(KEYINPUT68), .A3(G120gat), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n302), .A2(new_n303), .A3(new_n304), .A4(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n304), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n308), .B1(KEYINPUT1), .B2(new_n301), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n262), .B1(new_n300), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(G227gat), .A2(G233gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n300), .A2(new_n310), .ZN(new_n313));
  INV_X1    g112(.A(new_n310), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n314), .A2(new_n281), .A3(new_n299), .A4(KEYINPUT69), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n311), .A2(new_n312), .A3(new_n313), .A4(new_n315), .ZN(new_n316));
  XOR2_X1   g115(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT71), .ZN(new_n319));
  OR2_X1    g118(.A1(new_n316), .A2(KEYINPUT34), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT71), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n316), .A2(new_n321), .A3(new_n317), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n319), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT72), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT72), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n319), .A2(new_n320), .A3(new_n325), .A4(new_n322), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G15gat), .B(G43gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(G71gat), .B(G99gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n311), .A2(new_n313), .A3(new_n315), .ZN(new_n331));
  INV_X1    g130(.A(new_n312), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT33), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n330), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(KEYINPUT32), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n333), .B(KEYINPUT32), .C1(new_n334), .C2(new_n330), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n327), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n339), .B1(new_n326), .B2(new_n324), .ZN(new_n342));
  OR2_X1    g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT36), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT73), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n324), .A2(new_n345), .A3(new_n326), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n345), .B1(new_n324), .B2(new_n326), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n339), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n342), .A2(new_n344), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n343), .A2(new_n344), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT77), .ZN(new_n351));
  INV_X1    g150(.A(G204gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n251), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(G197gat), .A2(G204gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G211gat), .A2(G218gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n355), .B1(KEYINPUT22), .B2(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(G211gat), .A2(G218gat), .ZN(new_n359));
  OAI21_X1  g158(.A(KEYINPUT74), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n359), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT74), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n361), .A2(new_n362), .A3(new_n356), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n358), .A2(new_n360), .A3(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT75), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n363), .A2(new_n360), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT76), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT22), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n353), .A2(new_n354), .B1(new_n369), .B2(new_n356), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n367), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n368), .B1(new_n367), .B2(new_n370), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n351), .B1(new_n366), .B2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n364), .B(KEYINPUT75), .ZN(new_n376));
  INV_X1    g175(.A(new_n373), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n371), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n376), .A2(new_n378), .A3(KEYINPUT77), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n375), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(G226gat), .ZN(new_n382));
  INV_X1    g181(.A(G233gat), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n300), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n384), .ZN(new_n386));
  AND2_X1   g185(.A1(new_n281), .A2(new_n299), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n386), .B1(new_n387), .B2(KEYINPUT29), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n381), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT78), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n390), .B(new_n386), .C1(new_n387), .C2(KEYINPUT29), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT29), .B1(new_n281), .B2(new_n299), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT78), .B1(new_n392), .B2(new_n384), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n391), .A2(new_n385), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n380), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n389), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(KEYINPUT79), .B(G64gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(G92gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(G8gat), .B(G36gat), .ZN(new_n399));
  XOR2_X1   g198(.A(new_n398), .B(new_n399), .Z(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n389), .A2(new_n395), .A3(new_n400), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n402), .A2(KEYINPUT30), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT30), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n396), .A2(new_n405), .A3(new_n401), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT5), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT85), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT82), .ZN(new_n411));
  AND3_X1   g210(.A1(new_n307), .A2(new_n411), .A3(new_n309), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n411), .B1(new_n307), .B2(new_n309), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G141gat), .B(G148gat), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n415), .A2(KEYINPUT2), .ZN(new_n416));
  XNOR2_X1  g215(.A(G155gat), .B(G162gat), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  XOR2_X1   g217(.A(G141gat), .B(G148gat), .Z(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT80), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT80), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n415), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(G155gat), .A2(G162gat), .ZN(new_n423));
  AOI22_X1  g222(.A1(new_n420), .A2(new_n422), .B1(KEYINPUT2), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n417), .B(KEYINPUT81), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n418), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n410), .B1(new_n414), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n314), .ZN(new_n428));
  INV_X1    g227(.A(new_n418), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n423), .A2(KEYINPUT2), .ZN(new_n430));
  INV_X1    g229(.A(new_n422), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n415), .A2(new_n421), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT81), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n417), .B(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n429), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n436), .B(KEYINPUT85), .C1(new_n413), .C2(new_n412), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n427), .A2(new_n428), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(G225gat), .A2(G233gat), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n409), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT3), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n442), .B(new_n429), .C1(new_n433), .C2(new_n435), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT83), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n426), .A2(KEYINPUT83), .A3(new_n442), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n413), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n307), .A2(new_n411), .A3(new_n309), .ZN(new_n449));
  AOI22_X1  g248(.A1(new_n436), .A2(KEYINPUT3), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n428), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT4), .ZN(new_n453));
  XOR2_X1   g252(.A(KEYINPUT84), .B(KEYINPUT4), .Z(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n440), .B1(new_n428), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n451), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT4), .B1(new_n426), .B2(new_n314), .ZN(new_n459));
  NOR3_X1   g258(.A1(new_n436), .A2(new_n310), .A3(new_n455), .ZN(new_n460));
  AOI211_X1 g259(.A(new_n459), .B(new_n460), .C1(new_n447), .C2(new_n450), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n440), .A2(KEYINPUT5), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(G1gat), .B(G29gat), .ZN(new_n465));
  INV_X1    g264(.A(G85gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  XNOR2_X1  g266(.A(KEYINPUT0), .B(G57gat), .ZN(new_n468));
  XOR2_X1   g267(.A(new_n467), .B(new_n468), .Z(new_n469));
  NAND2_X1  g268(.A1(new_n464), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n427), .A2(new_n428), .A3(new_n439), .A4(new_n437), .ZN(new_n471));
  OAI211_X1 g270(.A(KEYINPUT39), .B(new_n471), .C1(new_n461), .C2(new_n439), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT39), .ZN(new_n473));
  INV_X1    g272(.A(new_n459), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n451), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n473), .B(new_n440), .C1(new_n475), .C2(new_n460), .ZN(new_n476));
  INV_X1    g275(.A(new_n469), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n472), .A2(new_n476), .A3(KEYINPUT40), .A4(new_n477), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n470), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n472), .A2(new_n477), .A3(new_n476), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT40), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n408), .A2(new_n479), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT37), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n389), .A2(new_n484), .A3(new_n395), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n484), .B1(new_n389), .B2(new_n395), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n400), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT38), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n464), .A2(KEYINPUT6), .A3(new_n469), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT87), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n441), .A2(new_n457), .B1(new_n461), .B2(new_n462), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT6), .B1(new_n491), .B2(new_n477), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(new_n470), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n477), .B1(new_n458), .B2(new_n463), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT87), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n494), .A2(new_n495), .A3(KEYINPUT6), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n488), .A2(new_n490), .A3(new_n493), .A4(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n400), .B1(new_n389), .B2(new_n395), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n394), .A2(new_n381), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n380), .A2(new_n385), .A3(new_n388), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(KEYINPUT37), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n501), .B1(new_n396), .B2(KEYINPUT37), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n401), .A2(KEYINPUT38), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n498), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n483), .B1(new_n497), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(G228gat), .A2(G233gat), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT29), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT88), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n377), .A2(new_n509), .A3(new_n371), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(new_n364), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n374), .A2(new_n509), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n508), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n426), .B1(new_n513), .B2(new_n442), .ZN(new_n514));
  AOI21_X1  g313(.A(KEYINPUT29), .B1(new_n445), .B2(new_n446), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n380), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n507), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(G22gat), .ZN(new_n518));
  INV_X1    g317(.A(new_n507), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n376), .A2(new_n378), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT3), .B1(new_n520), .B2(new_n508), .ZN(new_n521));
  OAI221_X1 g320(.A(new_n519), .B1(new_n521), .B2(new_n426), .C1(new_n380), .C2(new_n515), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n517), .A2(new_n518), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT89), .ZN(new_n524));
  XNOR2_X1  g323(.A(G78gat), .B(G106gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(KEYINPUT31), .B(G50gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n525), .B(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n517), .A2(new_n522), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(G22gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(new_n523), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT89), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n530), .A2(new_n533), .A3(new_n523), .A4(new_n527), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n506), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n495), .B1(new_n494), .B2(KEYINPUT6), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT6), .ZN(new_n538));
  NOR4_X1   g337(.A1(new_n491), .A2(KEYINPUT87), .A3(new_n538), .A4(new_n477), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT86), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n494), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT86), .B1(new_n491), .B2(new_n477), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n542), .A2(new_n543), .A3(new_n492), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n408), .B1(new_n540), .B2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n534), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n524), .A2(new_n527), .B1(new_n530), .B2(new_n523), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n350), .B1(new_n536), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n342), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n545), .A2(new_n535), .A3(new_n552), .A4(new_n348), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT35), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n490), .A2(new_n493), .A3(new_n496), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n555), .B(new_n407), .C1(new_n546), .C2(new_n547), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT35), .ZN(new_n558));
  INV_X1    g357(.A(new_n343), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n554), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n261), .B1(new_n551), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT105), .ZN(new_n563));
  XOR2_X1   g362(.A(G190gat), .B(G218gat), .Z(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(G99gat), .ZN(new_n566));
  INV_X1    g365(.A(G106gat), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(G99gat), .A2(G106gat), .ZN(new_n569));
  OAI21_X1  g368(.A(KEYINPUT101), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n568), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT8), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n573), .B1(new_n569), .B2(KEYINPUT101), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(KEYINPUT100), .B(G92gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(new_n466), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT99), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n579), .A2(G85gat), .A3(G92gat), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT7), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n571), .B1(new_n578), .B2(new_n582), .ZN(new_n583));
  AOI22_X1  g382(.A1(new_n572), .A2(new_n574), .B1(new_n576), .B2(new_n466), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n580), .B(KEYINPUT7), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n584), .A2(new_n570), .A3(new_n585), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(KEYINPUT102), .B1(new_n236), .B2(new_n237), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT102), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n589), .B1(new_n236), .B2(new_n237), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n587), .A2(new_n232), .ZN(new_n591));
  AOI22_X1  g390(.A1(new_n587), .A2(new_n588), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G232gat), .A2(G233gat), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n593), .B(KEYINPUT97), .Z(new_n594));
  INV_X1    g393(.A(KEYINPUT41), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n565), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT103), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n588), .A2(new_n587), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n586), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n242), .B(new_n600), .C1(KEYINPUT102), .C2(KEYINPUT17), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n596), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n602), .A2(new_n603), .A3(new_n564), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n597), .A2(new_n598), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n594), .A2(new_n595), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT98), .ZN(new_n607));
  XNOR2_X1  g406(.A(G134gat), .B(G162gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n602), .A2(KEYINPUT103), .A3(new_n603), .A4(new_n564), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n605), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT104), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n605), .A2(KEYINPUT104), .A3(new_n610), .A4(new_n609), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT95), .ZN(new_n616));
  XNOR2_X1  g415(.A(G57gat), .B(G64gat), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(G71gat), .B(G78gat), .Z(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT21), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n278), .B1(new_n208), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n208), .A2(new_n278), .A3(new_n622), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n624), .A2(G231gat), .A3(G233gat), .A4(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G231gat), .A2(G233gat), .ZN(new_n627));
  INV_X1    g426(.A(new_n625), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n627), .B1(new_n628), .B2(new_n623), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n621), .A2(KEYINPUT21), .ZN(new_n631));
  INV_X1    g430(.A(G211gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT96), .ZN(new_n636));
  XOR2_X1   g435(.A(G127gat), .B(G155gat), .Z(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n633), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n626), .A2(new_n639), .A3(new_n629), .ZN(new_n640));
  AND3_X1   g439(.A1(new_n634), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n638), .B1(new_n634), .B2(new_n640), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n609), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n597), .A2(new_n644), .A3(new_n604), .ZN(new_n645));
  AND4_X1   g444(.A1(new_n563), .A2(new_n615), .A3(new_n643), .A4(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n645), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(new_n613), .B2(new_n614), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n563), .B1(new_n648), .B2(new_n643), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n600), .A2(new_n621), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT10), .ZN(new_n653));
  OR2_X1    g452(.A1(new_n619), .A2(new_n620), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n619), .A2(new_n620), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n583), .A2(new_n654), .A3(new_n586), .A4(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n652), .A2(new_n653), .A3(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n600), .A2(KEYINPUT10), .A3(new_n621), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(G230gat), .A2(G233gat), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n652), .A2(new_n656), .ZN(new_n662));
  INV_X1    g461(.A(new_n660), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(G120gat), .B(G148gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(G176gat), .B(G204gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n665), .A2(new_n668), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n651), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n562), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n544), .A2(new_n496), .A3(new_n490), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g477(.A1(new_n673), .A2(new_n407), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT16), .B(G8gat), .Z(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT42), .ZN(new_n682));
  INV_X1    g481(.A(G8gat), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n682), .B1(new_n683), .B2(new_n679), .ZN(G1325gat));
  INV_X1    g483(.A(G15gat), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n348), .A2(new_n349), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n344), .B1(new_n341), .B2(new_n342), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT106), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n686), .A2(KEYINPUT106), .A3(new_n687), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n673), .A2(new_n685), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n674), .A2(new_n559), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n693), .B1(new_n685), .B2(new_n694), .ZN(G1326gat));
  NOR2_X1   g494(.A1(new_n673), .A2(new_n535), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT107), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT43), .B(G22gat), .Z(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1327gat));
  INV_X1    g498(.A(new_n648), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n556), .A2(KEYINPUT35), .ZN(new_n701));
  AOI22_X1  g500(.A1(new_n701), .A2(new_n559), .B1(new_n553), .B2(KEYINPUT35), .ZN(new_n702));
  OAI211_X1 g501(.A(KEYINPUT44), .B(new_n700), .C1(new_n702), .C2(new_n550), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n671), .B(KEYINPUT109), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n705), .A2(new_n261), .A3(new_n643), .ZN(new_n706));
  INV_X1    g505(.A(new_n691), .ZN(new_n707));
  AOI21_X1  g506(.A(KEYINPUT106), .B1(new_n686), .B2(new_n687), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n540), .A2(new_n493), .A3(new_n488), .A4(new_n504), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n548), .B1(new_n709), .B2(new_n483), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n545), .A2(new_n548), .ZN(new_n711));
  OAI22_X1  g510(.A1(new_n707), .A2(new_n708), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n648), .B1(new_n712), .B2(new_n561), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n703), .B(new_n706), .C1(new_n713), .C2(KEYINPUT44), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT110), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n536), .A2(new_n549), .ZN(new_n718));
  AOI22_X1  g517(.A1(new_n692), .A2(new_n718), .B1(new_n554), .B2(new_n560), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n717), .B1(new_n719), .B2(new_n648), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n720), .A2(KEYINPUT110), .A3(new_n703), .A4(new_n706), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n716), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(G29gat), .B1(new_n723), .B2(new_n675), .ZN(new_n724));
  INV_X1    g523(.A(new_n643), .ZN(new_n725));
  INV_X1    g524(.A(new_n671), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n700), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT108), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OR2_X1    g528(.A1(new_n727), .A2(new_n728), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n562), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n731), .A2(new_n216), .A3(new_n676), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT45), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n724), .A2(new_n733), .ZN(G1328gat));
  NOR2_X1   g533(.A1(new_n407), .A2(G36gat), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n562), .A2(new_n729), .A3(new_n730), .A4(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT46), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n407), .B1(new_n716), .B2(new_n721), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n739), .B2(new_n217), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT111), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n738), .B(KEYINPUT111), .C1(new_n739), .C2(new_n217), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(G1329gat));
  INV_X1    g543(.A(KEYINPUT47), .ZN(new_n745));
  INV_X1    g544(.A(new_n692), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n211), .B1(new_n722), .B2(new_n746), .ZN(new_n747));
  AND3_X1   g546(.A1(new_n731), .A2(new_n211), .A3(new_n559), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n745), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n714), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n211), .B1(new_n750), .B2(new_n746), .ZN(new_n751));
  OR3_X1    g550(.A1(new_n751), .A2(new_n748), .A3(new_n745), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n749), .A2(new_n752), .ZN(G1330gat));
  INV_X1    g552(.A(KEYINPUT48), .ZN(new_n754));
  INV_X1    g553(.A(G50gat), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n731), .A2(KEYINPUT112), .A3(new_n755), .A4(new_n548), .ZN(new_n756));
  OAI21_X1  g555(.A(G50gat), .B1(new_n714), .B2(new_n535), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n754), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI211_X1 g557(.A(new_n754), .B(G50gat), .C1(new_n723), .C2(new_n535), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n731), .A2(new_n548), .ZN(new_n760));
  AOI22_X1  g559(.A1(new_n760), .A2(new_n755), .B1(KEYINPUT112), .B2(KEYINPUT48), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n758), .B1(new_n759), .B2(new_n761), .ZN(G1331gat));
  NOR2_X1   g561(.A1(new_n719), .A2(new_n651), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n704), .A2(new_n260), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n676), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g567(.A1(new_n765), .A2(new_n407), .ZN(new_n769));
  NOR2_X1   g568(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n770));
  AND2_X1   g569(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n772), .B1(new_n769), .B2(new_n770), .ZN(G1333gat));
  NAND4_X1  g572(.A1(new_n763), .A2(G71gat), .A3(new_n746), .A4(new_n764), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT113), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n774), .B(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT115), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n343), .B(KEYINPUT114), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n765), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(G71gat), .ZN(new_n780));
  INV_X1    g579(.A(new_n778), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n763), .A2(KEYINPUT115), .A3(new_n764), .A4(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n779), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n776), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT50), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT50), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n776), .A2(new_n786), .A3(new_n783), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(G1334gat));
  NAND2_X1  g587(.A1(new_n766), .A2(new_n548), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g589(.A1(new_n643), .A2(new_n260), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n720), .A2(new_n671), .A3(new_n703), .A4(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n793));
  OR3_X1    g592(.A1(new_n792), .A2(new_n793), .A3(new_n675), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n793), .B1(new_n792), .B2(new_n675), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n794), .A2(G85gat), .A3(new_n795), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n713), .A2(KEYINPUT51), .A3(new_n791), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT51), .B1(new_n713), .B2(new_n791), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n671), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n676), .A2(new_n466), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n796), .B1(new_n799), .B2(new_n800), .ZN(G1336gat));
  INV_X1    g600(.A(new_n576), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n802), .B1(new_n792), .B2(new_n407), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT117), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n407), .A2(G92gat), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n705), .B(new_n806), .C1(new_n797), .C2(new_n798), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n803), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n805), .A2(new_n808), .A3(KEYINPUT52), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n803), .B(new_n807), .C1(new_n804), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(G1337gat));
  OAI21_X1  g611(.A(G99gat), .B1(new_n792), .B2(new_n692), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n559), .A2(new_n566), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n799), .B2(new_n814), .ZN(G1338gat));
  OAI21_X1  g614(.A(G106gat), .B1(new_n792), .B2(new_n535), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT118), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n535), .A2(G106gat), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n705), .B(new_n819), .C1(new_n797), .C2(new_n798), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n818), .A2(new_n821), .A3(KEYINPUT53), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT53), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n816), .B(new_n820), .C1(new_n817), .C2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(G1339gat));
  NAND4_X1  g624(.A1(new_n650), .A2(KEYINPUT119), .A3(new_n261), .A4(new_n726), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n615), .A2(new_n643), .A3(new_n645), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT105), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n648), .A2(new_n563), .A3(new_n643), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n828), .A2(new_n261), .A3(new_n829), .A4(new_n726), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT119), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n245), .B1(new_n244), .B2(new_n246), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n234), .B1(new_n233), .B2(new_n238), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n254), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n259), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n671), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT122), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n657), .A2(new_n658), .A3(new_n663), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(KEYINPUT120), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n657), .A2(new_n842), .A3(new_n658), .A4(new_n663), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n841), .A2(new_n661), .A3(KEYINPUT54), .A4(new_n843), .ZN(new_n844));
  XNOR2_X1  g643(.A(KEYINPUT121), .B(KEYINPUT54), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n659), .A2(new_n660), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n844), .A2(new_n846), .A3(new_n668), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT55), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n844), .A2(new_n846), .A3(KEYINPUT55), .A4(new_n668), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n849), .A2(new_n260), .A3(new_n669), .A4(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT122), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n852), .A3(new_n671), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n839), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n854), .A2(new_n648), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n849), .A2(new_n669), .A3(new_n850), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n648), .A2(new_n856), .A3(new_n836), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n725), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n826), .A2(new_n832), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n676), .ZN(new_n860));
  INV_X1    g659(.A(new_n348), .ZN(new_n861));
  NOR4_X1   g660(.A1(new_n860), .A2(new_n342), .A3(new_n861), .A4(new_n548), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n407), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n864), .A2(new_n305), .A3(new_n260), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n675), .A2(new_n408), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n859), .A2(new_n559), .A3(new_n535), .A4(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(G113gat), .B1(new_n867), .B2(new_n261), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n865), .A2(new_n868), .ZN(G1340gat));
  OAI21_X1  g668(.A(G120gat), .B1(new_n867), .B2(new_n704), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n863), .A2(G120gat), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n870), .B1(new_n871), .B2(new_n726), .ZN(G1341gat));
  INV_X1    g671(.A(G127gat), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n867), .A2(new_n873), .A3(new_n725), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n864), .A2(new_n643), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n874), .B1(new_n875), .B2(new_n873), .ZN(G1342gat));
  OR2_X1    g675(.A1(new_n648), .A2(G134gat), .ZN(new_n877));
  OR3_X1    g676(.A1(new_n863), .A2(KEYINPUT56), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(G134gat), .B1(new_n867), .B2(new_n648), .ZN(new_n879));
  OAI21_X1  g678(.A(KEYINPUT56), .B1(new_n863), .B2(new_n877), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(G1343gat));
  INV_X1    g680(.A(KEYINPUT124), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT58), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n860), .A2(new_n535), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n884), .A2(new_n407), .A3(new_n260), .A4(new_n692), .ZN(new_n885));
  INV_X1    g684(.A(G141gat), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n859), .A2(new_n548), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT57), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n692), .A2(new_n866), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n856), .A2(KEYINPUT123), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT123), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n849), .A2(new_n894), .A3(new_n669), .A4(new_n850), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n893), .A2(new_n260), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n700), .B1(new_n896), .B2(new_n838), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n725), .B1(new_n897), .B2(new_n857), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n826), .A2(new_n832), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n548), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n892), .B1(new_n900), .B2(KEYINPUT57), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n891), .A2(new_n901), .A3(G141gat), .A4(new_n260), .ZN(new_n902));
  AOI211_X1 g701(.A(new_n882), .B(new_n883), .C1(new_n887), .C2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(KEYINPUT124), .A2(KEYINPUT58), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n882), .A2(new_n883), .ZN(new_n905));
  AND4_X1   g704(.A1(new_n904), .A2(new_n887), .A3(new_n905), .A4(new_n902), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n903), .A2(new_n906), .ZN(G1344gat));
  NOR4_X1   g706(.A1(new_n860), .A2(new_n535), .A3(new_n408), .A4(new_n746), .ZN(new_n908));
  INV_X1    g707(.A(G148gat), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(new_n909), .A3(new_n671), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n891), .A2(new_n901), .ZN(new_n911));
  AOI211_X1 g710(.A(KEYINPUT59), .B(new_n909), .C1(new_n911), .C2(new_n671), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT59), .ZN(new_n913));
  AOI211_X1 g712(.A(KEYINPUT57), .B(new_n535), .C1(new_n898), .C2(new_n830), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n914), .B1(new_n888), .B2(KEYINPUT57), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n915), .A2(new_n671), .A3(new_n692), .A4(new_n866), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n913), .B1(new_n916), .B2(G148gat), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n910), .B1(new_n912), .B2(new_n917), .ZN(G1345gat));
  AOI21_X1  g717(.A(G155gat), .B1(new_n908), .B2(new_n643), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n911), .A2(G155gat), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n919), .B1(new_n920), .B2(new_n643), .ZN(G1346gat));
  INV_X1    g720(.A(G162gat), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n908), .A2(new_n922), .A3(new_n700), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n911), .A2(new_n700), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n923), .B1(new_n924), .B2(new_n922), .ZN(G1347gat));
  NAND2_X1  g724(.A1(new_n675), .A2(new_n408), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n859), .A2(new_n535), .A3(new_n927), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n861), .A2(new_n342), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n931), .A2(new_n271), .A3(new_n260), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n928), .A2(new_n781), .ZN(new_n933));
  OAI21_X1  g732(.A(G169gat), .B1(new_n933), .B2(new_n261), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(G1348gat));
  NOR3_X1   g734(.A1(new_n933), .A2(new_n272), .A3(new_n704), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n931), .A2(new_n671), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n936), .B1(new_n272), .B2(new_n937), .ZN(G1349gat));
  NAND3_X1  g737(.A1(new_n931), .A2(new_n263), .A3(new_n643), .ZN(new_n939));
  OAI21_X1  g738(.A(G183gat), .B1(new_n933), .B2(new_n725), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g741(.A(G190gat), .B1(new_n933), .B2(new_n648), .ZN(new_n943));
  XOR2_X1   g742(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n944));
  XNOR2_X1  g743(.A(new_n943), .B(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n931), .A2(new_n264), .A3(new_n700), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1351gat));
  NOR2_X1   g746(.A1(new_n746), .A2(new_n926), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n889), .A2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n950), .A2(new_n251), .A3(new_n260), .ZN(new_n951));
  OR2_X1    g750(.A1(new_n915), .A2(KEYINPUT126), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n915), .A2(KEYINPUT126), .ZN(new_n953));
  AND4_X1   g752(.A1(new_n260), .A2(new_n952), .A3(new_n948), .A4(new_n953), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n951), .B1(new_n954), .B2(new_n251), .ZN(G1352gat));
  NOR3_X1   g754(.A1(new_n949), .A2(G204gat), .A3(new_n726), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n956), .B(KEYINPUT62), .ZN(new_n957));
  AND4_X1   g756(.A1(new_n705), .A2(new_n952), .A3(new_n948), .A4(new_n953), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n957), .B1(new_n352), .B2(new_n958), .ZN(G1353gat));
  NAND3_X1  g758(.A1(new_n950), .A2(new_n632), .A3(new_n643), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT63), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n746), .A2(new_n725), .A3(new_n926), .ZN(new_n962));
  AOI211_X1 g761(.A(new_n961), .B(new_n632), .C1(new_n915), .C2(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n888), .A2(KEYINPUT57), .ZN(new_n964));
  INV_X1    g763(.A(new_n914), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n964), .A2(new_n965), .A3(new_n962), .ZN(new_n966));
  AOI21_X1  g765(.A(KEYINPUT63), .B1(new_n966), .B2(G211gat), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n960), .B1(new_n963), .B2(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI211_X1 g769(.A(KEYINPUT127), .B(new_n960), .C1(new_n963), .C2(new_n967), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(G1354gat));
  INV_X1    g771(.A(G218gat), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n950), .A2(new_n973), .A3(new_n700), .ZN(new_n974));
  AND4_X1   g773(.A1(new_n700), .A2(new_n952), .A3(new_n948), .A4(new_n953), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n974), .B1(new_n975), .B2(new_n973), .ZN(G1355gat));
endmodule


