//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 0 1 0 0 0 0 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n762, new_n763, new_n764,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n832, new_n833, new_n834, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953;
  XNOR2_X1  g000(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g002(.A(G155gat), .B(G162gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT2), .ZN(new_n205));
  XOR2_X1   g004(.A(KEYINPUT80), .B(G155gat), .Z(new_n206));
  AOI21_X1  g005(.A(new_n205), .B1(new_n206), .B2(G162gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT79), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n204), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NOR2_X1   g008(.A1(KEYINPUT78), .A2(KEYINPUT2), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n204), .A2(new_n210), .ZN(new_n211));
  XOR2_X1   g010(.A(G141gat), .B(G148gat), .Z(new_n212));
  OR2_X1    g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NOR3_X1   g012(.A1(new_n204), .A2(new_n208), .A3(KEYINPUT2), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n214), .A2(KEYINPUT78), .A3(new_n212), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n209), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n217));
  AOI21_X1  g016(.A(KEYINPUT29), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(G197gat), .B(G204gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT22), .ZN(new_n220));
  INV_X1    g019(.A(G211gat), .ZN(new_n221));
  INV_X1    g020(.A(G218gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n219), .A2(new_n223), .ZN(new_n224));
  XOR2_X1   g023(.A(G211gat), .B(G218gat), .Z(new_n225));
  XOR2_X1   g024(.A(new_n224), .B(new_n225), .Z(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT74), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n224), .B(new_n225), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT74), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n218), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT29), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n228), .A2(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n216), .B1(new_n217), .B2(new_n234), .ZN(new_n235));
  OAI211_X1 g034(.A(G228gat), .B(G233gat), .C1(new_n232), .C2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n216), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n217), .B1(new_n234), .B2(KEYINPUT84), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT84), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n239), .B1(new_n228), .B2(new_n233), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n237), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G228gat), .A2(G233gat), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n241), .B(new_n242), .C1(new_n231), .C2(new_n218), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n236), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT85), .B(G50gat), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G78gat), .B(G106gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(G22gat), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n236), .A2(new_n243), .A3(new_n245), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n247), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n250), .B1(new_n247), .B2(new_n251), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n203), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n247), .A2(new_n251), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(new_n249), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n247), .A2(new_n250), .A3(new_n251), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n256), .A2(new_n257), .A3(new_n202), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(G226gat), .A2(G233gat), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(G183gat), .A2(G190gat), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT24), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n265));
  AND2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(G183gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT66), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT66), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(G183gat), .ZN(new_n270));
  INV_X1    g069(.A(G190gat), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n268), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  AND2_X1   g071(.A1(new_n266), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g072(.A1(G169gat), .A2(G176gat), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(G169gat), .A2(G176gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT23), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n274), .A2(KEYINPUT23), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(KEYINPUT25), .B1(new_n273), .B2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT65), .B(G169gat), .ZN(new_n282));
  INV_X1    g081(.A(G176gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(KEYINPUT23), .A3(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n267), .A2(new_n271), .A3(KEYINPUT64), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT64), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n286), .B1(G183gat), .B2(G190gat), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n264), .A2(new_n285), .A3(new_n287), .A4(new_n265), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT25), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n284), .A2(new_n288), .A3(new_n289), .A4(new_n278), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT28), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT27), .B(G183gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT68), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n267), .A2(KEYINPUT27), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT27), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n296), .A2(G183gat), .ZN(new_n297));
  OAI21_X1  g096(.A(KEYINPUT68), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n291), .B1(new_n299), .B2(new_n271), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n275), .A2(KEYINPUT26), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT26), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n274), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n301), .A2(new_n276), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n295), .A2(KEYINPUT67), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n305), .A2(new_n291), .A3(new_n271), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n269), .A2(KEYINPUT67), .A3(G183gat), .ZN(new_n307));
  AND3_X1   g106(.A1(new_n307), .A2(KEYINPUT27), .A3(new_n268), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n304), .B(new_n262), .C1(new_n306), .C2(new_n308), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n281), .B(new_n290), .C1(new_n300), .C2(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n261), .B1(new_n310), .B2(new_n233), .ZN(new_n311));
  OR2_X1    g110(.A1(new_n300), .A2(new_n309), .ZN(new_n312));
  INV_X1    g111(.A(new_n280), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n266), .A2(new_n272), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n289), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n290), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n260), .B1(new_n312), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(KEYINPUT75), .B1(new_n311), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT75), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT29), .B1(new_n312), .B2(new_n317), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n320), .B1(new_n321), .B2(new_n261), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n319), .A2(new_n231), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT76), .ZN(new_n324));
  INV_X1    g123(.A(new_n231), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n325), .B1(new_n311), .B2(new_n318), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT76), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n319), .A2(new_n327), .A3(new_n322), .A4(new_n231), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n324), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G8gat), .B(G36gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(G92gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n331), .B(KEYINPUT77), .ZN(new_n332));
  INV_X1    g131(.A(G64gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n332), .B(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  OR3_X1    g134(.A1(new_n329), .A2(KEYINPUT30), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n329), .A2(new_n335), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n324), .A2(new_n326), .A3(new_n334), .A4(new_n328), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(KEYINPUT30), .A3(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(KEYINPUT0), .B(G57gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n340), .B(G85gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(G1gat), .B(G29gat), .ZN(new_n342));
  XOR2_X1   g141(.A(new_n341), .B(new_n342), .Z(new_n343));
  XNOR2_X1  g142(.A(G127gat), .B(G134gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(G113gat), .B(G120gat), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n344), .B1(new_n345), .B2(KEYINPUT69), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(KEYINPUT1), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n346), .A2(new_n347), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n216), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT4), .ZN(new_n353));
  NAND2_X1  g152(.A1(G225gat), .A2(G233gat), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n352), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n216), .A2(new_n217), .ZN(new_n357));
  INV_X1    g156(.A(new_n351), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n209), .A2(KEYINPUT3), .A3(new_n213), .A4(new_n215), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n216), .A2(KEYINPUT4), .A3(new_n351), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n356), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n237), .A2(KEYINPUT81), .A3(new_n358), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT81), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n364), .B1(new_n216), .B2(new_n351), .ZN(new_n365));
  AOI22_X1  g164(.A1(new_n363), .A2(new_n365), .B1(new_n351), .B2(new_n216), .ZN(new_n366));
  OAI211_X1 g165(.A(KEYINPUT5), .B(new_n362), .C1(new_n366), .C2(new_n354), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT82), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n216), .A2(new_n368), .A3(new_n351), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n368), .B1(new_n216), .B2(new_n351), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n353), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n371), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n373), .A2(KEYINPUT4), .A3(new_n369), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n355), .A2(KEYINPUT5), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n372), .A2(new_n374), .A3(new_n360), .A4(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n343), .B1(new_n367), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT88), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n372), .A2(new_n374), .A3(new_n360), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT39), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(new_n381), .A3(new_n355), .ZN(new_n382));
  AND2_X1   g181(.A1(new_n382), .A2(new_n343), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n363), .A2(new_n365), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n384), .A2(new_n354), .A3(new_n352), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT39), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT86), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n380), .A2(new_n355), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT86), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n385), .A2(new_n389), .A3(KEYINPUT39), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n387), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n383), .A2(new_n391), .A3(KEYINPUT40), .ZN(new_n392));
  AND4_X1   g191(.A1(new_n336), .A2(new_n339), .A3(new_n379), .A4(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT40), .B1(new_n383), .B2(new_n391), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n394), .A2(KEYINPUT87), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT87), .ZN(new_n396));
  AOI211_X1 g195(.A(new_n396), .B(KEYINPUT40), .C1(new_n383), .C2(new_n391), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n259), .B1(new_n393), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT37), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n324), .A2(new_n326), .A3(new_n400), .A4(new_n328), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT38), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n319), .A2(new_n325), .A3(new_n322), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n231), .B1(new_n311), .B2(new_n318), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n403), .A2(KEYINPUT37), .A3(new_n404), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n401), .A2(new_n402), .A3(new_n335), .A4(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT89), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  AND2_X1   g207(.A1(new_n329), .A2(KEYINPUT37), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n401), .A2(new_n335), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT38), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT90), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n329), .A2(KEYINPUT37), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n413), .A2(new_n335), .A3(new_n401), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT90), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n414), .A2(new_n415), .A3(KEYINPUT38), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n408), .A2(new_n412), .A3(new_n338), .A4(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n377), .A2(KEYINPUT6), .ZN(new_n418));
  INV_X1    g217(.A(new_n379), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT6), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n367), .A2(new_n376), .ZN(new_n421));
  INV_X1    g220(.A(new_n343), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n418), .B1(new_n419), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n399), .B1(new_n417), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n310), .A2(KEYINPUT70), .A3(new_n351), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT70), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n349), .A2(new_n427), .A3(new_n350), .ZN(new_n428));
  INV_X1    g227(.A(new_n350), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT70), .B1(new_n429), .B2(new_n348), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n312), .A2(new_n317), .A3(new_n428), .A4(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(G227gat), .A2(G233gat), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT34), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n434), .A2(KEYINPUT71), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n432), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n433), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n437), .B1(new_n426), .B2(new_n431), .ZN(new_n438));
  XOR2_X1   g237(.A(KEYINPUT71), .B(KEYINPUT34), .Z(new_n439));
  OAI21_X1  g238(.A(new_n436), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n426), .A2(new_n431), .A3(new_n437), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT33), .ZN(new_n442));
  XNOR2_X1  g241(.A(G15gat), .B(G43gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(G71gat), .B(G99gat), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n443), .B(new_n444), .Z(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n441), .B(KEYINPUT32), .C1(new_n442), .C2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n441), .A2(KEYINPUT32), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n441), .A2(new_n442), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n449), .A3(new_n445), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n440), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n450), .A2(new_n440), .A3(new_n447), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT72), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT73), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT72), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n450), .A2(new_n440), .A3(new_n456), .A4(new_n447), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n454), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n455), .B1(new_n454), .B2(new_n457), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n452), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT36), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n451), .B1(new_n454), .B2(new_n457), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT36), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n339), .A2(new_n336), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n418), .B1(new_n423), .B2(new_n377), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n462), .A2(new_n464), .B1(new_n467), .B2(new_n259), .ZN(new_n468));
  AND2_X1   g267(.A1(new_n339), .A2(new_n336), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n460), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT35), .ZN(new_n471));
  AND2_X1   g270(.A1(new_n254), .A2(new_n258), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n470), .A2(new_n471), .A3(new_n472), .A4(new_n424), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n254), .A2(new_n258), .A3(new_n463), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT35), .B1(new_n475), .B2(new_n467), .ZN(new_n476));
  AOI22_X1  g275(.A1(new_n425), .A2(new_n468), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G127gat), .B(G155gat), .ZN(new_n478));
  XOR2_X1   g277(.A(new_n478), .B(KEYINPUT20), .Z(new_n479));
  XNOR2_X1  g278(.A(G15gat), .B(G22gat), .ZN(new_n480));
  INV_X1    g279(.A(G1gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT16), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT95), .ZN(new_n484));
  OR2_X1    g283(.A1(G15gat), .A2(G22gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(G15gat), .A2(G22gat), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n485), .A2(new_n481), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n484), .A2(new_n488), .A3(G8gat), .ZN(new_n489));
  INV_X1    g288(.A(G8gat), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n483), .B(new_n487), .C1(KEYINPUT95), .C2(new_n490), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(G71gat), .A2(G78gat), .ZN(new_n493));
  NOR2_X1   g292(.A1(G71gat), .A2(G78gat), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n493), .B1(new_n494), .B2(KEYINPUT99), .ZN(new_n495));
  OR2_X1    g294(.A1(new_n493), .A2(KEYINPUT99), .ZN(new_n496));
  XNOR2_X1  g295(.A(G57gat), .B(G64gat), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n495), .B(new_n496), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT101), .ZN(new_n500));
  NAND3_X1  g299(.A1(KEYINPUT100), .A2(G57gat), .A3(G64gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(KEYINPUT100), .A2(G57gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(new_n333), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT9), .ZN(new_n504));
  NOR3_X1   g303(.A1(new_n504), .A2(G71gat), .A3(G78gat), .ZN(new_n505));
  INV_X1    g304(.A(new_n493), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n501), .B(new_n503), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  AND3_X1   g306(.A1(new_n499), .A2(new_n500), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n500), .B1(new_n499), .B2(new_n507), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT21), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n492), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OR2_X1    g311(.A1(new_n512), .A2(G183gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(G183gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(G231gat), .A2(G233gat), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n513), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n516), .B1(new_n513), .B2(new_n514), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n479), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n513), .A2(new_n514), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(new_n515), .ZN(new_n522));
  INV_X1    g321(.A(new_n479), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(new_n517), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n511), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT102), .B(KEYINPUT19), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(G211gat), .ZN(new_n528));
  XOR2_X1   g327(.A(new_n526), .B(new_n528), .Z(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n525), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n520), .A2(new_n524), .A3(new_n529), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT14), .ZN(new_n535));
  OR3_X1    g334(.A1(new_n535), .A2(G29gat), .A3(G36gat), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n535), .B1(G29gat), .B2(G36gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(KEYINPUT92), .B(G29gat), .ZN(new_n538));
  INV_X1    g337(.A(G36gat), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n536), .B(new_n537), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(G43gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(G50gat), .ZN(new_n542));
  INV_X1    g341(.A(G50gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(G43gat), .ZN(new_n544));
  AND3_X1   g343(.A1(new_n542), .A2(new_n544), .A3(KEYINPUT15), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n540), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(KEYINPUT93), .B1(new_n541), .B2(G50gat), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT94), .B1(new_n543), .B2(G43gat), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT93), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n550), .A2(new_n543), .A3(G43gat), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT94), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n552), .A2(new_n541), .A3(G50gat), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n548), .A2(new_n549), .A3(new_n551), .A4(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT15), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n545), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n547), .B1(new_n556), .B2(new_n540), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT17), .ZN(new_n558));
  NAND2_X1  g357(.A1(G99gat), .A2(G106gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g359(.A1(G85gat), .A2(G92gat), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT7), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(G85gat), .ZN(new_n564));
  INV_X1    g363(.A(G92gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n560), .A2(new_n563), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G99gat), .B(G106gat), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  AOI22_X1  g370(.A1(KEYINPUT8), .A2(new_n559), .B1(new_n564), .B2(new_n565), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n572), .A2(new_n569), .A3(new_n563), .A4(new_n567), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT17), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n547), .B(new_n575), .C1(new_n556), .C2(new_n540), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n558), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n556), .A2(new_n540), .ZN(new_n579));
  INV_X1    g378(.A(new_n574), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n579), .A2(new_n580), .A3(new_n547), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n577), .A2(new_n578), .A3(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G134gat), .B(G162gat), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n583), .B(KEYINPUT103), .Z(new_n584));
  OR2_X1    g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G190gat), .B(G218gat), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n582), .A2(new_n584), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n585), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n588), .B1(new_n585), .B2(new_n589), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR3_X1   g391(.A1(new_n477), .A2(new_n534), .A3(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n558), .A2(new_n492), .A3(new_n576), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n489), .A2(new_n491), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n595), .A3(new_n547), .ZN(new_n596));
  AND2_X1   g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT98), .ZN(new_n598));
  NAND2_X1  g397(.A1(G229gat), .A2(G233gat), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n599), .B(KEYINPUT96), .Z(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n597), .A2(new_n598), .A3(KEYINPUT18), .A4(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n594), .A2(new_n596), .A3(new_n601), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT18), .ZN(new_n604));
  OAI21_X1  g403(.A(KEYINPUT98), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n492), .A2(new_n557), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(new_n596), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n600), .B(KEYINPUT13), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n602), .A2(KEYINPUT97), .A3(new_n605), .A4(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n603), .A2(new_n604), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n602), .A2(new_n609), .A3(new_n605), .A4(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G113gat), .B(G141gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(G169gat), .B(G197gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(KEYINPUT91), .B(KEYINPUT11), .Z(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT12), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  AND3_X1   g418(.A1(new_n610), .A2(new_n612), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n612), .B1(new_n610), .B2(new_n619), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G120gat), .B(G148gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(new_n283), .ZN(new_n624));
  INV_X1    g423(.A(G204gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(G230gat), .A2(G233gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT104), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n499), .A2(new_n507), .ZN(new_n631));
  AND3_X1   g430(.A1(new_n631), .A2(new_n573), .A3(new_n571), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(KEYINPUT101), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n499), .A2(new_n500), .A3(new_n507), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n632), .B1(new_n635), .B2(new_n574), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT105), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n580), .B(KEYINPUT10), .C1(new_n508), .C2(new_n509), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n639), .B1(new_n636), .B2(KEYINPUT10), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n638), .B1(new_n640), .B2(new_n630), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n574), .B1(new_n508), .B2(new_n509), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n580), .A2(new_n631), .ZN(new_n643));
  AOI21_X1  g442(.A(KEYINPUT10), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n639), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n638), .B(new_n630), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  OAI221_X1 g446(.A(new_n627), .B1(new_n630), .B2(new_n637), .C1(new_n641), .C2(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n644), .A2(new_n645), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n649), .A2(new_n629), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n637), .A2(new_n630), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n626), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n622), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n593), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n655), .A2(new_n466), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(new_n481), .ZN(G1324gat));
  NOR2_X1   g456(.A1(new_n655), .A2(new_n465), .ZN(new_n658));
  NAND2_X1  g457(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n659));
  OR2_X1    g458(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT42), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n663), .B(new_n664), .C1(new_n490), .C2(new_n658), .ZN(G1325gat));
  INV_X1    g464(.A(G15gat), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n454), .A2(new_n457), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(KEYINPUT73), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n454), .A2(new_n455), .A3(new_n457), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n451), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n464), .B1(new_n670), .B2(KEYINPUT36), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n655), .A2(new_n666), .A3(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n593), .A2(new_n670), .A3(new_n654), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n672), .B1(new_n666), .B2(new_n673), .ZN(G1326gat));
  NOR2_X1   g473(.A1(new_n655), .A2(new_n472), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT43), .B(G22gat), .Z(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1327gat));
  INV_X1    g476(.A(new_n592), .ZN(new_n678));
  INV_X1    g477(.A(new_n653), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n602), .A2(new_n609), .A3(new_n605), .ZN(new_n680));
  OAI211_X1 g479(.A(new_n680), .B(new_n611), .C1(KEYINPUT97), .C2(new_n618), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n610), .A2(new_n612), .A3(new_n619), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n534), .A2(new_n679), .A3(new_n683), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n477), .A2(new_n678), .A3(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n466), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n685), .A2(new_n686), .A3(new_n538), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT45), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n689), .B1(new_n477), .B2(new_n678), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n467), .A2(new_n259), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n671), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n416), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n415), .B1(new_n414), .B2(KEYINPUT38), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n424), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n695), .A2(new_n696), .A3(new_n338), .A4(new_n408), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n692), .B1(new_n697), .B2(new_n399), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n469), .A2(new_n686), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n471), .B1(new_n699), .B2(new_n474), .ZN(new_n700));
  AND4_X1   g499(.A1(new_n471), .A2(new_n424), .A3(new_n670), .A4(new_n465), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n700), .B1(new_n472), .B2(new_n701), .ZN(new_n702));
  OAI211_X1 g501(.A(KEYINPUT44), .B(new_n592), .C1(new_n698), .C2(new_n702), .ZN(new_n703));
  XOR2_X1   g502(.A(new_n653), .B(KEYINPUT106), .Z(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n705), .A2(new_n533), .A3(new_n622), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n690), .A2(new_n703), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(KEYINPUT107), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n690), .A2(new_n703), .A3(new_n709), .A4(new_n706), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n466), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n688), .B1(new_n711), .B2(new_n538), .ZN(G1328gat));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n708), .A2(new_n710), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n539), .B1(new_n714), .B2(new_n469), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n685), .A2(new_n539), .A3(new_n469), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT46), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n713), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT46), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n716), .B(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n465), .B1(new_n708), .B2(new_n710), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n720), .B(KEYINPUT108), .C1(new_n721), .C2(new_n539), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n718), .A2(new_n722), .ZN(G1329gat));
  INV_X1    g522(.A(KEYINPUT47), .ZN(new_n724));
  INV_X1    g523(.A(new_n671), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n541), .B1(new_n714), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n685), .A2(new_n541), .A3(new_n670), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT109), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n724), .B1(new_n726), .B2(new_n729), .ZN(new_n730));
  OAI211_X1 g529(.A(KEYINPUT47), .B(G43gat), .C1(new_n707), .C2(new_n671), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n731), .B(new_n727), .C1(new_n728), .C2(KEYINPUT47), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n730), .A2(new_n732), .ZN(G1330gat));
  NAND4_X1  g532(.A1(new_n690), .A2(new_n703), .A3(new_n259), .A4(new_n706), .ZN(new_n734));
  OR2_X1    g533(.A1(new_n734), .A2(KEYINPUT112), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(KEYINPUT112), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n735), .A2(G50gat), .A3(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n685), .A2(new_n543), .A3(new_n259), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT111), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n737), .A2(KEYINPUT48), .A3(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n738), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n714), .A2(new_n259), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n742), .B1(new_n743), .B2(G50gat), .ZN(new_n744));
  XNOR2_X1  g543(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n741), .B1(new_n744), .B2(new_n745), .ZN(G1331gat));
  INV_X1    g545(.A(KEYINPUT114), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n533), .A2(new_n678), .A3(new_n622), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(new_n704), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n749), .B(KEYINPUT113), .Z(new_n750));
  OR3_X1    g549(.A1(new_n477), .A2(new_n747), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n747), .B1(new_n477), .B2(new_n750), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n686), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g554(.A1(new_n751), .A2(new_n752), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n756), .A2(new_n465), .ZN(new_n757));
  NOR2_X1   g556(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n758));
  AND2_X1   g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(new_n757), .B2(new_n758), .ZN(G1333gat));
  NOR2_X1   g560(.A1(new_n756), .A2(new_n460), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n725), .A2(G71gat), .ZN(new_n763));
  OAI22_X1  g562(.A1(new_n762), .A2(G71gat), .B1(new_n756), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g564(.A1(new_n753), .A2(new_n259), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g566(.A1(new_n533), .A2(new_n683), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n592), .B(new_n768), .C1(new_n698), .C2(new_n702), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT51), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n773), .A2(new_n679), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n774), .A2(new_n564), .A3(new_n686), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n690), .A2(new_n703), .A3(new_n653), .A4(new_n768), .ZN(new_n776));
  OAI21_X1  g575(.A(G85gat), .B1(new_n776), .B2(new_n466), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(G1336gat));
  OAI21_X1  g577(.A(G92gat), .B1(new_n776), .B2(new_n465), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n704), .A2(new_n465), .A3(G92gat), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT115), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n779), .B1(new_n773), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g581(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n782), .B(new_n784), .ZN(G1337gat));
  INV_X1    g584(.A(G99gat), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n774), .A2(new_n786), .A3(new_n670), .ZN(new_n787));
  OAI21_X1  g586(.A(G99gat), .B1(new_n776), .B2(new_n671), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(G1338gat));
  OAI21_X1  g588(.A(G106gat), .B1(new_n776), .B2(new_n472), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n472), .A2(new_n704), .A3(G106gat), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n790), .B(new_n791), .C1(new_n773), .C2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(KEYINPUT117), .ZN(new_n795));
  OR2_X1    g594(.A1(new_n793), .A2(KEYINPUT117), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n795), .B(new_n796), .C1(new_n771), .C2(new_n772), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n797), .A2(new_n790), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n794), .B1(new_n798), .B2(new_n791), .ZN(G1339gat));
  NAND4_X1  g598(.A1(new_n533), .A2(new_n622), .A3(new_n678), .A4(new_n679), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT118), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n649), .A2(new_n629), .ZN(new_n803));
  OAI211_X1 g602(.A(KEYINPUT54), .B(new_n803), .C1(new_n641), .C2(new_n647), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n627), .B1(new_n650), .B2(new_n806), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n804), .A2(new_n805), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n805), .B1(new_n804), .B2(new_n807), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n648), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n680), .A2(new_n618), .A3(new_n611), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n597), .A2(new_n601), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n607), .A2(new_n608), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n617), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n811), .A2(new_n592), .A3(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n810), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n653), .A2(new_n811), .A3(new_n814), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n817), .B1(new_n810), .B2(new_n622), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n816), .B1(new_n818), .B2(new_n678), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n802), .B1(new_n533), .B2(new_n819), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n820), .A2(new_n686), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(new_n472), .A3(new_n470), .ZN(new_n822));
  OAI21_X1  g621(.A(G113gat), .B1(new_n822), .B2(new_n622), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n475), .A2(new_n469), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n622), .A2(G113gat), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(KEYINPUT119), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n823), .B1(new_n825), .B2(new_n827), .ZN(G1340gat));
  OAI21_X1  g627(.A(G120gat), .B1(new_n822), .B2(new_n704), .ZN(new_n829));
  OR2_X1    g628(.A1(new_n825), .A2(G120gat), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n829), .B1(new_n830), .B2(new_n679), .ZN(G1341gat));
  INV_X1    g630(.A(new_n825), .ZN(new_n832));
  AOI21_X1  g631(.A(G127gat), .B1(new_n832), .B2(new_n533), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n822), .A2(new_n534), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n833), .B1(G127gat), .B2(new_n834), .ZN(G1342gat));
  NOR3_X1   g634(.A1(new_n825), .A2(G134gat), .A3(new_n678), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(KEYINPUT56), .ZN(new_n837));
  OAI21_X1  g636(.A(G134gat), .B1(new_n822), .B2(new_n678), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(G1343gat));
  NAND2_X1  g638(.A1(new_n820), .A2(new_n259), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n725), .A2(new_n466), .A3(new_n469), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(G141gat), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n843), .A2(new_n844), .A3(new_n683), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(KEYINPUT58), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n805), .A2(KEYINPUT121), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n804), .A2(new_n807), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n848), .B1(new_n804), .B2(new_n807), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n648), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n817), .B1(new_n851), .B2(new_n622), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n816), .B1(new_n852), .B2(new_n678), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT122), .B1(new_n853), .B2(new_n533), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT122), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n804), .A2(new_n807), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n847), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n804), .A2(new_n807), .A3(new_n848), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(new_n683), .A3(new_n648), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n592), .B1(new_n860), .B2(new_n817), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n855), .B(new_n534), .C1(new_n861), .C2(new_n816), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n854), .A2(new_n802), .A3(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n472), .A2(new_n864), .ZN(new_n865));
  AND3_X1   g664(.A1(new_n863), .A2(KEYINPUT123), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT123), .B1(new_n863), .B2(new_n865), .ZN(new_n867));
  AOI21_X1  g666(.A(KEYINPUT57), .B1(new_n820), .B2(new_n259), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n842), .B(KEYINPUT120), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n869), .A2(new_n622), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n846), .B1(new_n844), .B2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT124), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n869), .A2(new_n873), .A3(new_n870), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n863), .A2(new_n865), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT123), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n840), .A2(new_n864), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n863), .A2(KEYINPUT123), .A3(new_n865), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n842), .B(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT124), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n683), .B1(new_n874), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n845), .B1(new_n884), .B2(G141gat), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT58), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n872), .B1(new_n885), .B2(new_n886), .ZN(G1344gat));
  INV_X1    g686(.A(G148gat), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n843), .A2(new_n888), .A3(new_n653), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n873), .B1(new_n869), .B2(new_n870), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n880), .A2(KEYINPUT124), .A3(new_n882), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n679), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n892), .A2(KEYINPUT59), .A3(new_n888), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n853), .A2(new_n533), .ZN(new_n895));
  INV_X1    g694(.A(new_n800), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n259), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n864), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n898), .B1(new_n840), .B2(new_n864), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n882), .A2(new_n653), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n894), .B1(new_n900), .B2(G148gat), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n889), .B1(new_n893), .B2(new_n901), .ZN(G1345gat));
  AOI21_X1  g701(.A(new_n206), .B1(new_n843), .B2(new_n533), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n534), .B1(new_n890), .B2(new_n891), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n903), .B1(new_n904), .B2(new_n206), .ZN(G1346gat));
  NOR3_X1   g704(.A1(new_n725), .A2(G162gat), .A3(new_n466), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n841), .A2(new_n465), .A3(new_n592), .A4(new_n906), .ZN(new_n907));
  XOR2_X1   g706(.A(new_n907), .B(KEYINPUT125), .Z(new_n908));
  AOI21_X1  g707(.A(new_n678), .B1(new_n890), .B2(new_n891), .ZN(new_n909));
  INV_X1    g708(.A(G162gat), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(G1347gat));
  NOR2_X1   g710(.A1(new_n465), .A2(new_n686), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n820), .A2(new_n472), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n670), .ZN(new_n914));
  OAI21_X1  g713(.A(G169gat), .B1(new_n914), .B2(new_n622), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n463), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n683), .A2(new_n282), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(G1348gat));
  NOR3_X1   g717(.A1(new_n914), .A2(new_n283), .A3(new_n704), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n913), .A2(new_n463), .A3(new_n653), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n919), .B1(new_n283), .B2(new_n920), .ZN(G1349gat));
  NAND2_X1  g720(.A1(new_n268), .A2(new_n270), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n922), .B1(new_n914), .B2(new_n534), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n533), .A2(new_n299), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n923), .B1(new_n916), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g725(.A(G190gat), .B1(new_n914), .B2(new_n678), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT61), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n913), .A2(new_n271), .A3(new_n463), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n928), .B1(new_n678), .B2(new_n929), .ZN(G1351gat));
  AND2_X1   g729(.A1(new_n899), .A2(new_n912), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(new_n671), .ZN(new_n932));
  OAI21_X1  g731(.A(G197gat), .B1(new_n932), .B2(new_n622), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n671), .A2(new_n912), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n841), .A2(new_n934), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n935), .A2(G197gat), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n933), .B1(new_n622), .B2(new_n936), .ZN(G1352gat));
  OR3_X1    g736(.A1(new_n932), .A2(KEYINPUT127), .A3(new_n704), .ZN(new_n938));
  OAI21_X1  g737(.A(KEYINPUT127), .B1(new_n932), .B2(new_n704), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n938), .A2(G204gat), .A3(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT126), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n935), .B1(new_n941), .B2(KEYINPUT62), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n942), .A2(new_n625), .A3(new_n653), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n941), .A2(KEYINPUT62), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n943), .B(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n940), .A2(new_n945), .ZN(G1353gat));
  NAND3_X1  g745(.A1(new_n931), .A2(new_n671), .A3(new_n533), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n947), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n948));
  AOI21_X1  g747(.A(KEYINPUT63), .B1(new_n947), .B2(G211gat), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n533), .A2(new_n221), .ZN(new_n950));
  OAI22_X1  g749(.A1(new_n948), .A2(new_n949), .B1(new_n935), .B2(new_n950), .ZN(G1354gat));
  NOR3_X1   g750(.A1(new_n932), .A2(new_n222), .A3(new_n678), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n841), .A2(new_n592), .A3(new_n934), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n952), .B1(new_n222), .B2(new_n953), .ZN(G1355gat));
endmodule


