//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 1 0 1 0 1 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n805, new_n806,
    new_n807, new_n808, new_n810, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n968, new_n969,
    new_n970, new_n971, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT12), .Z(new_n206));
  INV_X1    g005(.A(KEYINPUT18), .ZN(new_n207));
  NAND2_X1  g006(.A1(G229gat), .A2(G233gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT15), .ZN(new_n210));
  OR2_X1    g009(.A1(G43gat), .A2(G50gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(G43gat), .A2(G50gat), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(G29gat), .A2(G36gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n214), .B(KEYINPUT14), .ZN(new_n215));
  INV_X1    g014(.A(G29gat), .ZN(new_n216));
  INV_X1    g015(.A(G36gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n213), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n213), .A2(KEYINPUT91), .ZN(new_n220));
  INV_X1    g019(.A(new_n212), .ZN(new_n221));
  NOR2_X1   g020(.A1(G43gat), .A2(G50gat), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT15), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT91), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n221), .A2(KEYINPUT15), .ZN(new_n227));
  XNOR2_X1  g026(.A(KEYINPUT92), .B(G50gat), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n227), .B1(new_n228), .B2(G43gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT93), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT93), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n227), .B(new_n231), .C1(new_n228), .C2(G43gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n226), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n215), .A2(KEYINPUT94), .ZN(new_n234));
  OR2_X1    g033(.A1(new_n214), .A2(KEYINPUT14), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT94), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n214), .A2(KEYINPUT14), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n234), .B(new_n238), .C1(new_n216), .C2(new_n217), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n219), .B1(new_n233), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(G8gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(G15gat), .B(G22gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n242), .A2(G1gat), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G1gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT16), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n242), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n241), .B1(new_n244), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n247), .ZN(new_n249));
  NOR3_X1   g048(.A1(new_n249), .A2(new_n243), .A3(G8gat), .ZN(new_n250));
  OR2_X1    g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  AOI211_X1 g050(.A(new_n207), .B(new_n209), .C1(new_n240), .C2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT95), .B(KEYINPUT17), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n240), .A2(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n248), .A2(new_n250), .ZN(new_n256));
  OAI211_X1 g055(.A(KEYINPUT17), .B(new_n219), .C1(new_n233), .C2(new_n239), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n252), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n240), .A2(new_n251), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n256), .B(new_n219), .C1(new_n233), .C2(new_n239), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(new_n208), .B(KEYINPUT13), .Z(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n209), .B1(new_n240), .B2(new_n251), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT18), .B1(new_n258), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n206), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT96), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI211_X1 g069(.A(KEYINPUT96), .B(new_n206), .C1(new_n265), .C2(new_n267), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n258), .A2(new_n266), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(new_n207), .ZN(new_n274));
  AOI22_X1  g073(.A1(new_n252), .A2(new_n258), .B1(new_n262), .B2(new_n263), .ZN(new_n275));
  INV_X1    g074(.A(new_n206), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT97), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT97), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n274), .A2(new_n275), .A3(new_n279), .A4(new_n276), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n272), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT98), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n272), .A2(new_n281), .A3(KEYINPUT98), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(G57gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n288), .A2(KEYINPUT99), .ZN(new_n289));
  INV_X1    g088(.A(G64gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G71gat), .A2(G78gat), .ZN(new_n292));
  OR2_X1    g091(.A1(G71gat), .A2(G78gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT9), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n297), .B1(new_n288), .B2(new_n290), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n293), .A2(new_n292), .ZN(new_n299));
  AOI22_X1  g098(.A1(new_n291), .A2(new_n295), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n300), .A2(KEYINPUT21), .ZN(new_n301));
  XOR2_X1   g100(.A(G127gat), .B(G155gat), .Z(new_n302));
  XOR2_X1   g101(.A(new_n301), .B(new_n302), .Z(new_n303));
  AOI21_X1  g102(.A(new_n251), .B1(KEYINPUT21), .B2(new_n300), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n303), .B(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G231gat), .A2(G233gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n306), .B(KEYINPUT100), .ZN(new_n307));
  XOR2_X1   g106(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G183gat), .B(G211gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n309), .B(new_n310), .ZN(new_n311));
  OR2_X1    g110(.A1(new_n305), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n305), .A2(new_n311), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(KEYINPUT101), .B(G85gat), .ZN(new_n315));
  INV_X1    g114(.A(G92gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(G99gat), .A2(G106gat), .ZN(new_n317));
  AOI22_X1  g116(.A1(new_n315), .A2(new_n316), .B1(KEYINPUT8), .B2(new_n317), .ZN(new_n318));
  XOR2_X1   g117(.A(G99gat), .B(G106gat), .Z(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G85gat), .A2(G92gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n321), .B(KEYINPUT7), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n318), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n320), .B1(new_n318), .B2(new_n322), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n255), .B(new_n257), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G190gat), .B(G218gat), .ZN(new_n327));
  XOR2_X1   g126(.A(new_n327), .B(KEYINPUT102), .Z(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n324), .A2(new_n325), .ZN(new_n330));
  AND2_X1   g129(.A1(G232gat), .A2(G233gat), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n240), .A2(new_n330), .B1(KEYINPUT41), .B2(new_n331), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n326), .A2(new_n329), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n329), .B1(new_n326), .B2(new_n332), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n331), .A2(KEYINPUT41), .ZN(new_n335));
  XNOR2_X1  g134(.A(G134gat), .B(G162gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n335), .B(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  OR3_X1    g137(.A1(new_n333), .A2(new_n334), .A3(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n338), .B1(new_n333), .B2(new_n334), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(G230gat), .ZN(new_n342));
  INV_X1    g141(.A(G233gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AND2_X1   g143(.A1(new_n291), .A2(new_n295), .ZN(new_n345));
  AND2_X1   g144(.A1(new_n298), .A2(new_n299), .ZN(new_n346));
  OAI22_X1  g145(.A1(new_n324), .A2(new_n325), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n325), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n348), .A2(new_n300), .A3(new_n323), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT10), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n347), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n330), .A2(KEYINPUT10), .A3(new_n300), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n344), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n347), .A2(new_n349), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(new_n344), .ZN(new_n356));
  XNOR2_X1  g155(.A(G120gat), .B(G148gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(G176gat), .B(G204gat), .ZN(new_n358));
  XOR2_X1   g157(.A(new_n357), .B(new_n358), .Z(new_n359));
  NAND3_X1  g158(.A1(new_n354), .A2(new_n356), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n359), .B1(new_n354), .B2(new_n356), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n314), .A2(new_n341), .A3(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n364), .B(KEYINPUT103), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT90), .ZN(new_n366));
  XOR2_X1   g165(.A(G1gat), .B(G29gat), .Z(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G57gat), .B(G85gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n369), .B(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT78), .ZN(new_n372));
  NAND2_X1  g171(.A1(G225gat), .A2(G233gat), .ZN(new_n373));
  INV_X1    g172(.A(G120gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(G113gat), .ZN(new_n375));
  INV_X1    g174(.A(G113gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(G120gat), .ZN(new_n377));
  AOI21_X1  g176(.A(KEYINPUT1), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(G127gat), .A2(G134gat), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(G127gat), .A2(G134gat), .ZN(new_n381));
  NOR3_X1   g180(.A1(new_n380), .A2(new_n381), .A3(KEYINPUT67), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT67), .ZN(new_n383));
  INV_X1    g182(.A(G127gat), .ZN(new_n384));
  INV_X1    g183(.A(G134gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n383), .B1(new_n386), .B2(new_n379), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n378), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT1), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n376), .A2(G120gat), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n374), .A2(G113gat), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n386), .A2(KEYINPUT66), .A3(new_n379), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT66), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n394), .B1(new_n380), .B2(new_n381), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n392), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n388), .A2(new_n396), .ZN(new_n397));
  XOR2_X1   g196(.A(G141gat), .B(G148gat), .Z(new_n398));
  INV_X1    g197(.A(G155gat), .ZN(new_n399));
  INV_X1    g198(.A(G162gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(G155gat), .A2(G162gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(KEYINPUT2), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n398), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G141gat), .B(G148gat), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n402), .B(new_n401), .C1(new_n406), .C2(KEYINPUT2), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n397), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n388), .A2(new_n396), .A3(new_n407), .A4(new_n405), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n373), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT77), .ZN(new_n412));
  OAI21_X1  g211(.A(KEYINPUT5), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  AOI211_X1 g212(.A(KEYINPUT77), .B(new_n373), .C1(new_n409), .C2(new_n410), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n372), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n397), .A2(new_n408), .ZN(new_n416));
  AOI22_X1  g215(.A1(new_n388), .A2(new_n396), .B1(new_n407), .B2(new_n405), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT77), .B1(new_n418), .B2(new_n373), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n411), .A2(new_n412), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n419), .A2(new_n420), .A3(KEYINPUT78), .A4(KEYINPUT5), .ZN(new_n421));
  INV_X1    g220(.A(new_n373), .ZN(new_n422));
  AOI22_X1  g221(.A1(new_n408), .A2(KEYINPUT3), .B1(new_n388), .B2(new_n396), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT3), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n405), .A2(new_n407), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n422), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n397), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT75), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n408), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n405), .A2(new_n407), .A3(KEYINPUT75), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n427), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT76), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(new_n432), .A3(KEYINPUT4), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n431), .A2(KEYINPUT4), .ZN(new_n434));
  OAI21_X1  g233(.A(KEYINPUT76), .B1(new_n410), .B2(KEYINPUT4), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n426), .B(new_n433), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n415), .A2(new_n421), .A3(new_n436), .ZN(new_n437));
  AOI211_X1 g236(.A(KEYINPUT5), .B(new_n422), .C1(new_n423), .C2(new_n425), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT80), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT4), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n427), .A2(new_n429), .A3(new_n440), .A4(new_n430), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n410), .A2(KEYINPUT4), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n438), .A2(new_n439), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n439), .B1(new_n438), .B2(new_n443), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n371), .B1(new_n437), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT6), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT6), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n437), .A2(new_n446), .A3(new_n371), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n449), .B(new_n450), .C1(new_n447), .C2(KEYINPUT81), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n437), .A2(new_n446), .ZN(new_n452));
  INV_X1    g251(.A(new_n371), .ZN(new_n453));
  AND3_X1   g252(.A1(new_n452), .A2(KEYINPUT81), .A3(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n448), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(G8gat), .B(G36gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(G64gat), .B(G92gat), .ZN(new_n457));
  XOR2_X1   g256(.A(new_n456), .B(new_n457), .Z(new_n458));
  NAND2_X1  g257(.A1(G226gat), .A2(G233gat), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(KEYINPUT27), .B(G183gat), .ZN(new_n461));
  INV_X1    g260(.A(G190gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT28), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n461), .A2(KEYINPUT28), .A3(new_n462), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g266(.A1(G169gat), .A2(G176gat), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT26), .ZN(new_n470));
  NAND2_X1  g269(.A1(G169gat), .A2(G176gat), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n468), .A2(KEYINPUT26), .ZN(new_n473));
  NAND2_X1  g272(.A1(G183gat), .A2(G190gat), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n467), .A2(new_n472), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT24), .ZN(new_n477));
  INV_X1    g276(.A(G183gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(G190gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n462), .A2(G183gat), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n468), .B1(KEYINPUT23), .B2(new_n471), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n474), .A2(KEYINPUT24), .ZN(new_n483));
  NOR3_X1   g282(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(G169gat), .ZN(new_n485));
  INV_X1    g284(.A(G176gat), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n485), .A2(new_n486), .A3(KEYINPUT23), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT64), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT64), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n468), .A2(new_n489), .A3(KEYINPUT23), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT25), .B1(new_n484), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n471), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT23), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n469), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n495), .A2(KEYINPUT25), .A3(new_n487), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT65), .B1(new_n481), .B2(new_n483), .ZN(new_n497));
  INV_X1    g296(.A(new_n483), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT65), .ZN(new_n499));
  XNOR2_X1  g298(.A(G183gat), .B(G190gat), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n498), .B(new_n499), .C1(new_n500), .C2(new_n477), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n496), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n476), .B1(new_n492), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT29), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n460), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n475), .A2(new_n472), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n506), .B1(new_n465), .B2(new_n466), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n497), .A2(new_n501), .ZN(new_n508));
  INV_X1    g307(.A(new_n496), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n479), .A2(new_n480), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n483), .B1(new_n511), .B2(KEYINPUT24), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n512), .A2(new_n491), .A3(new_n495), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT25), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n507), .B1(new_n510), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n516), .A2(new_n459), .ZN(new_n517));
  NOR2_X1   g316(.A1(G197gat), .A2(G204gat), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(G197gat), .A2(G204gat), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT22), .ZN(new_n521));
  NAND2_X1  g320(.A1(G211gat), .A2(G218gat), .ZN(new_n522));
  AOI22_X1  g321(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AND2_X1   g322(.A1(G211gat), .A2(G218gat), .ZN(new_n524));
  NOR2_X1   g323(.A1(G211gat), .A2(G218gat), .ZN(new_n525));
  NOR3_X1   g324(.A1(new_n524), .A2(new_n525), .A3(KEYINPUT72), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT72), .ZN(new_n527));
  OR2_X1    g326(.A1(G211gat), .A2(G218gat), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n527), .B1(new_n528), .B2(new_n522), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n523), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT73), .ZN(new_n531));
  INV_X1    g330(.A(new_n520), .ZN(new_n532));
  OAI22_X1  g331(.A1(new_n532), .A2(new_n518), .B1(new_n524), .B2(KEYINPUT22), .ZN(new_n533));
  OAI21_X1  g332(.A(KEYINPUT72), .B1(new_n524), .B2(new_n525), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n528), .A2(new_n527), .A3(new_n522), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n530), .A2(new_n531), .A3(new_n536), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n533), .A2(KEYINPUT73), .A3(new_n534), .A4(new_n535), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NOR3_X1   g339(.A1(new_n505), .A2(new_n517), .A3(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n459), .B1(new_n516), .B2(KEYINPUT29), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n503), .A2(new_n460), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n539), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n458), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT30), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n540), .B1(new_n505), .B2(new_n517), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n542), .A2(new_n539), .A3(new_n543), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n550), .A2(KEYINPUT30), .A3(new_n458), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT74), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n548), .A2(new_n549), .A3(KEYINPUT74), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n458), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n455), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT82), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n455), .A2(KEYINPUT82), .A3(new_n557), .ZN(new_n561));
  XNOR2_X1  g360(.A(G78gat), .B(G106gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(G22gat), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(G228gat), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n565), .A2(new_n343), .ZN(new_n566));
  INV_X1    g365(.A(new_n425), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n539), .B1(KEYINPUT29), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n408), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n537), .A2(new_n504), .A3(new_n538), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT3), .B1(new_n570), .B2(KEYINPUT83), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT83), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n537), .A2(new_n572), .A3(new_n504), .A4(new_n538), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n569), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT84), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n568), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AOI211_X1 g375(.A(KEYINPUT84), .B(new_n569), .C1(new_n571), .C2(new_n573), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n566), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n429), .A2(new_n430), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT29), .B1(new_n530), .B2(new_n536), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n579), .B1(KEYINPUT3), .B2(new_n580), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n581), .B(new_n568), .C1(new_n565), .C2(new_n343), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT31), .B(G50gat), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  AND3_X1   g383(.A1(new_n578), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n584), .B1(new_n578), .B2(new_n582), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n564), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n578), .A2(new_n582), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(new_n583), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n578), .A2(new_n582), .A3(new_n584), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n589), .A2(new_n563), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n587), .A2(new_n591), .A3(KEYINPUT85), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n587), .A2(new_n591), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT85), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n560), .A2(new_n561), .B1(new_n592), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT38), .ZN(new_n597));
  INV_X1    g396(.A(new_n555), .ZN(new_n598));
  AOI21_X1  g397(.A(KEYINPUT74), .B1(new_n548), .B2(new_n549), .ZN(new_n599));
  OAI21_X1  g398(.A(KEYINPUT37), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(KEYINPUT89), .B(KEYINPUT37), .Z(new_n601));
  AOI21_X1  g400(.A(new_n458), .B1(new_n550), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n597), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n548), .A2(new_n549), .A3(KEYINPUT37), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n602), .A2(new_n597), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n545), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n450), .A2(new_n449), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n452), .A2(KEYINPUT87), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(new_n453), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT87), .ZN(new_n611));
  AND3_X1   g410(.A1(new_n437), .A2(new_n446), .A3(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n608), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n607), .A2(new_n613), .A3(new_n448), .ZN(new_n614));
  INV_X1    g413(.A(new_n593), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n418), .A2(new_n373), .ZN(new_n616));
  AOI22_X1  g415(.A1(new_n441), .A2(new_n442), .B1(new_n425), .B2(new_n423), .ZN(new_n617));
  OAI211_X1 g416(.A(KEYINPUT39), .B(new_n616), .C1(new_n617), .C2(new_n373), .ZN(new_n618));
  XNOR2_X1  g417(.A(KEYINPUT86), .B(KEYINPUT39), .ZN(new_n619));
  AND2_X1   g418(.A1(new_n441), .A2(new_n442), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n423), .A2(new_n425), .ZN(new_n621));
  OAI211_X1 g420(.A(new_n422), .B(new_n619), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n618), .A2(new_n622), .A3(KEYINPUT40), .A4(new_n371), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT88), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n617), .A2(new_n373), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n453), .B1(new_n625), .B2(new_n619), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT88), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n626), .A2(new_n627), .A3(KEYINPUT40), .A4(new_n618), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(new_n618), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT40), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n629), .B(new_n632), .C1(new_n552), .C2(new_n556), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n611), .B1(new_n437), .B2(new_n446), .ZN(new_n634));
  NOR3_X1   g433(.A1(new_n612), .A2(new_n634), .A3(new_n371), .ZN(new_n635));
  OR2_X1    g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n614), .A2(new_n615), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT36), .ZN(new_n638));
  AOI22_X1  g437(.A1(new_n508), .A2(new_n509), .B1(new_n513), .B2(new_n514), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n427), .B1(new_n639), .B2(new_n507), .ZN(new_n640));
  NAND2_X1  g439(.A1(G227gat), .A2(G233gat), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  OAI211_X1 g441(.A(new_n476), .B(new_n397), .C1(new_n492), .C2(new_n502), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n640), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(KEYINPUT32), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT68), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n644), .A2(KEYINPUT68), .A3(KEYINPUT32), .ZN(new_n648));
  XNOR2_X1  g447(.A(G15gat), .B(G43gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(G71gat), .B(G99gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT33), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n651), .B1(new_n644), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n647), .A2(new_n648), .A3(new_n653), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n651), .A2(new_n652), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n644), .A2(KEYINPUT32), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT69), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n644), .A2(KEYINPUT69), .A3(KEYINPUT32), .A4(new_n655), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n642), .B1(new_n640), .B2(new_n643), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT34), .ZN(new_n662));
  AND3_X1   g461(.A1(new_n654), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n662), .B1(new_n654), .B2(new_n660), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n638), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT71), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI211_X1 g466(.A(KEYINPUT71), .B(new_n638), .C1(new_n663), .C2(new_n664), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT70), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n663), .A2(new_n664), .A3(new_n670), .ZN(new_n671));
  AOI211_X1 g470(.A(KEYINPUT70), .B(new_n662), .C1(new_n654), .C2(new_n660), .ZN(new_n672));
  OAI21_X1  g471(.A(KEYINPUT36), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n637), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n596), .A2(new_n675), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n613), .A2(new_n448), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n663), .A2(new_n664), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT35), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n678), .A2(new_n679), .A3(new_n557), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n677), .A2(new_n680), .A3(new_n593), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n672), .B1(new_n678), .B2(KEYINPUT70), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n682), .A2(new_n593), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n560), .A2(new_n683), .A3(new_n561), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n681), .B1(new_n684), .B2(KEYINPUT35), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n366), .B1(new_n676), .B2(new_n685), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n591), .B(new_n587), .C1(new_n633), .C2(new_n635), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  AOI22_X1  g487(.A1(new_n688), .A2(new_n614), .B1(new_n669), .B2(new_n673), .ZN(new_n689));
  AND3_X1   g488(.A1(new_n455), .A2(KEYINPUT82), .A3(new_n557), .ZN(new_n690));
  AOI21_X1  g489(.A(KEYINPUT82), .B1(new_n455), .B2(new_n557), .ZN(new_n691));
  INV_X1    g490(.A(new_n592), .ZN(new_n692));
  AOI21_X1  g491(.A(KEYINPUT85), .B1(new_n587), .B2(new_n591), .ZN(new_n693));
  OAI22_X1  g492(.A1(new_n690), .A2(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n689), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n690), .A2(new_n691), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n679), .B1(new_n696), .B2(new_n683), .ZN(new_n697));
  OAI211_X1 g496(.A(new_n695), .B(KEYINPUT90), .C1(new_n697), .C2(new_n681), .ZN(new_n698));
  AOI211_X1 g497(.A(new_n287), .B(new_n365), .C1(new_n686), .C2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(new_n455), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(new_n245), .ZN(G1324gat));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n703));
  INV_X1    g502(.A(new_n557), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n241), .B1(new_n699), .B2(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n287), .B1(new_n686), .B2(new_n698), .ZN(new_n706));
  INV_X1    g505(.A(new_n365), .ZN(new_n707));
  XOR2_X1   g506(.A(KEYINPUT16), .B(G8gat), .Z(new_n708));
  AND4_X1   g507(.A1(new_n704), .A2(new_n706), .A3(new_n707), .A4(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT42), .B1(new_n705), .B2(new_n709), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n706), .A2(new_n704), .A3(new_n707), .A4(new_n708), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT42), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n703), .B1(new_n710), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n686), .A2(new_n698), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n715), .A2(new_n704), .A3(new_n286), .A4(new_n707), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(G8gat), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n712), .B1(new_n717), .B2(new_n711), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n711), .A2(new_n712), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n718), .A2(new_n719), .A3(KEYINPUT104), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n714), .A2(new_n720), .ZN(G1325gat));
  OAI21_X1  g520(.A(G15gat), .B1(new_n700), .B2(new_n674), .ZN(new_n722));
  INV_X1    g521(.A(new_n678), .ZN(new_n723));
  OR2_X1    g522(.A1(new_n723), .A2(G15gat), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n722), .B1(new_n700), .B2(new_n724), .ZN(G1326gat));
  NOR2_X1   g524(.A1(new_n692), .A2(new_n693), .ZN(new_n726));
  OAI21_X1  g525(.A(KEYINPUT105), .B1(new_n700), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT105), .ZN(new_n728));
  INV_X1    g527(.A(new_n726), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n699), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(KEYINPUT43), .B(G22gat), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n727), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n731), .B1(new_n727), .B2(new_n730), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(G1327gat));
  INV_X1    g533(.A(new_n314), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n363), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n736), .A2(new_n341), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n706), .A2(new_n737), .ZN(new_n738));
  OR3_X1    g537(.A1(new_n738), .A2(G29gat), .A3(new_n455), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT45), .ZN(new_n740));
  OR2_X1    g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n341), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n744), .B1(new_n686), .B2(new_n698), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n695), .B1(new_n697), .B2(new_n681), .ZN(new_n746));
  INV_X1    g545(.A(new_n341), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT44), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n282), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n736), .A2(new_n750), .ZN(new_n751));
  XOR2_X1   g550(.A(new_n751), .B(KEYINPUT106), .Z(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(G29gat), .B1(new_n754), .B2(new_n455), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n741), .A2(new_n755), .A3(new_n756), .ZN(G1328gat));
  AND2_X1   g556(.A1(new_n706), .A2(new_n737), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n758), .A2(new_n217), .A3(new_n704), .ZN(new_n759));
  OR2_X1    g558(.A1(new_n759), .A2(KEYINPUT46), .ZN(new_n760));
  OAI21_X1  g559(.A(G36gat), .B1(new_n754), .B2(new_n557), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(KEYINPUT46), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(G1329gat));
  NOR2_X1   g562(.A1(new_n723), .A2(G43gat), .ZN(new_n764));
  AND4_X1   g563(.A1(new_n715), .A2(new_n286), .A3(new_n737), .A4(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NOR4_X1   g565(.A1(new_n745), .A2(new_n748), .A3(new_n674), .A4(new_n752), .ZN(new_n767));
  INV_X1    g566(.A(G43gat), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT47), .B1(new_n769), .B2(KEYINPUT107), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n715), .A2(new_n743), .ZN(new_n771));
  INV_X1    g570(.A(new_n748), .ZN(new_n772));
  INV_X1    g571(.A(new_n674), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n771), .A2(new_n772), .A3(new_n773), .A4(new_n753), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n765), .B1(new_n774), .B2(G43gat), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT107), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT47), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n770), .A2(new_n778), .ZN(G1330gat));
  NOR2_X1   g578(.A1(new_n726), .A2(new_n228), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n758), .A2(new_n780), .ZN(new_n781));
  NOR4_X1   g580(.A1(new_n745), .A2(new_n748), .A3(new_n726), .A4(new_n752), .ZN(new_n782));
  INV_X1    g581(.A(new_n228), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT48), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n785), .B1(new_n758), .B2(new_n780), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n771), .A2(new_n772), .A3(new_n593), .A4(new_n753), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n228), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT108), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n787), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n790), .B1(new_n787), .B2(new_n789), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n786), .B1(new_n791), .B2(new_n792), .ZN(G1331gat));
  NOR4_X1   g592(.A1(new_n282), .A2(new_n735), .A3(new_n747), .A4(new_n363), .ZN(new_n794));
  XOR2_X1   g593(.A(new_n794), .B(KEYINPUT109), .Z(new_n795));
  AND2_X1   g594(.A1(new_n746), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n455), .B(KEYINPUT110), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g598(.A(new_n557), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(KEYINPUT111), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n796), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n803));
  XOR2_X1   g602(.A(new_n802), .B(new_n803), .Z(G1333gat));
  NAND2_X1  g603(.A1(new_n796), .A2(new_n773), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n723), .A2(G71gat), .ZN(new_n806));
  AOI22_X1  g605(.A1(new_n805), .A2(G71gat), .B1(new_n796), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g606(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n807), .B(new_n808), .ZN(G1334gat));
  NAND2_X1  g608(.A1(new_n796), .A2(new_n729), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(G78gat), .ZN(G1335gat));
  INV_X1    g610(.A(new_n749), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n282), .A2(new_n314), .ZN(new_n813));
  INV_X1    g612(.A(new_n363), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n812), .A2(new_n455), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n746), .A2(new_n747), .A3(new_n813), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT51), .ZN(new_n818));
  OR2_X1    g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n818), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n814), .A2(new_n315), .ZN(new_n823));
  OR2_X1    g622(.A1(new_n455), .A2(new_n823), .ZN(new_n824));
  OAI22_X1  g623(.A1(new_n816), .A2(new_n315), .B1(new_n822), .B2(new_n824), .ZN(G1336gat));
  NAND3_X1  g624(.A1(new_n704), .A2(new_n316), .A3(new_n814), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(KEYINPUT113), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n821), .A2(new_n827), .ZN(new_n828));
  NOR4_X1   g627(.A1(new_n745), .A2(new_n748), .A3(new_n557), .A4(new_n815), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n828), .B1(new_n829), .B2(new_n316), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT114), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n831), .B1(new_n829), .B2(new_n316), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n830), .A2(KEYINPUT52), .A3(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n834));
  OAI221_X1 g633(.A(new_n828), .B1(new_n831), .B2(new_n834), .C1(new_n829), .C2(new_n316), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(G1337gat));
  NOR3_X1   g635(.A1(new_n812), .A2(new_n674), .A3(new_n815), .ZN(new_n837));
  INV_X1    g636(.A(G99gat), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n678), .A2(new_n838), .A3(new_n814), .ZN(new_n839));
  XOR2_X1   g638(.A(new_n839), .B(KEYINPUT115), .Z(new_n840));
  OAI22_X1  g639(.A1(new_n837), .A2(new_n838), .B1(new_n822), .B2(new_n840), .ZN(G1338gat));
  NOR3_X1   g640(.A1(new_n615), .A2(G106gat), .A3(new_n363), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT53), .B1(new_n821), .B2(new_n842), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n812), .A2(new_n615), .A3(new_n815), .ZN(new_n844));
  INV_X1    g643(.A(G106gat), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n749), .A2(new_n729), .A3(new_n814), .A4(new_n813), .ZN(new_n847));
  AOI22_X1  g646(.A1(new_n847), .A2(G106gat), .B1(new_n821), .B2(new_n842), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n846), .B1(new_n848), .B2(new_n849), .ZN(G1339gat));
  NOR2_X1   g649(.A1(new_n364), .A2(new_n282), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n208), .B1(new_n258), .B2(new_n260), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n262), .A2(new_n263), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n205), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n281), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n747), .B1(new_n855), .B2(KEYINPUT118), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n857), .B1(new_n281), .B2(new_n854), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n351), .A2(new_n352), .A3(new_n344), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n354), .A2(KEYINPUT54), .A3(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n353), .A2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n359), .ZN(new_n864));
  AOI21_X1  g663(.A(KEYINPUT116), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT116), .ZN(new_n866));
  AOI211_X1 g665(.A(new_n866), .B(new_n359), .C1(new_n353), .C2(new_n862), .ZN(new_n867));
  OAI211_X1 g666(.A(KEYINPUT55), .B(new_n861), .C1(new_n865), .C2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n360), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(KEYINPUT117), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT117), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n868), .A2(new_n871), .A3(new_n360), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n861), .B1(new_n865), .B2(new_n867), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT55), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n870), .A2(new_n872), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n859), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n855), .A2(new_n363), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n878), .B1(new_n876), .B2(new_n282), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n877), .B1(new_n879), .B2(new_n747), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n851), .B1(new_n880), .B2(new_n735), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n678), .A2(new_n557), .ZN(new_n882));
  OR4_X1    g681(.A1(new_n455), .A2(new_n881), .A3(new_n882), .A4(new_n729), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n883), .A2(new_n376), .A3(new_n287), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n880), .A2(new_n735), .ZN(new_n885));
  INV_X1    g684(.A(new_n851), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n887), .A2(new_n797), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(new_n557), .A3(new_n683), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n889), .A2(new_n750), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n884), .B1(new_n890), .B2(new_n376), .ZN(G1340gat));
  NOR3_X1   g690(.A1(new_n883), .A2(new_n374), .A3(new_n363), .ZN(new_n892));
  OR2_X1    g691(.A1(new_n889), .A2(new_n363), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n892), .B1(new_n893), .B2(new_n374), .ZN(G1341gat));
  NOR3_X1   g693(.A1(new_n883), .A2(new_n384), .A3(new_n735), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n889), .A2(new_n735), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n896), .A2(KEYINPUT119), .ZN(new_n897));
  AOI21_X1  g696(.A(G127gat), .B1(new_n896), .B2(KEYINPUT119), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n895), .B1(new_n897), .B2(new_n898), .ZN(G1342gat));
  OR3_X1    g698(.A1(new_n889), .A2(G134gat), .A3(new_n341), .ZN(new_n900));
  OR2_X1    g699(.A1(new_n900), .A2(KEYINPUT56), .ZN(new_n901));
  OAI21_X1  g700(.A(G134gat), .B1(new_n883), .B2(new_n341), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(KEYINPUT56), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(G1343gat));
  NOR3_X1   g703(.A1(new_n773), .A2(new_n704), .A3(new_n615), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n888), .A2(new_n905), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n906), .A2(G141gat), .A3(new_n287), .ZN(new_n907));
  XOR2_X1   g706(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n908));
  NOR2_X1   g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n875), .A2(new_n360), .A3(new_n868), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n910), .B1(new_n284), .B2(new_n285), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n341), .B1(new_n911), .B2(new_n878), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n314), .B1(new_n912), .B2(new_n877), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n913), .A2(new_n851), .ZN(new_n914));
  OAI21_X1  g713(.A(KEYINPUT57), .B1(new_n914), .B2(new_n726), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n773), .A2(new_n455), .A3(new_n704), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n887), .A2(new_n593), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n915), .B(new_n916), .C1(KEYINPUT57), .C2(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(G141gat), .B1(new_n918), .B2(new_n287), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n909), .A2(new_n919), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n918), .A2(new_n750), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n907), .B1(new_n921), .B2(G141gat), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT58), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(G1344gat));
  OAI21_X1  g723(.A(G148gat), .B1(new_n918), .B2(new_n363), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT59), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OR3_X1    g726(.A1(new_n906), .A2(G148gat), .A3(new_n363), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT121), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n365), .A2(new_n286), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n929), .B1(new_n913), .B2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(new_n930), .ZN(new_n932));
  INV_X1    g731(.A(new_n910), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n272), .A2(new_n281), .A3(KEYINPUT98), .ZN(new_n934));
  AOI21_X1  g733(.A(KEYINPUT98), .B1(new_n272), .B2(new_n281), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(new_n878), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI22_X1  g737(.A1(new_n938), .A2(new_n341), .B1(new_n876), .B2(new_n859), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n932), .B(KEYINPUT121), .C1(new_n939), .C2(new_n314), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n726), .A2(KEYINPUT57), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n931), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g741(.A(KEYINPUT57), .B1(new_n881), .B2(new_n615), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AND3_X1   g743(.A1(new_n944), .A2(new_n814), .A3(new_n916), .ZN(new_n945));
  NAND2_X1  g744(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n927), .B(new_n928), .C1(new_n945), .C2(new_n946), .ZN(G1345gat));
  OAI21_X1  g746(.A(G155gat), .B1(new_n918), .B2(new_n735), .ZN(new_n948));
  INV_X1    g747(.A(new_n906), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n949), .A2(new_n399), .A3(new_n314), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(G1346gat));
  OAI21_X1  g750(.A(G162gat), .B1(new_n918), .B2(new_n341), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n949), .A2(new_n400), .A3(new_n747), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(G1347gat));
  OR2_X1    g753(.A1(new_n797), .A2(new_n557), .ZN(new_n955));
  OR4_X1    g754(.A1(new_n723), .A2(new_n881), .A3(new_n729), .A4(new_n955), .ZN(new_n956));
  OAI21_X1  g755(.A(G169gat), .B1(new_n956), .B2(new_n287), .ZN(new_n957));
  XOR2_X1   g756(.A(new_n957), .B(KEYINPUT122), .Z(new_n958));
  AND2_X1   g757(.A1(new_n887), .A2(new_n455), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n682), .A2(new_n593), .A3(new_n557), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n962), .A2(new_n485), .A3(new_n282), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n958), .A2(new_n963), .ZN(G1348gat));
  OAI21_X1  g763(.A(G176gat), .B1(new_n956), .B2(new_n363), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n814), .A2(new_n486), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n965), .B1(new_n961), .B2(new_n966), .ZN(G1349gat));
  OAI21_X1  g766(.A(G183gat), .B1(new_n956), .B2(new_n735), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n314), .A2(new_n461), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n968), .B1(new_n961), .B2(new_n969), .ZN(new_n970));
  XOR2_X1   g769(.A(KEYINPUT123), .B(KEYINPUT60), .Z(new_n971));
  XNOR2_X1  g770(.A(new_n970), .B(new_n971), .ZN(G1350gat));
  OAI21_X1  g771(.A(G190gat), .B1(new_n956), .B2(new_n341), .ZN(new_n973));
  XNOR2_X1  g772(.A(new_n973), .B(KEYINPUT61), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n962), .A2(new_n462), .A3(new_n747), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(G1351gat));
  NOR3_X1   g775(.A1(new_n773), .A2(new_n557), .A3(new_n615), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n959), .A2(new_n977), .ZN(new_n978));
  NOR3_X1   g777(.A1(new_n978), .A2(G197gat), .A3(new_n750), .ZN(new_n979));
  XNOR2_X1  g778(.A(new_n979), .B(KEYINPUT124), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT125), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n955), .A2(new_n773), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n944), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n981), .B1(new_n983), .B2(new_n287), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n984), .A2(G197gat), .ZN(new_n985));
  NOR3_X1   g784(.A1(new_n983), .A2(new_n981), .A3(new_n287), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n980), .B1(new_n985), .B2(new_n986), .ZN(G1352gat));
  OAI21_X1  g786(.A(G204gat), .B1(new_n983), .B2(new_n363), .ZN(new_n988));
  NOR3_X1   g787(.A1(new_n978), .A2(G204gat), .A3(new_n363), .ZN(new_n989));
  NAND2_X1  g788(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  XOR2_X1   g790(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n992));
  OAI211_X1 g791(.A(new_n988), .B(new_n991), .C1(new_n989), .C2(new_n992), .ZN(G1353gat));
  OR3_X1    g792(.A1(new_n978), .A2(G211gat), .A3(new_n735), .ZN(new_n994));
  NAND4_X1  g793(.A1(new_n942), .A2(new_n314), .A3(new_n943), .A4(new_n982), .ZN(new_n995));
  AND3_X1   g794(.A1(new_n995), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n996));
  AOI21_X1  g795(.A(KEYINPUT63), .B1(new_n995), .B2(G211gat), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n994), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n998), .A2(KEYINPUT127), .ZN(new_n999));
  INV_X1    g798(.A(KEYINPUT127), .ZN(new_n1000));
  OAI211_X1 g799(.A(new_n994), .B(new_n1000), .C1(new_n996), .C2(new_n997), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n999), .A2(new_n1001), .ZN(G1354gat));
  OAI21_X1  g801(.A(G218gat), .B1(new_n983), .B2(new_n341), .ZN(new_n1003));
  OR2_X1    g802(.A1(new_n341), .A2(G218gat), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n1003), .B1(new_n978), .B2(new_n1004), .ZN(G1355gat));
endmodule


