//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 0 0 1 0 0 0 0 1 1 0 1 0 0 1 1 0 0 1 0 1 1 1 0 0 0 0 0 0 1 0 0 1 0 0 0 1 0 1 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n221, new_n222, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n230, new_n231, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(new_n204));
  AOI22_X1  g0004(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n208));
  NAND4_X1  g0008(.A1(new_n205), .A2(new_n206), .A3(new_n207), .A4(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n204), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT1), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n204), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT0), .Z(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  AOI211_X1 g0019(.A(new_n211), .B(new_n214), .C1(new_n217), .C2(new_n219), .ZN(G361));
  XNOR2_X1  g0020(.A(G238), .B(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G232), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n221), .B(new_n222), .ZN(new_n223));
  XOR2_X1   g0023(.A(KEYINPUT2), .B(G226), .Z(new_n224));
  XNOR2_X1  g0024(.A(new_n223), .B(new_n224), .ZN(new_n225));
  XOR2_X1   g0025(.A(G264), .B(G270), .Z(new_n226));
  XNOR2_X1  g0026(.A(G250), .B(G257), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n225), .B(new_n228), .ZN(G358));
  INV_X1    g0029(.A(G50), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G68), .ZN(new_n231));
  INV_X1    g0031(.A(G68), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G50), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G58), .B(G77), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  INV_X1    g0036(.A(G107), .ZN(new_n237));
  NAND2_X1  g0037(.A1(new_n237), .A2(G97), .ZN(new_n238));
  INV_X1    g0038(.A(G97), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n239), .A2(G107), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G87), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n236), .B(new_n243), .ZN(G351));
  NAND3_X1  g0044(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(new_n215), .ZN(new_n246));
  NOR2_X1   g0046(.A1(G58), .A2(G68), .ZN(new_n247));
  AOI21_X1  g0047(.A(new_n216), .B1(new_n247), .B2(new_n230), .ZN(new_n248));
  OR2_X1    g0048(.A1(new_n248), .A2(KEYINPUT68), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(KEYINPUT68), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G150), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT8), .B(G58), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n216), .A2(G33), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT67), .ZN(new_n256));
  OAI211_X1 g0056(.A(new_n249), .B(new_n250), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  AND2_X1   g0057(.A1(new_n255), .A2(new_n256), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n246), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT69), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT69), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n261), .B(new_n246), .C1(new_n257), .C2(new_n258), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(G13), .A3(G20), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(new_n246), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n230), .B1(new_n263), .B2(G20), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n266), .A2(new_n267), .B1(new_n230), .B2(new_n265), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n260), .A2(new_n262), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT9), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n260), .A2(KEYINPUT9), .A3(new_n262), .A4(new_n268), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT66), .ZN(new_n273));
  INV_X1    g0073(.A(G41), .ZN(new_n274));
  INV_X1    g0074(.A(G45), .ZN(new_n275));
  AOI21_X1  g0075(.A(G1), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(G1), .A3(G13), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n276), .A2(new_n278), .A3(G274), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n263), .B1(G41), .B2(G45), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n280), .B1(G226), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT3), .ZN(new_n285));
  INV_X1    g0085(.A(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G1698), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n289), .A2(G222), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(KEYINPUT65), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT65), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n289), .A2(new_n293), .A3(G222), .A4(new_n290), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n290), .B1(new_n287), .B2(new_n288), .ZN(new_n296));
  AND2_X1   g0096(.A1(KEYINPUT3), .A2(G33), .ZN(new_n297));
  NOR2_X1   g0097(.A1(KEYINPUT3), .A2(G33), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n296), .A2(G223), .B1(new_n299), .B2(G77), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n295), .A2(new_n300), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n273), .B(new_n284), .C1(new_n301), .C2(new_n278), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n278), .B1(new_n295), .B2(new_n300), .ZN(new_n303));
  INV_X1    g0103(.A(new_n284), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT66), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n302), .A2(G200), .A3(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n271), .A2(new_n272), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT10), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT70), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n302), .A2(new_n305), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n310), .B1(new_n311), .B2(G190), .ZN(new_n312));
  INV_X1    g0112(.A(G190), .ZN(new_n313));
  AOI211_X1 g0113(.A(KEYINPUT70), .B(new_n313), .C1(new_n302), .C2(new_n305), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n308), .B(new_n309), .C1(new_n312), .C2(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n312), .A2(new_n314), .ZN(new_n316));
  OAI21_X1  g0116(.A(KEYINPUT10), .B1(new_n316), .B2(new_n307), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G179), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n311), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G169), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n305), .A2(new_n302), .A3(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n320), .A2(new_n269), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  NOR3_X1   g0124(.A1(new_n230), .A2(G20), .A3(G33), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n325), .B(KEYINPUT72), .ZN(new_n326));
  INV_X1    g0126(.A(G77), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n254), .A2(new_n327), .B1(new_n216), .B2(G68), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n246), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT11), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI211_X1 g0131(.A(KEYINPUT11), .B(new_n246), .C1(new_n326), .C2(new_n328), .ZN(new_n332));
  OAI21_X1  g0132(.A(KEYINPUT12), .B1(new_n264), .B2(G68), .ZN(new_n333));
  OR3_X1    g0133(.A1(new_n264), .A2(KEYINPUT12), .A3(G68), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n232), .B1(new_n263), .B2(G20), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n333), .A2(new_n334), .B1(new_n266), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n331), .A2(new_n332), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n222), .A2(G1698), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n289), .B(new_n338), .C1(G226), .C2(G1698), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n286), .A2(new_n239), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n278), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(G238), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n279), .B1(new_n343), .B2(new_n282), .ZN(new_n344));
  OAI21_X1  g0144(.A(KEYINPUT13), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n345), .A2(G190), .ZN(new_n346));
  INV_X1    g0146(.A(new_n342), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT13), .ZN(new_n348));
  INV_X1    g0148(.A(new_n344), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n337), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n350), .A2(KEYINPUT71), .A3(new_n345), .ZN(new_n352));
  OR4_X1    g0152(.A1(KEYINPUT71), .A2(new_n342), .A3(KEYINPUT13), .A4(new_n344), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n352), .A2(new_n353), .A3(G200), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n352), .A2(new_n353), .A3(G169), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT14), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT14), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n352), .A2(new_n353), .A3(new_n358), .A4(G169), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n350), .A2(G179), .A3(new_n345), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n357), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n355), .B1(new_n361), .B2(new_n337), .ZN(new_n362));
  INV_X1    g0162(.A(new_n246), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n264), .ZN(new_n364));
  OAI21_X1  g0164(.A(G77), .B1(new_n216), .B2(G1), .ZN(new_n365));
  OAI22_X1  g0165(.A1(new_n364), .A2(new_n365), .B1(G77), .B2(new_n264), .ZN(new_n366));
  XOR2_X1   g0166(.A(KEYINPUT8), .B(G58), .Z(new_n367));
  AOI22_X1  g0167(.A1(new_n367), .A2(new_n251), .B1(G20), .B2(G77), .ZN(new_n368));
  XNOR2_X1  g0168(.A(KEYINPUT15), .B(G87), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n368), .B1(new_n254), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n366), .B1(new_n370), .B2(new_n246), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n296), .A2(G238), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n289), .A2(G232), .A3(new_n290), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n372), .B(new_n373), .C1(new_n237), .C2(new_n289), .ZN(new_n374));
  INV_X1    g0174(.A(new_n278), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n280), .B1(G244), .B2(new_n283), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n371), .B1(new_n378), .B2(new_n321), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n376), .A2(new_n319), .A3(new_n377), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n376), .A2(G190), .A3(new_n377), .ZN(new_n383));
  INV_X1    g0183(.A(new_n371), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(G200), .B2(new_n378), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n382), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n362), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT17), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n253), .B1(new_n263), .B2(G20), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n389), .A2(new_n266), .B1(new_n253), .B2(new_n265), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT7), .B1(new_n299), .B2(new_n216), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n287), .A2(KEYINPUT7), .A3(new_n216), .A4(new_n288), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(G68), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G58), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n395), .A2(new_n232), .ZN(new_n396));
  OAI21_X1  g0196(.A(G20), .B1(new_n396), .B2(new_n247), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n251), .A2(G159), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(KEYINPUT16), .B1(new_n394), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n287), .A2(new_n216), .A3(new_n288), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT7), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n232), .B1(new_n404), .B2(new_n392), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n397), .A2(KEYINPUT16), .A3(new_n398), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n246), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n390), .B1(new_n401), .B2(new_n407), .ZN(new_n408));
  OR2_X1    g0208(.A1(G223), .A2(G1698), .ZN(new_n409));
  OAI221_X1 g0209(.A(new_n409), .B1(G226), .B2(new_n290), .C1(new_n297), .C2(new_n298), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G33), .A2(G87), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n278), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n279), .B1(new_n222), .B2(new_n282), .ZN(new_n413));
  OAI21_X1  g0213(.A(G200), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n410), .A2(new_n411), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n375), .ZN(new_n416));
  INV_X1    g0216(.A(new_n413), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n414), .B1(new_n418), .B2(new_n313), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n388), .B1(new_n408), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n416), .A2(G190), .A3(new_n417), .ZN(new_n421));
  AND2_X1   g0221(.A1(new_n421), .A2(new_n414), .ZN(new_n422));
  INV_X1    g0222(.A(new_n390), .ZN(new_n423));
  INV_X1    g0223(.A(new_n406), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n363), .B1(new_n394), .B2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT16), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(new_n405), .B2(new_n399), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n423), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n422), .A2(new_n428), .A3(KEYINPUT17), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n420), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT73), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n408), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n428), .A2(KEYINPUT73), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n418), .A2(G169), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n416), .A2(G179), .A3(new_n417), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n432), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n430), .B1(KEYINPUT18), .B2(new_n437), .ZN(new_n438));
  OR2_X1    g0238(.A1(new_n437), .A2(KEYINPUT18), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n324), .A2(new_n387), .A3(new_n440), .ZN(new_n441));
  OAI211_X1 g0241(.A(G257), .B(G1698), .C1(new_n297), .C2(new_n298), .ZN(new_n442));
  OAI211_X1 g0242(.A(G250), .B(new_n290), .C1(new_n297), .C2(new_n298), .ZN(new_n443));
  NAND2_X1  g0243(.A1(G33), .A2(G294), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n375), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT76), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT5), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n447), .B1(new_n448), .B2(G41), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n274), .A2(KEYINPUT76), .A3(KEYINPUT5), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n275), .A2(G1), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n448), .A2(G41), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n449), .A2(new_n450), .A3(new_n451), .A4(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n278), .A2(G274), .ZN(new_n454));
  OR2_X1    g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n453), .A2(G264), .A3(new_n278), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n446), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G169), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n446), .A2(G179), .A3(new_n455), .A4(new_n456), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT85), .ZN(new_n461));
  OR3_X1    g0261(.A1(new_n264), .A2(KEYINPUT25), .A3(G107), .ZN(new_n462));
  OAI21_X1  g0262(.A(KEYINPUT25), .B1(new_n264), .B2(G107), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n263), .A2(G33), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n264), .A2(new_n464), .A3(new_n215), .A4(new_n245), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n462), .B(new_n463), .C1(new_n237), .C2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT84), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n465), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G107), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n470), .A2(KEYINPUT84), .A3(new_n462), .A4(new_n463), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT23), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n473), .B1(new_n216), .B2(G107), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n237), .A2(KEYINPUT23), .A3(G20), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(G33), .A2(G116), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n216), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n216), .B(G87), .C1(new_n297), .C2(new_n298), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT22), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT22), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n289), .A2(new_n483), .A3(new_n216), .A4(G87), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n480), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  AND2_X1   g0285(.A1(new_n485), .A2(KEYINPUT24), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n246), .B1(new_n485), .B2(KEYINPUT24), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n472), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT85), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n458), .A2(new_n489), .A3(new_n459), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n461), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT86), .ZN(new_n492));
  OR2_X1    g0292(.A1(new_n485), .A2(KEYINPUT24), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n485), .A2(KEYINPUT24), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n493), .A2(new_n246), .A3(new_n494), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n446), .A2(new_n455), .A3(new_n456), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G190), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n457), .A2(G200), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n495), .A2(new_n472), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n491), .A2(new_n492), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n492), .B1(new_n491), .B2(new_n499), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g0302(.A(G264), .B(G1698), .C1(new_n297), .C2(new_n298), .ZN(new_n503));
  OAI211_X1 g0303(.A(G257), .B(new_n290), .C1(new_n297), .C2(new_n298), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n287), .A2(G303), .A3(new_n288), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n375), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n453), .A2(G270), .A3(new_n278), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n507), .A2(new_n455), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n469), .A2(G116), .ZN(new_n510));
  INV_X1    g0310(.A(G116), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n263), .A2(new_n511), .A3(G13), .A4(G20), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT82), .ZN(new_n513));
  XNOR2_X1  g0313(.A(new_n512), .B(new_n513), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n245), .A2(new_n215), .B1(G20), .B2(new_n511), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G33), .A2(G283), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n516), .B(new_n216), .C1(G33), .C2(new_n239), .ZN(new_n517));
  AND3_X1   g0317(.A1(new_n515), .A2(KEYINPUT20), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(KEYINPUT20), .B1(new_n515), .B2(new_n517), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n510), .B(new_n514), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n509), .A2(new_n520), .A3(G169), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT83), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT21), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n521), .A2(new_n522), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT21), .ZN(new_n526));
  INV_X1    g0326(.A(new_n520), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n507), .A2(G179), .A3(new_n455), .A4(new_n508), .ZN(new_n528));
  OR2_X1    g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n520), .B1(new_n509), .B2(G200), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(new_n313), .B2(new_n509), .ZN(new_n531));
  AND4_X1   g0331(.A1(new_n524), .A2(new_n526), .A3(new_n529), .A4(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n216), .A2(G33), .A3(G97), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT19), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(KEYINPUT78), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT78), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(KEYINPUT19), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n533), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT80), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT80), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n533), .A2(new_n535), .A3(new_n537), .A4(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n216), .B(G68), .C1(new_n297), .C2(new_n298), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n539), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n536), .A2(KEYINPUT19), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n534), .A2(KEYINPUT78), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n340), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(G97), .A2(G107), .ZN(new_n547));
  AND2_X1   g0347(.A1(KEYINPUT79), .A2(G87), .ZN(new_n548));
  NOR2_X1   g0348(.A1(KEYINPUT79), .A2(G87), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n546), .A2(new_n216), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n246), .B1(new_n543), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n369), .A2(new_n265), .ZN(new_n553));
  INV_X1    g0353(.A(new_n369), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n469), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n552), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n278), .A2(G274), .A3(new_n451), .ZN(new_n557));
  NOR2_X1   g0357(.A1(G238), .A2(G1698), .ZN(new_n558));
  INV_X1    g0358(.A(G244), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n558), .B1(new_n559), .B2(G1698), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n478), .B1(new_n560), .B2(new_n289), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n557), .B1(new_n561), .B2(new_n278), .ZN(new_n562));
  INV_X1    g0362(.A(G250), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n563), .B1(new_n263), .B2(G45), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT77), .ZN(new_n565));
  AND3_X1   g0365(.A1(new_n564), .A2(new_n278), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n565), .B1(new_n564), .B2(new_n278), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(G169), .B1(new_n562), .B2(new_n568), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n278), .A2(G274), .A3(new_n451), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n343), .A2(new_n290), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n559), .A2(G1698), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n571), .B(new_n572), .C1(new_n297), .C2(new_n298), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n477), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n570), .B1(new_n574), .B2(new_n375), .ZN(new_n575));
  INV_X1    g0375(.A(new_n567), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n564), .A2(new_n278), .A3(new_n565), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n575), .A2(G179), .A3(new_n578), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n556), .A2(KEYINPUT81), .B1(new_n569), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT81), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n552), .A2(new_n555), .A3(new_n581), .A4(new_n553), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n469), .A2(G87), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n552), .A2(new_n553), .A3(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(G200), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n585), .B1(new_n575), .B2(new_n578), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n562), .A2(new_n568), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n586), .B1(G190), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n580), .A2(new_n582), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n453), .A2(G257), .A3(new_n278), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n455), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n516), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n592), .B1(new_n296), .B2(G250), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT4), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n594), .A2(G1698), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n595), .B(G244), .C1(new_n298), .C2(new_n297), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT74), .ZN(new_n597));
  OAI211_X1 g0397(.A(G244), .B(new_n290), .C1(new_n297), .C2(new_n298), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n594), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT74), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n289), .A2(new_n600), .A3(G244), .A4(new_n595), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n593), .A2(new_n597), .A3(new_n599), .A4(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT75), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n278), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n597), .A2(new_n601), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n559), .B1(new_n287), .B2(new_n288), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT4), .B1(new_n606), .B2(new_n290), .ZN(new_n607));
  OAI211_X1 g0407(.A(G250), .B(G1698), .C1(new_n297), .C2(new_n298), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n516), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n605), .A2(new_n610), .A3(KEYINPUT75), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n591), .B1(new_n604), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n319), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n264), .A2(G97), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n465), .B2(new_n239), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT6), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n239), .A2(new_n237), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n617), .B1(new_n618), .B2(new_n547), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(new_n617), .B2(new_n238), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(G20), .ZN(new_n621));
  OAI21_X1  g0421(.A(G107), .B1(new_n391), .B2(new_n393), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n251), .A2(G77), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n616), .B1(new_n624), .B2(new_n246), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n613), .B(new_n626), .C1(G169), .C2(new_n612), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n612), .A2(G190), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n628), .B(new_n625), .C1(new_n585), .C2(new_n612), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n532), .A2(new_n589), .A3(new_n627), .A4(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n502), .A2(new_n630), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n441), .A2(new_n631), .ZN(G372));
  INV_X1    g0432(.A(new_n323), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n425), .A2(new_n427), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n634), .A2(new_n390), .B1(new_n434), .B2(new_n435), .ZN(new_n635));
  XNOR2_X1  g0435(.A(new_n635), .B(KEYINPUT18), .ZN(new_n636));
  INV_X1    g0436(.A(new_n355), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n637), .A2(new_n382), .B1(new_n361), .B2(new_n337), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n636), .B1(new_n638), .B2(new_n430), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n633), .B1(new_n639), .B2(new_n318), .ZN(new_n640));
  INV_X1    g0440(.A(new_n441), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n562), .A2(new_n319), .A3(new_n568), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n321), .B1(new_n575), .B2(new_n578), .ZN(new_n643));
  OAI21_X1  g0443(.A(KEYINPUT87), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT87), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n569), .A2(new_n645), .A3(new_n579), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n644), .A2(new_n556), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n588), .A2(new_n584), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n647), .A2(new_n499), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n488), .A2(new_n460), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n526), .A2(new_n650), .A3(new_n529), .A4(new_n524), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n649), .A2(new_n627), .A3(new_n629), .A4(new_n651), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n652), .A2(new_n647), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n602), .A2(new_n603), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n611), .A2(new_n654), .A3(new_n375), .ZN(new_n655));
  INV_X1    g0455(.A(new_n591), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n625), .B1(new_n657), .B2(new_n321), .ZN(new_n658));
  XNOR2_X1  g0458(.A(KEYINPUT88), .B(KEYINPUT26), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n589), .A2(new_n613), .A3(new_n658), .A4(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT89), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n658), .A2(new_n648), .A3(new_n613), .A4(new_n647), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n613), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n626), .B1(new_n612), .B2(G169), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n669), .A2(KEYINPUT89), .A3(new_n589), .A4(new_n660), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n663), .A2(new_n666), .A3(new_n670), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n653), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n640), .B1(new_n641), .B2(new_n672), .ZN(G369));
  NAND3_X1  g0473(.A1(new_n263), .A2(new_n216), .A3(G13), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(new_n676), .A3(G213), .ZN(new_n677));
  INV_X1    g0477(.A(G343), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n491), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n488), .A2(new_n679), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n500), .B2(new_n501), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT91), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OAI211_X1 g0485(.A(KEYINPUT91), .B(new_n682), .C1(new_n500), .C2(new_n501), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n681), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n526), .A2(new_n529), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n524), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n527), .A2(new_n680), .ZN(new_n690));
  MUX2_X1   g0490(.A(new_n532), .B(new_n689), .S(new_n690), .Z(new_n691));
  XOR2_X1   g0491(.A(KEYINPUT90), .B(G330), .Z(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n687), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n679), .B1(new_n688), .B2(new_n524), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n685), .A2(new_n686), .A3(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n488), .A2(new_n460), .A3(new_n680), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n695), .A2(new_n699), .ZN(G399));
  INV_X1    g0500(.A(new_n212), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(G41), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n550), .A2(new_n511), .A3(new_n547), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(new_n263), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n218), .B2(new_n703), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT28), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n679), .B1(new_n653), .B2(new_n671), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT29), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n556), .A2(KEYINPUT81), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n569), .A2(new_n579), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(new_n582), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n648), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n659), .B1(new_n627), .B2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT96), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT95), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n664), .B2(new_n665), .ZN(new_n720));
  OAI211_X1 g0520(.A(KEYINPUT96), .B(new_n659), .C1(new_n627), .C2(new_n715), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n647), .A2(new_n648), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n669), .A2(new_n722), .A3(KEYINPUT95), .A4(KEYINPUT26), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n718), .A2(new_n720), .A3(new_n721), .A4(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n647), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n649), .A2(new_n627), .A3(new_n629), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n688), .A2(new_n491), .A3(new_n524), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n679), .B1(new_n724), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n711), .B1(new_n710), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n496), .B1(new_n655), .B2(new_n656), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT92), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n732), .B1(new_n562), .B2(new_n568), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n575), .A2(KEYINPUT92), .A3(new_n578), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n733), .A2(new_n319), .A3(new_n509), .A4(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT93), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n455), .A2(new_n508), .ZN(new_n738));
  AOI21_X1  g0538(.A(G179), .B1(new_n738), .B2(new_n507), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n739), .A2(KEYINPUT93), .A3(new_n734), .A4(new_n733), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n731), .A2(new_n737), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n575), .A2(new_n578), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n446), .A2(new_n456), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n528), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n612), .A2(KEYINPUT30), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n612), .A2(new_n744), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT30), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n741), .A2(new_n745), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(KEYINPUT94), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT94), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n741), .A2(new_n748), .A3(new_n751), .A4(new_n745), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n750), .A2(new_n679), .A3(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT31), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n631), .A2(new_n680), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n749), .A2(KEYINPUT31), .A3(new_n679), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n692), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n730), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n708), .B1(new_n758), .B2(G1), .ZN(G364));
  INV_X1    g0559(.A(G13), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(G20), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n263), .B1(new_n761), .B2(G45), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n702), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n701), .A2(new_n299), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n766), .A2(G355), .B1(new_n511), .B2(new_n701), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n767), .A2(KEYINPUT97), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(KEYINPUT97), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n701), .A2(new_n289), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n219), .A2(new_n275), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n770), .B(new_n771), .C1(new_n275), .C2(new_n236), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n768), .A2(new_n769), .A3(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G13), .A2(G33), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(G20), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n215), .B1(G20), .B2(new_n321), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n778), .B(KEYINPUT98), .Z(new_n779));
  AND2_X1   g0579(.A1(new_n773), .A2(new_n779), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n313), .A2(G179), .A3(G200), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n216), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G97), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n216), .A2(new_n319), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n786), .A2(new_n585), .A3(G190), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n784), .B1(new_n788), .B2(new_n232), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n789), .B(KEYINPUT99), .Z(new_n790));
  NOR2_X1   g0590(.A1(new_n216), .A2(G179), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G190), .A2(G200), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G159), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT32), .ZN(new_n796));
  NOR3_X1   g0596(.A1(new_n786), .A2(new_n313), .A3(G200), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n395), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n785), .A2(new_n792), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n289), .B1(new_n800), .B2(new_n327), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n313), .A2(new_n585), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n785), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n791), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n803), .A2(new_n230), .B1(new_n804), .B2(new_n550), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n791), .A2(new_n313), .A3(G200), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(new_n237), .ZN(new_n807));
  NOR4_X1   g0607(.A1(new_n799), .A2(new_n801), .A3(new_n805), .A4(new_n807), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n790), .A2(new_n796), .A3(new_n808), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT100), .Z(new_n810));
  INV_X1    g0610(.A(new_n793), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G329), .ZN(new_n812));
  INV_X1    g0612(.A(G322), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n812), .B1(new_n798), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n803), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n814), .B1(G326), .B2(new_n815), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n804), .B(KEYINPUT101), .Z(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(G303), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n783), .A2(G294), .ZN(new_n819));
  INV_X1    g0619(.A(G283), .ZN(new_n820));
  INV_X1    g0620(.A(G311), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n820), .A2(new_n806), .B1(new_n800), .B2(new_n821), .ZN(new_n822));
  XNOR2_X1  g0622(.A(KEYINPUT33), .B(G317), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n289), .B(new_n822), .C1(new_n787), .C2(new_n823), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n816), .A2(new_n818), .A3(new_n819), .A4(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(KEYINPUT102), .B1(new_n810), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n777), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n810), .A2(KEYINPUT102), .A3(new_n825), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n765), .B(new_n780), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n776), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n830), .B1(new_n691), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n694), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n833), .A2(new_n764), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n693), .B2(new_n691), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(G396));
  NAND2_X1  g0637(.A1(new_n384), .A2(new_n679), .ZN(new_n838));
  OR3_X1    g0638(.A1(new_n381), .A2(KEYINPUT103), .A3(new_n680), .ZN(new_n839));
  OAI21_X1  g0639(.A(KEYINPUT103), .B1(new_n381), .B2(new_n680), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n386), .A2(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n709), .B(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n757), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n764), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n844), .B2(new_n843), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n827), .A2(new_n775), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n764), .B1(G77), .B2(new_n847), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n788), .A2(new_n820), .B1(new_n800), .B2(new_n511), .ZN(new_n849));
  INV_X1    g0649(.A(new_n806), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n289), .B(new_n849), .C1(G87), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n817), .A2(G107), .ZN(new_n852));
  INV_X1    g0652(.A(G303), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n803), .A2(new_n853), .B1(new_n793), .B2(new_n821), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(G294), .B2(new_n797), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n851), .A2(new_n784), .A3(new_n852), .A4(new_n855), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n787), .A2(G150), .B1(new_n815), .B2(G137), .ZN(new_n857));
  INV_X1    g0657(.A(G143), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n857), .B1(new_n858), .B2(new_n798), .C1(new_n794), .C2(new_n800), .ZN(new_n859));
  XOR2_X1   g0659(.A(new_n859), .B(KEYINPUT34), .Z(new_n860));
  NOR2_X1   g0660(.A1(new_n806), .A2(new_n232), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n299), .B(new_n861), .C1(G132), .C2(new_n811), .ZN(new_n862));
  INV_X1    g0662(.A(new_n817), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n862), .B1(new_n395), .B2(new_n782), .C1(new_n863), .C2(new_n230), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n856), .B1(new_n860), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n848), .B1(new_n865), .B2(new_n777), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n842), .B2(new_n775), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n846), .A2(new_n867), .ZN(G384));
  NOR2_X1   g0668(.A1(new_n761), .A2(new_n263), .ZN(new_n869));
  INV_X1    g0669(.A(new_n677), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n432), .A2(new_n433), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT37), .B1(new_n422), .B2(new_n428), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n437), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT105), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n437), .A2(new_n871), .A3(KEYINPUT105), .A4(new_n872), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT104), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n408), .A2(new_n419), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n878), .B1(new_n635), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n436), .A2(new_n408), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n422), .A2(new_n428), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n881), .A2(new_n882), .A3(KEYINPUT104), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n408), .A2(new_n870), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n880), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(KEYINPUT37), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n877), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n884), .B1(new_n438), .B2(new_n439), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n887), .A2(KEYINPUT38), .A3(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT38), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n875), .A2(new_n876), .B1(new_n885), .B2(KEYINPUT37), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n891), .B1(new_n892), .B2(new_n888), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n337), .A2(new_n679), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n362), .A2(new_n896), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n337), .B(new_n679), .C1(new_n361), .C2(new_n355), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI211_X1 g0699(.A(new_n679), .B(new_n841), .C1(new_n653), .C2(new_n671), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n381), .A2(new_n679), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n894), .B(new_n899), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n636), .A2(new_n870), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT38), .B1(new_n887), .B2(new_n889), .ZN(new_n905));
  NOR3_X1   g0705(.A1(new_n892), .A2(new_n891), .A3(new_n888), .ZN(new_n906));
  OAI21_X1  g0706(.A(KEYINPUT39), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(KEYINPUT106), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT107), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n635), .B2(new_n879), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n881), .A2(new_n882), .A3(KEYINPUT107), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n910), .A2(new_n871), .A3(new_n911), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n875), .A2(new_n876), .B1(new_n912), .B2(KEYINPUT37), .ZN(new_n913));
  INV_X1    g0713(.A(new_n430), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n871), .B1(new_n636), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n891), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT39), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n890), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT106), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n919), .B(KEYINPUT39), .C1(new_n905), .C2(new_n906), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n908), .A2(new_n918), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n361), .A2(new_n337), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n922), .A2(new_n679), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n904), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n730), .A2(new_n441), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n640), .ZN(new_n926));
  XOR2_X1   g0726(.A(new_n924), .B(new_n926), .Z(new_n927));
  NAND2_X1  g0727(.A1(new_n890), .A2(new_n916), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n753), .A2(new_n754), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n491), .A2(new_n499), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(KEYINPUT86), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n491), .A2(new_n492), .A3(new_n499), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AND3_X1   g0733(.A1(new_n627), .A2(new_n629), .A3(new_n589), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n933), .A2(new_n934), .A3(new_n532), .A4(new_n680), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n750), .A2(KEYINPUT31), .A3(new_n679), .A4(new_n752), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n929), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n898), .ZN(new_n938));
  AOI211_X1 g0738(.A(new_n895), .B(new_n355), .C1(new_n361), .C2(new_n337), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n842), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n928), .A2(new_n937), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n940), .B1(new_n755), .B2(new_n936), .ZN(new_n943));
  AOI21_X1  g0743(.A(KEYINPUT40), .B1(new_n890), .B2(new_n893), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n942), .A2(KEYINPUT40), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n441), .A2(new_n937), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n945), .B(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n947), .A2(new_n692), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n869), .B1(new_n927), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n927), .B2(new_n949), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n620), .A2(KEYINPUT35), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n620), .A2(KEYINPUT35), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n952), .A2(G116), .A3(new_n217), .A4(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT36), .ZN(new_n955));
  OAI21_X1  g0755(.A(G77), .B1(new_n395), .B2(new_n232), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n231), .B1(new_n956), .B2(new_n218), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n957), .A2(G1), .A3(new_n760), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n951), .A2(new_n955), .A3(new_n958), .ZN(G367));
  INV_X1    g0759(.A(new_n695), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n627), .B(new_n629), .C1(new_n625), .C2(new_n680), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n669), .A2(new_n679), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n960), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n685), .A2(new_n963), .A3(new_n686), .A4(new_n696), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n967), .A2(KEYINPUT42), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n627), .B1(new_n961), .B2(new_n491), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n967), .A2(KEYINPUT42), .B1(new_n680), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(KEYINPUT108), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n584), .A2(new_n680), .ZN(new_n973));
  MUX2_X1   g0773(.A(new_n722), .B(new_n725), .S(new_n973), .Z(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT43), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT108), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n968), .A2(new_n970), .A3(new_n976), .ZN(new_n977));
  AND3_X1   g0777(.A1(new_n972), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(new_n972), .B2(new_n977), .ZN(new_n980));
  NOR3_X1   g0780(.A1(new_n978), .A2(new_n980), .A3(KEYINPUT109), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT109), .ZN(new_n982));
  INV_X1    g0782(.A(new_n977), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n976), .B1(new_n968), .B2(new_n970), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n983), .A2(new_n984), .B1(KEYINPUT43), .B2(new_n974), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n972), .A2(new_n975), .A3(new_n977), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n982), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n966), .B1(new_n981), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(KEYINPUT109), .B1(new_n978), .B2(new_n980), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n985), .A2(new_n982), .A3(new_n986), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n989), .A2(new_n965), .A3(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n702), .B(KEYINPUT41), .Z(new_n992));
  NAND3_X1  g0792(.A1(new_n697), .A2(new_n698), .A3(new_n963), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT45), .ZN(new_n994));
  AND2_X1   g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n993), .A2(new_n994), .ZN(new_n996));
  AOI21_X1  g0796(.A(KEYINPUT44), .B1(new_n699), .B2(new_n964), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT44), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n998), .B(new_n963), .C1(new_n697), .C2(new_n698), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n995), .A2(new_n996), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n1000), .A2(KEYINPUT110), .A3(new_n695), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n681), .B(new_n696), .C1(new_n685), .C2(new_n686), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n697), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n833), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n696), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n687), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1006), .A2(new_n694), .A3(new_n697), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n758), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n960), .B1(new_n997), .B2(new_n999), .C1(new_n996), .C2(new_n995), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n695), .A2(KEYINPUT110), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1001), .A2(new_n1010), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n992), .B1(new_n1013), .B2(new_n758), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n988), .B(new_n991), .C1(new_n1014), .C2(new_n763), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n770), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1016), .A2(new_n228), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n778), .B1(new_n212), .B2(new_n369), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n764), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n800), .A2(new_n230), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n788), .A2(new_n794), .B1(new_n804), .B2(new_n395), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n1020), .B(new_n1021), .C1(G137), .C2(new_n811), .ZN(new_n1022));
  INV_X1    g0822(.A(G150), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n798), .A2(new_n1023), .B1(new_n803), .B2(new_n858), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(G68), .B2(new_n783), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n850), .A2(G77), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n289), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1027), .A2(KEYINPUT113), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(KEYINPUT113), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1022), .A2(new_n1025), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(G294), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(KEYINPUT112), .B(G317), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n788), .A2(new_n1031), .B1(new_n793), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(G97), .B2(new_n850), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n817), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n797), .A2(G303), .B1(new_n815), .B2(G311), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1036), .A2(KEYINPUT111), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(KEYINPUT111), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1034), .A2(new_n1035), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n800), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n289), .B1(new_n1040), .B2(G283), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n804), .A2(new_n511), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1041), .B1(KEYINPUT46), .B2(new_n1042), .C1(new_n237), .C2(new_n782), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1030), .B1(new_n1039), .B2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT47), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1019), .B1(new_n1045), .B2(new_n777), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n974), .B2(new_n831), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1015), .A2(new_n1047), .ZN(G387));
  NAND2_X1  g0848(.A1(new_n1009), .A2(new_n702), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT114), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n758), .A2(new_n1008), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1009), .A2(KEYINPUT114), .A3(new_n702), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n804), .A2(new_n327), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n289), .B1(new_n806), .B2(new_n239), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n1055), .B(new_n1056), .C1(G68), .C2(new_n1040), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n815), .A2(G159), .B1(new_n811), .B2(G150), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n367), .A2(new_n787), .B1(new_n797), .B2(G50), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n783), .A2(new_n554), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n787), .A2(G311), .B1(G303), .B2(new_n1040), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1062), .B1(new_n813), .B2(new_n803), .C1(new_n798), .C2(new_n1032), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT48), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n782), .A2(new_n820), .B1(new_n804), .B2(new_n1031), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1065), .A2(KEYINPUT49), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n289), .B1(new_n811), .B2(G326), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1068), .B(new_n1069), .C1(new_n511), .C2(new_n806), .ZN(new_n1070));
  AOI21_X1  g0870(.A(KEYINPUT49), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1061), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n777), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n225), .A2(new_n275), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n1074), .A2(new_n770), .B1(new_n704), .B2(new_n766), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n367), .A2(new_n230), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT50), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n275), .B1(new_n232), .B2(new_n327), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n1077), .A2(new_n704), .A3(new_n1078), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n1075), .A2(new_n1079), .B1(G107), .B2(new_n212), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n765), .B1(new_n1080), .B2(new_n779), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1073), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n687), .B2(new_n776), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n1008), .B2(new_n763), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1054), .A2(new_n1084), .ZN(G393));
  NAND2_X1  g0885(.A1(new_n1000), .A2(new_n695), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT115), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1086), .A2(new_n1011), .A3(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1000), .A2(KEYINPUT115), .A3(new_n695), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n762), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n964), .A2(new_n776), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n778), .B1(new_n239), .B2(new_n212), .C1(new_n1016), .C2(new_n243), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n764), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n788), .A2(new_n230), .B1(new_n793), .B2(new_n858), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n299), .B1(new_n850), .B2(G87), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n327), .B2(new_n782), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n232), .A2(new_n804), .B1(new_n800), .B2(new_n253), .ZN(new_n1097));
  OR3_X1    g0897(.A1(new_n1094), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n797), .A2(G159), .B1(new_n815), .B2(G150), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT51), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n797), .A2(G311), .B1(new_n815), .B2(G317), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT52), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n289), .B(new_n807), .C1(G116), .C2(new_n783), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n804), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(G283), .A2(new_n1104), .B1(new_n811), .B2(G322), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n787), .A2(G303), .B1(G294), .B2(new_n1040), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1103), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n1098), .A2(new_n1100), .B1(new_n1102), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1093), .B1(new_n1108), .B2(new_n777), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1091), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  OR3_X1    g0911(.A1(new_n1090), .A2(KEYINPUT116), .A3(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(KEYINPUT116), .B1(new_n1090), .B2(new_n1111), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1088), .A2(new_n1009), .A3(new_n1089), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1115), .A2(new_n702), .A3(new_n1013), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1114), .A2(new_n1116), .ZN(G390));
  INV_X1    g0917(.A(new_n923), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n901), .B1(new_n709), .B2(new_n842), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n899), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1118), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1121), .A2(new_n908), .A3(new_n918), .A4(new_n920), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n901), .B1(new_n729), .B2(new_n842), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1118), .B(new_n928), .C1(new_n1123), .C2(new_n1120), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n929), .A2(new_n935), .A3(new_n756), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1125), .A2(new_n693), .A3(new_n842), .A4(new_n899), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1122), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n928), .A2(new_n1118), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n729), .A2(new_n842), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n901), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1128), .B1(new_n1131), .B2(new_n899), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n920), .A2(new_n918), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n919), .B1(new_n894), .B2(KEYINPUT39), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1132), .B1(new_n1135), .B2(new_n1121), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n941), .A2(G330), .A3(new_n937), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1127), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n441), .A2(G330), .A3(new_n937), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n925), .A2(new_n640), .A3(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n937), .A2(G330), .A3(new_n842), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n1141), .A2(KEYINPUT117), .A3(new_n1120), .ZN(new_n1142));
  AOI21_X1  g0942(.A(KEYINPUT117), .B1(new_n1141), .B2(new_n1120), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1125), .A2(new_n693), .A3(new_n842), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n1120), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1119), .B1(new_n1147), .B2(new_n1137), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1140), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1138), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1137), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1141), .A2(new_n1120), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT117), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1141), .A2(KEYINPUT117), .A3(new_n1120), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1147), .A2(new_n1137), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1119), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1159), .A2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1153), .A2(new_n1127), .A3(new_n1163), .A4(new_n1140), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1150), .A2(new_n702), .A3(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n921), .A2(new_n775), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n289), .B1(new_n817), .B2(G87), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT119), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n861), .B1(new_n787), .B2(G107), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n327), .B2(new_n782), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n798), .A2(new_n511), .B1(new_n800), .B2(new_n239), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n803), .A2(new_n820), .B1(new_n793), .B2(new_n1031), .ZN(new_n1172));
  NOR3_X1   g0972(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n797), .A2(G132), .B1(new_n815), .B2(G128), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1174), .B(KEYINPUT118), .Z(new_n1175));
  AOI22_X1  g0975(.A1(new_n787), .A2(G137), .B1(G125), .B2(new_n811), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n230), .B2(new_n806), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(KEYINPUT54), .B(G143), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n804), .A2(new_n1023), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT53), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n289), .B1(new_n800), .B2(new_n1178), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n794), .B2(new_n782), .ZN(new_n1183));
  NOR3_X1   g0983(.A1(new_n1177), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n1168), .A2(new_n1173), .B1(new_n1175), .B2(new_n1184), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n764), .B1(new_n367), .B2(new_n847), .C1(new_n1185), .C2(new_n827), .ZN(new_n1186));
  OAI21_X1  g0986(.A(KEYINPUT120), .B1(new_n1166), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1186), .B1(new_n1135), .B2(new_n774), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT120), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1187), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1153), .A2(new_n763), .A3(new_n1127), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1165), .A2(new_n1193), .ZN(G378));
  OAI21_X1  g0994(.A(new_n1140), .B1(new_n1138), .B2(new_n1149), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n269), .A2(new_n870), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(new_n318), .B2(new_n323), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n318), .A2(new_n323), .A3(new_n1196), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1200), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1196), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n633), .B(new_n1203), .C1(new_n315), .C2(new_n317), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1202), .B1(new_n1197), .B2(new_n1204), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n1201), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(G330), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1206), .B1(new_n945), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1201), .A2(new_n1205), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT40), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n943), .B2(new_n928), .ZN(new_n1211));
  AND4_X1   g1011(.A1(new_n1210), .A2(new_n894), .A3(new_n937), .A4(new_n941), .ZN(new_n1212));
  OAI211_X1 g1012(.A(G330), .B(new_n1209), .C1(new_n1211), .C2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1208), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n924), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n924), .A2(new_n1208), .A3(new_n1213), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1195), .A2(KEYINPUT57), .A3(new_n1218), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1195), .A2(new_n1218), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n702), .B(new_n1219), .C1(new_n1220), .C2(KEYINPUT57), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1206), .A2(new_n774), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n764), .B1(G50), .B2(new_n847), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n230), .B1(G33), .B2(G41), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n299), .B2(new_n274), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n798), .A2(new_n237), .B1(new_n369), .B2(new_n800), .ZN(new_n1226));
  NOR4_X1   g1026(.A1(new_n1226), .A2(G41), .A3(new_n289), .A4(new_n1055), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n803), .A2(new_n511), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n806), .A2(new_n395), .B1(new_n793), .B2(new_n820), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1228), .B(new_n1229), .C1(G97), .C2(new_n787), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1227), .B(new_n1230), .C1(new_n232), .C2(new_n782), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT58), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1225), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(KEYINPUT122), .B(G124), .ZN(new_n1234));
  AOI211_X1 g1034(.A(G33), .B(G41), .C1(new_n811), .C2(new_n1234), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n787), .A2(G132), .B1(G137), .B2(new_n1040), .ZN(new_n1236));
  INV_X1    g1036(.A(G125), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1236), .B1(new_n1237), .B2(new_n803), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n804), .A2(new_n1178), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(new_n797), .B2(G128), .ZN(new_n1240));
  XOR2_X1   g1040(.A(new_n1240), .B(KEYINPUT121), .Z(new_n1241));
  AOI211_X1 g1041(.A(new_n1238), .B(new_n1241), .C1(G150), .C2(new_n783), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT59), .ZN(new_n1243));
  OAI221_X1 g1043(.A(new_n1235), .B1(new_n794), .B2(new_n806), .C1(new_n1242), .C2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  OAI221_X1 g1046(.A(new_n1233), .B1(new_n1232), .B2(new_n1231), .C1(new_n1244), .C2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1223), .B1(new_n1247), .B2(new_n777), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n1218), .A2(new_n763), .B1(new_n1222), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1221), .A2(new_n1249), .ZN(G375));
  NAND2_X1  g1050(.A1(new_n1120), .A2(new_n774), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n764), .B1(G68), .B2(new_n847), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(G150), .A2(new_n1040), .B1(new_n811), .B2(G128), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n299), .B1(new_n850), .B2(G58), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1253), .B(new_n1254), .C1(new_n230), .C2(new_n782), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n797), .A2(G137), .B1(new_n815), .B2(G132), .ZN(new_n1256));
  OAI221_X1 g1056(.A(new_n1256), .B1(new_n788), .B2(new_n1178), .C1(new_n863), .C2(new_n794), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(G116), .A2(new_n787), .B1(new_n797), .B2(G283), .ZN(new_n1258));
  OAI221_X1 g1058(.A(new_n1258), .B1(new_n1031), .B2(new_n803), .C1(new_n863), .C2(new_n239), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(G107), .A2(new_n1040), .B1(new_n811), .B2(G303), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1260), .A2(new_n299), .A3(new_n1060), .A4(new_n1026), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n1255), .A2(new_n1257), .B1(new_n1259), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT123), .ZN(new_n1263));
  OR2_X1    g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n827), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1252), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n1163), .A2(new_n763), .B1(new_n1251), .B2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n992), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1149), .A2(new_n1268), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1163), .A2(new_n1140), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1267), .B1(new_n1269), .B2(new_n1270), .ZN(G381));
  AND2_X1   g1071(.A1(new_n1221), .A2(new_n1249), .ZN(new_n1272));
  INV_X1    g1072(.A(G387), .ZN(new_n1273));
  INV_X1    g1073(.A(G390), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1054), .A2(new_n836), .A3(new_n1084), .ZN(new_n1275));
  NOR4_X1   g1075(.A1(G378), .A2(G381), .A3(G384), .A4(new_n1275), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1272), .A2(new_n1273), .A3(new_n1274), .A4(new_n1276), .ZN(G407));
  INV_X1    g1077(.A(G213), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(G378), .A2(G343), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1278), .B1(new_n1272), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(G407), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1281), .B(KEYINPUT124), .ZN(G409));
  NAND3_X1  g1082(.A1(new_n925), .A2(new_n640), .A3(new_n1139), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1159), .A2(new_n1162), .A3(new_n1283), .A4(KEYINPUT60), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1149), .A2(new_n1284), .A3(new_n702), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1148), .B1(new_n1286), .B2(new_n1156), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT60), .B1(new_n1287), .B2(new_n1283), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1267), .B1(new_n1285), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(G384), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  OAI211_X1 g1091(.A(G384), .B(new_n1267), .C1(new_n1285), .C2(new_n1288), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1278), .A2(G343), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  OR2_X1    g1094(.A1(new_n1294), .A2(KEYINPUT125), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1291), .A2(new_n1292), .A3(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1293), .A2(G2897), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1296), .A2(new_n1298), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1291), .A2(new_n1292), .A3(new_n1297), .A4(new_n1295), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1122), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1137), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1283), .B1(new_n1305), .B2(new_n1163), .ZN(new_n1306));
  AND3_X1   g1106(.A1(new_n924), .A2(new_n1208), .A3(new_n1213), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n921), .A2(new_n923), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n904), .ZN(new_n1309));
  AOI22_X1  g1109(.A1(new_n1208), .A2(new_n1213), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  OAI21_X1  g1110(.A(KEYINPUT57), .B1(new_n1307), .B2(new_n1310), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n702), .B1(new_n1306), .B2(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(KEYINPUT57), .B1(new_n1195), .B2(new_n1218), .ZN(new_n1313));
  OAI211_X1 g1113(.A(G378), .B(new_n1249), .C1(new_n1312), .C2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1195), .A2(new_n1268), .A3(new_n1218), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(new_n1249), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n703), .B1(new_n1138), .B2(new_n1149), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1317), .B1(new_n1164), .B2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1316), .A2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1314), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n1294), .ZN(new_n1322));
  AOI21_X1  g1122(.A(KEYINPUT61), .B1(new_n1302), .B2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT63), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1324), .B1(new_n1322), .B2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1275), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n836), .B1(new_n1054), .B2(new_n1084), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1329), .B1(G387), .B2(KEYINPUT126), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(G393), .A2(G396), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(new_n1275), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1332), .B1(new_n1047), .B2(new_n1015), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1274), .B1(new_n1330), .B2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(G387), .A2(new_n1329), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT126), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1336), .B1(new_n1015), .B2(new_n1047), .ZN(new_n1337));
  OAI211_X1 g1137(.A(new_n1335), .B(G390), .C1(new_n1329), .C2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1334), .A2(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1293), .B1(new_n1314), .B2(new_n1320), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1325), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1340), .A2(KEYINPUT63), .A3(new_n1341), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1323), .A2(new_n1326), .A3(new_n1339), .A4(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT62), .ZN(new_n1344));
  AND3_X1   g1144(.A1(new_n1340), .A2(new_n1344), .A3(new_n1341), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT61), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1346), .B1(new_n1340), .B2(new_n1301), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1344), .B1(new_n1340), .B2(new_n1341), .ZN(new_n1348));
  NOR3_X1   g1148(.A1(new_n1345), .A2(new_n1347), .A3(new_n1348), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1343), .B1(new_n1349), .B2(new_n1339), .ZN(G405));
  NAND2_X1  g1150(.A1(new_n1339), .A2(KEYINPUT127), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(G375), .A2(new_n1319), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1352), .A2(new_n1325), .A3(new_n1314), .ZN(new_n1353));
  AOI21_X1  g1153(.A(G378), .B1(new_n1221), .B2(new_n1249), .ZN(new_n1354));
  INV_X1    g1154(.A(new_n1314), .ZN(new_n1355));
  OAI21_X1  g1155(.A(new_n1341), .B1(new_n1354), .B2(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1353), .A2(new_n1356), .ZN(new_n1357));
  INV_X1    g1157(.A(KEYINPUT127), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1334), .A2(new_n1338), .A3(new_n1358), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1351), .A2(new_n1357), .A3(new_n1359), .ZN(new_n1360));
  NAND4_X1  g1160(.A1(new_n1339), .A2(new_n1353), .A3(KEYINPUT127), .A4(new_n1356), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1360), .A2(new_n1361), .ZN(G402));
endmodule


