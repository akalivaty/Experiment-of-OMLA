//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 1 1 0 1 0 1 1 0 1 1 0 0 1 1 1 1 1 1 0 0 0 1 0 1 0 1 0 1 0 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n777, new_n778,
    new_n779, new_n780, new_n782, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n860, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n984, new_n985, new_n986;
  XNOR2_X1  g000(.A(KEYINPUT77), .B(G211gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G218gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT76), .B(KEYINPUT22), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G197gat), .B(G204gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n205), .A2(new_n206), .A3(new_n208), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT78), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT78), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n210), .A2(new_n214), .A3(new_n211), .ZN(new_n215));
  NOR2_X1   g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XOR2_X1   g018(.A(G141gat), .B(G148gat), .Z(new_n220));
  INV_X1    g019(.A(KEYINPUT2), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT80), .ZN(new_n223));
  INV_X1    g022(.A(G141gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(KEYINPUT80), .A2(G141gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(G148gat), .A3(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT81), .B1(new_n224), .B2(G148gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n225), .A2(KEYINPUT81), .A3(G148gat), .A4(new_n226), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n218), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n232), .B1(new_n221), .B2(new_n216), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n222), .B1(new_n231), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  XOR2_X1   g036(.A(KEYINPUT79), .B(KEYINPUT29), .Z(new_n238));
  AOI22_X1  g037(.A1(new_n213), .A2(new_n215), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G228gat), .A2(G233gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT87), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n210), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n207), .A2(KEYINPUT87), .A3(new_n209), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n243), .A2(new_n211), .A3(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT3), .B1(new_n245), .B2(new_n238), .ZN(new_n246));
  OAI211_X1 g045(.A(new_n240), .B(new_n241), .C1(new_n246), .C2(new_n235), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT29), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n212), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n235), .B1(new_n249), .B2(new_n236), .ZN(new_n250));
  OAI211_X1 g049(.A(G228gat), .B(G233gat), .C1(new_n239), .C2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(G22gat), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT86), .ZN(new_n254));
  INV_X1    g053(.A(G22gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n247), .A2(new_n251), .A3(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n253), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G78gat), .B(G106gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT31), .B(G50gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(KEYINPUT88), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n257), .A2(new_n262), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n253), .A2(new_n254), .A3(new_n256), .A4(new_n261), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(G183gat), .A2(G190gat), .ZN(new_n268));
  MUX2_X1   g067(.A(KEYINPUT24), .B(new_n267), .S(new_n268), .Z(new_n269));
  NOR2_X1   g068(.A1(G169gat), .A2(G176gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT23), .ZN(new_n271));
  OR2_X1    g070(.A1(new_n270), .A2(KEYINPUT23), .ZN(new_n272));
  NAND2_X1  g071(.A1(G169gat), .A2(G176gat), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n269), .A2(new_n271), .A3(new_n272), .A4(new_n273), .ZN(new_n274));
  XOR2_X1   g073(.A(KEYINPUT65), .B(KEYINPUT25), .Z(new_n275));
  NAND2_X1  g074(.A1(new_n272), .A2(KEYINPUT25), .ZN(new_n276));
  INV_X1    g075(.A(new_n273), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n271), .B1(new_n277), .B2(KEYINPUT66), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT66), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n273), .A2(new_n279), .ZN(new_n280));
  NOR3_X1   g079(.A1(new_n276), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  AOI22_X1  g080(.A1(new_n274), .A2(new_n275), .B1(new_n281), .B2(new_n269), .ZN(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT27), .B(G183gat), .ZN(new_n283));
  INV_X1    g082(.A(G190gat), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(KEYINPUT28), .A3(new_n284), .ZN(new_n285));
  AND2_X1   g084(.A1(KEYINPUT67), .A2(KEYINPUT27), .ZN(new_n286));
  NOR2_X1   g085(.A1(KEYINPUT67), .A2(KEYINPUT27), .ZN(new_n287));
  OAI21_X1  g086(.A(G183gat), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT68), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT68), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n290), .B(G183gat), .C1(new_n286), .C2(new_n287), .ZN(new_n291));
  INV_X1    g090(.A(G183gat), .ZN(new_n292));
  AOI21_X1  g091(.A(G190gat), .B1(new_n292), .B2(KEYINPUT27), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n289), .A2(KEYINPUT69), .A3(new_n291), .A4(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT28), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n293), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n297), .B1(new_n288), .B2(KEYINPUT68), .ZN(new_n298));
  AOI21_X1  g097(.A(KEYINPUT69), .B1(new_n298), .B2(new_n291), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n285), .B1(new_n296), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n270), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n277), .B1(new_n301), .B2(KEYINPUT26), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT70), .ZN(new_n303));
  OR2_X1    g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(KEYINPUT71), .B(KEYINPUT26), .ZN(new_n305));
  AOI22_X1  g104(.A1(new_n302), .A2(new_n303), .B1(new_n305), .B2(new_n270), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  AND2_X1   g106(.A1(new_n307), .A2(new_n268), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n282), .B1(new_n300), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(G113gat), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n310), .A2(KEYINPUT72), .A3(G120gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT72), .ZN(new_n312));
  INV_X1    g111(.A(G120gat), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n312), .B1(G113gat), .B2(new_n313), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n313), .A2(G113gat), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n311), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G134gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G127gat), .ZN(new_n318));
  INV_X1    g117(.A(G127gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G134gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT1), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n318), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n310), .A2(G120gat), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n321), .B1(new_n324), .B2(new_n315), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n318), .A2(new_n320), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n316), .A2(new_n323), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n309), .B(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G227gat), .A2(G233gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT34), .ZN(new_n332));
  XOR2_X1   g131(.A(new_n330), .B(KEYINPUT64), .Z(new_n333));
  OR3_X1    g132(.A1(new_n328), .A2(KEYINPUT34), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT32), .ZN(new_n336));
  AND2_X1   g135(.A1(new_n328), .A2(new_n333), .ZN(new_n337));
  XOR2_X1   g136(.A(G15gat), .B(G43gat), .Z(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(KEYINPUT73), .ZN(new_n339));
  XOR2_X1   g138(.A(G71gat), .B(G99gat), .Z(new_n340));
  XNOR2_X1  g139(.A(new_n340), .B(KEYINPUT74), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n339), .B(new_n341), .ZN(new_n342));
  AOI211_X1 g141(.A(new_n336), .B(new_n337), .C1(KEYINPUT33), .C2(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n342), .B1(new_n337), .B2(KEYINPUT33), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n337), .A2(new_n336), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n335), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  AND2_X1   g146(.A1(new_n332), .A2(new_n334), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n344), .A2(new_n345), .ZN(new_n349));
  INV_X1    g148(.A(new_n333), .ZN(new_n350));
  OAI21_X1  g149(.A(KEYINPUT32), .B1(new_n329), .B2(new_n350), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n351), .B(new_n342), .C1(KEYINPUT33), .C2(new_n337), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n348), .A2(new_n349), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n266), .A2(new_n347), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT5), .ZN(new_n355));
  NAND2_X1  g154(.A1(G225gat), .A2(G233gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G113gat), .B(G120gat), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n326), .B1(new_n358), .B2(KEYINPUT1), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n310), .A2(KEYINPUT72), .A3(G120gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n315), .ZN(new_n361));
  OAI21_X1  g160(.A(KEYINPUT72), .B1(new_n310), .B2(G120gat), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n359), .B1(new_n363), .B2(new_n322), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n233), .B1(new_n229), .B2(new_n230), .ZN(new_n365));
  NOR3_X1   g164(.A1(new_n364), .A2(new_n365), .A3(new_n222), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT81), .ZN(new_n367));
  INV_X1    g166(.A(G148gat), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n367), .B1(G141gat), .B2(new_n368), .ZN(new_n369));
  AND2_X1   g168(.A1(KEYINPUT80), .A2(G141gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(KEYINPUT80), .A2(G141gat), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n369), .B1(new_n372), .B2(G148gat), .ZN(new_n373));
  INV_X1    g172(.A(new_n230), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n234), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n222), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n316), .A2(new_n323), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n375), .A2(new_n376), .B1(new_n359), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n357), .B1(new_n366), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n355), .B1(new_n379), .B2(KEYINPUT83), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n375), .A2(new_n327), .A3(new_n376), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n364), .B1(new_n365), .B2(new_n222), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n356), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT83), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT4), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n375), .A2(new_n327), .A3(new_n376), .A4(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT82), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n389), .B1(new_n366), .B2(new_n386), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n381), .A2(KEYINPUT82), .A3(KEYINPUT4), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n388), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n364), .B1(new_n235), .B2(new_n236), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n375), .A2(new_n376), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n394), .A2(KEYINPUT3), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n356), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n380), .B(new_n385), .C1(new_n392), .C2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n387), .A2(KEYINPUT84), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT84), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n235), .A2(new_n399), .A3(new_n386), .A4(new_n327), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n381), .A2(KEYINPUT4), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n327), .B1(new_n394), .B2(KEYINPUT3), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n237), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n357), .A2(KEYINPUT5), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n403), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n397), .A2(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(G1gat), .B(G29gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(KEYINPUT0), .ZN(new_n410));
  XNOR2_X1  g209(.A(G57gat), .B(G85gat), .ZN(new_n411));
  XOR2_X1   g210(.A(new_n410), .B(new_n411), .Z(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n414), .A2(KEYINPUT6), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT6), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT85), .ZN(new_n417));
  OAI21_X1  g216(.A(KEYINPUT5), .B1(new_n383), .B2(new_n384), .ZN(new_n418));
  AOI211_X1 g217(.A(KEYINPUT83), .B(new_n356), .C1(new_n381), .C2(new_n382), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n381), .A2(KEYINPUT82), .A3(KEYINPUT4), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT82), .B1(new_n381), .B2(KEYINPUT4), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n387), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n357), .B1(new_n404), .B2(new_n237), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI22_X1  g224(.A1(new_n401), .A2(new_n402), .B1(new_n237), .B2(new_n404), .ZN(new_n426));
  AOI22_X1  g225(.A1(new_n420), .A2(new_n425), .B1(new_n426), .B2(new_n406), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n417), .B1(new_n427), .B2(new_n412), .ZN(new_n428));
  AND4_X1   g227(.A1(new_n417), .A2(new_n397), .A3(new_n412), .A4(new_n407), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n416), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n415), .B1(new_n430), .B2(new_n414), .ZN(new_n431));
  NAND2_X1  g230(.A1(G226gat), .A2(G233gat), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n432), .B1(new_n309), .B2(KEYINPUT29), .ZN(new_n433));
  INV_X1    g232(.A(new_n432), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n307), .A2(new_n268), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n298), .A2(new_n291), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT69), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n438), .A2(new_n295), .A3(new_n294), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n435), .B1(new_n439), .B2(new_n285), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n434), .B1(new_n440), .B2(new_n282), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n213), .A2(new_n215), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n433), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n238), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n432), .B1(new_n309), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n443), .B1(new_n446), .B2(new_n441), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT30), .ZN(new_n449));
  XNOR2_X1  g248(.A(G8gat), .B(G36gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(G64gat), .B(G92gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n448), .A2(new_n449), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n446), .A2(new_n441), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n442), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n433), .A2(new_n441), .A3(new_n443), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n457), .A3(new_n453), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT30), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n453), .B1(new_n456), .B2(new_n457), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n454), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n431), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT35), .B1(new_n354), .B2(new_n462), .ZN(new_n463));
  AND4_X1   g262(.A1(new_n347), .A2(new_n353), .A3(new_n264), .A4(new_n263), .ZN(new_n464));
  XOR2_X1   g263(.A(KEYINPUT92), .B(KEYINPUT35), .Z(new_n465));
  NAND2_X1  g264(.A1(new_n431), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n461), .A2(KEYINPUT89), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n456), .A2(new_n457), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n452), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n470), .A2(new_n458), .A3(KEYINPUT30), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT89), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n471), .A2(new_n472), .A3(new_n454), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n464), .A2(new_n467), .A3(new_n475), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n463), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n414), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n416), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n390), .A2(new_n391), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n396), .B1(new_n480), .B2(new_n387), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n379), .A2(KEYINPUT83), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n482), .A2(KEYINPUT5), .A3(new_n385), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n412), .B(new_n407), .C1(new_n481), .C2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT85), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n397), .A2(new_n417), .A3(new_n412), .A4(new_n407), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT6), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n479), .B1(new_n487), .B2(new_n478), .ZN(new_n488));
  INV_X1    g287(.A(new_n458), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT37), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n453), .B1(new_n448), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT38), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n433), .A2(new_n441), .A3(new_n442), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT37), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n442), .B1(new_n446), .B2(new_n441), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n492), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n489), .B1(new_n491), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n488), .A2(new_n498), .A3(KEYINPUT90), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n452), .B1(new_n469), .B2(KEYINPUT37), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n448), .A2(new_n490), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT38), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT90), .B1(new_n488), .B2(new_n498), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OR2_X1    g304(.A1(new_n426), .A2(new_n356), .ZN(new_n506));
  OR2_X1    g305(.A1(new_n506), .A2(KEYINPUT39), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT39), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n366), .A2(new_n378), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n508), .B1(new_n509), .B2(new_n356), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n413), .B1(new_n506), .B2(new_n510), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n507), .A2(KEYINPUT40), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT40), .B1(new_n507), .B2(new_n511), .ZN(new_n513));
  NOR3_X1   g312(.A1(new_n512), .A2(new_n513), .A3(new_n478), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n461), .A2(KEYINPUT89), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n472), .B1(new_n471), .B2(new_n454), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n266), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT91), .B1(new_n505), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT90), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n458), .B1(new_n500), .B2(new_n496), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n520), .B1(new_n431), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n522), .A2(new_n499), .A3(new_n502), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n265), .B1(new_n474), .B2(new_n514), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT91), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n519), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n347), .A2(new_n353), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT36), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n529), .A2(KEYINPUT75), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(KEYINPUT75), .B(KEYINPUT36), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n347), .A2(new_n353), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n462), .A2(new_n265), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n477), .B1(new_n527), .B2(new_n536), .ZN(new_n537));
  XOR2_X1   g336(.A(G43gat), .B(G50gat), .Z(new_n538));
  INV_X1    g337(.A(KEYINPUT15), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(KEYINPUT95), .B(G36gat), .Z(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(G29gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n538), .A2(new_n539), .ZN(new_n543));
  OR3_X1    g342(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n544));
  OAI21_X1  g343(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AND4_X1   g345(.A1(new_n540), .A2(new_n542), .A3(new_n543), .A4(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n545), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT94), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n544), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n550), .B1(new_n549), .B2(new_n544), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n540), .B1(new_n551), .B2(new_n542), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n547), .B1(KEYINPUT96), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n553), .B1(KEYINPUT96), .B2(new_n552), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT17), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT16), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n556), .A2(G1gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(G15gat), .B(G22gat), .ZN(new_n558));
  MUX2_X1   g357(.A(G1gat), .B(new_n557), .S(new_n558), .Z(new_n559));
  INV_X1    g358(.A(G8gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n555), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n554), .A2(new_n561), .ZN(new_n564));
  NAND2_X1  g363(.A1(G229gat), .A2(G233gat), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT18), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G113gat), .B(G141gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT11), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G169gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT93), .B(G197gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT12), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n568), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n563), .A2(KEYINPUT18), .A3(new_n564), .A4(new_n565), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n565), .B(KEYINPUT13), .Z(new_n577));
  NOR2_X1   g376(.A1(new_n554), .A2(new_n561), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT98), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n578), .B1(new_n579), .B2(new_n564), .ZN(new_n580));
  NOR3_X1   g379(.A1(new_n554), .A2(KEYINPUT98), .A3(new_n561), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n577), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n576), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(KEYINPUT99), .B1(new_n575), .B2(new_n583), .ZN(new_n584));
  AND2_X1   g383(.A1(new_n576), .A2(new_n582), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT99), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n585), .A2(new_n586), .A3(new_n568), .A4(new_n574), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n574), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT97), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n568), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(new_n585), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n568), .A2(new_n590), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n589), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT100), .ZN(new_n595));
  AND3_X1   g394(.A1(new_n588), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n595), .B1(new_n588), .B2(new_n594), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n537), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G57gat), .B(G64gat), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n601));
  OR2_X1    g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(G71gat), .B(G78gat), .Z(new_n603));
  OR2_X1    g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n603), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT21), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G231gat), .A2(G233gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G127gat), .B(G155gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n562), .B1(new_n607), .B2(new_n606), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G183gat), .B(G211gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(G232gat), .A2(G233gat), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n620), .A2(KEYINPUT41), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT101), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(G85gat), .A2(G92gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT7), .ZN(new_n625));
  INV_X1    g424(.A(G99gat), .ZN(new_n626));
  INV_X1    g425(.A(G106gat), .ZN(new_n627));
  OAI21_X1  g426(.A(KEYINPUT8), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n625), .B(new_n628), .C1(G85gat), .C2(G92gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(G99gat), .B(G106gat), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n629), .B(new_n630), .Z(new_n631));
  NAND2_X1  g430(.A1(new_n555), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n629), .B(new_n630), .ZN(new_n633));
  AOI22_X1  g432(.A1(new_n554), .A2(new_n633), .B1(KEYINPUT41), .B2(new_n620), .ZN(new_n634));
  XNOR2_X1  g433(.A(G190gat), .B(G218gat), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n632), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n636), .B1(new_n632), .B2(new_n634), .ZN(new_n639));
  XNOR2_X1  g438(.A(G134gat), .B(G162gat), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NOR3_X1   g440(.A1(new_n638), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n632), .A2(new_n634), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n635), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n640), .B1(new_n644), .B2(new_n637), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n623), .B1(new_n642), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n641), .B1(new_n638), .B2(new_n639), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n644), .A2(new_n637), .A3(new_n640), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n647), .A2(new_n622), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n618), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n631), .A2(new_n606), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n633), .A2(new_n605), .A3(new_n604), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT10), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n654), .A2(KEYINPUT102), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n652), .A2(new_n653), .A3(new_n655), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT102), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n653), .A2(new_n655), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(G230gat), .A2(G233gat), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(G120gat), .B(G148gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(G176gat), .B(G204gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n665), .B(new_n669), .C1(new_n654), .C2(new_n664), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n654), .A2(new_n664), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT103), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n663), .A2(new_n672), .A3(new_n664), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n661), .B1(new_n656), .B2(new_n659), .ZN(new_n674));
  INV_X1    g473(.A(new_n664), .ZN(new_n675));
  OAI21_X1  g474(.A(KEYINPUT103), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n671), .B1(new_n673), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n670), .B1(new_n677), .B2(new_n669), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n651), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n599), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n682), .A2(new_n431), .ZN(new_n683));
  XOR2_X1   g482(.A(new_n683), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g483(.A1(new_n682), .A2(new_n475), .ZN(new_n685));
  OAI21_X1  g484(.A(KEYINPUT42), .B1(new_n685), .B2(new_n560), .ZN(new_n686));
  XOR2_X1   g485(.A(KEYINPUT16), .B(G8gat), .Z(new_n687));
  NAND2_X1  g486(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  MUX2_X1   g487(.A(KEYINPUT42), .B(new_n686), .S(new_n688), .Z(G1325gat));
  INV_X1    g488(.A(new_n534), .ZN(new_n690));
  OAI21_X1  g489(.A(G15gat), .B1(new_n682), .B2(new_n690), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n528), .A2(G15gat), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n691), .B1(new_n682), .B2(new_n692), .ZN(G1326gat));
  NOR2_X1   g492(.A1(new_n682), .A2(new_n266), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT43), .B(G22gat), .Z(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1327gat));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697));
  AND3_X1   g496(.A1(new_n523), .A2(new_n525), .A3(new_n524), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n525), .B1(new_n523), .B2(new_n524), .ZN(new_n699));
  OAI211_X1 g498(.A(new_n536), .B(KEYINPUT107), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n463), .A2(new_n476), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(KEYINPUT107), .B1(new_n527), .B2(new_n536), .ZN(new_n703));
  OAI211_X1 g502(.A(new_n697), .B(new_n650), .C1(new_n702), .C2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT108), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n650), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n536), .B1(new_n698), .B2(new_n699), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n707), .B1(new_n708), .B2(new_n701), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT106), .B1(new_n709), .B2(new_n697), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n711), .B(KEYINPUT44), .C1(new_n537), .C2(new_n707), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n708), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n715), .A2(new_n701), .A3(new_n700), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n716), .A2(KEYINPUT108), .A3(new_n697), .A4(new_n650), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n706), .A2(new_n713), .A3(new_n717), .ZN(new_n718));
  XOR2_X1   g517(.A(new_n678), .B(KEYINPUT105), .Z(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n588), .A2(new_n594), .ZN(new_n721));
  INV_X1    g520(.A(new_n618), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n718), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT109), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n718), .A2(KEYINPUT109), .A3(new_n723), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(G29gat), .B1(new_n728), .B2(new_n431), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n618), .A2(new_n650), .A3(new_n679), .ZN(new_n730));
  XOR2_X1   g529(.A(new_n730), .B(KEYINPUT104), .Z(new_n731));
  NAND2_X1  g530(.A1(new_n599), .A2(new_n731), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n732), .A2(G29gat), .A3(new_n431), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n733), .B(KEYINPUT45), .Z(new_n734));
  NAND2_X1  g533(.A1(new_n729), .A2(new_n734), .ZN(G1328gat));
  OAI21_X1  g534(.A(new_n541), .B1(new_n728), .B2(new_n475), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n732), .A2(new_n475), .A3(new_n541), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT46), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(G1329gat));
  OR3_X1    g538(.A1(new_n732), .A2(G43gat), .A3(new_n528), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT47), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n718), .A2(KEYINPUT109), .A3(new_n723), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT109), .B1(new_n718), .B2(new_n723), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n744), .A2(new_n745), .A3(new_n690), .ZN(new_n746));
  INV_X1    g545(.A(G43gat), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n743), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT110), .ZN(new_n749));
  OAI21_X1  g548(.A(G43gat), .B1(new_n724), .B2(new_n690), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n741), .B1(new_n750), .B2(new_n740), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n748), .A2(new_n749), .A3(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n726), .A2(new_n534), .A3(new_n727), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n742), .B1(new_n754), .B2(G43gat), .ZN(new_n755));
  OAI21_X1  g554(.A(KEYINPUT110), .B1(new_n755), .B2(new_n751), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n753), .A2(new_n756), .ZN(G1330gat));
  INV_X1    g556(.A(KEYINPUT48), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n732), .A2(G50gat), .A3(new_n266), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n718), .A2(new_n265), .A3(new_n723), .ZN(new_n760));
  AOI211_X1 g559(.A(new_n758), .B(new_n759), .C1(new_n760), .C2(G50gat), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n761), .A2(KEYINPUT111), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n761), .A2(KEYINPUT111), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n726), .A2(new_n265), .A3(new_n727), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n759), .B1(new_n764), .B2(G50gat), .ZN(new_n765));
  OAI22_X1  g564(.A1(new_n762), .A2(new_n763), .B1(new_n765), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g565(.A1(new_n716), .A2(new_n721), .A3(new_n651), .A4(new_n720), .ZN(new_n767));
  OR2_X1    g566(.A1(new_n767), .A2(new_n431), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G57gat), .ZN(G1332gat));
  OR2_X1    g568(.A1(new_n767), .A2(KEYINPUT112), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n767), .A2(KEYINPUT112), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n770), .A2(new_n474), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n773));
  AND2_X1   g572(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n775), .B1(new_n773), .B2(new_n772), .ZN(G1333gat));
  NAND4_X1  g575(.A1(new_n770), .A2(G71gat), .A3(new_n534), .A4(new_n771), .ZN(new_n777));
  INV_X1    g576(.A(G71gat), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n778), .B1(new_n767), .B2(new_n528), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT50), .ZN(G1334gat));
  NAND3_X1  g580(.A1(new_n770), .A2(new_n265), .A3(new_n771), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(G78gat), .ZN(G1335gat));
  INV_X1    g582(.A(new_n721), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n784), .A2(new_n722), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n718), .A2(new_n678), .A3(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n787));
  OR2_X1    g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(G85gat), .B1(new_n790), .B2(new_n431), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n716), .A2(new_n650), .A3(new_n785), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT51), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n679), .A2(G85gat), .A3(new_n431), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n791), .A2(new_n796), .ZN(G1336gat));
  OAI21_X1  g596(.A(G92gat), .B1(new_n786), .B2(new_n475), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n719), .A2(G92gat), .A3(new_n475), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n794), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(KEYINPUT115), .A2(KEYINPUT52), .ZN(new_n801));
  AND2_X1   g600(.A1(KEYINPUT115), .A2(KEYINPUT52), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n798), .B(new_n800), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT114), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n800), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n794), .A2(KEYINPUT114), .A3(new_n799), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n788), .A2(new_n474), .A3(new_n789), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n807), .B1(new_n808), .B2(G92gat), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n803), .B1(new_n809), .B2(new_n810), .ZN(G1337gat));
  OAI21_X1  g610(.A(G99gat), .B1(new_n790), .B2(new_n690), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n679), .A2(new_n528), .A3(G99gat), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n794), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(G1338gat));
  AND4_X1   g614(.A1(new_n627), .A2(new_n794), .A3(new_n265), .A4(new_n720), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n816), .A2(KEYINPUT53), .ZN(new_n817));
  OAI21_X1  g616(.A(G106gat), .B1(new_n786), .B2(new_n266), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n788), .A2(new_n265), .A3(new_n789), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n816), .B1(new_n820), .B2(G106gat), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n819), .B1(new_n821), .B2(new_n822), .ZN(G1339gat));
  NAND3_X1  g622(.A1(new_n651), .A2(new_n721), .A3(new_n679), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825));
  XOR2_X1   g624(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n826));
  AND3_X1   g625(.A1(new_n673), .A2(new_n676), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n674), .A2(new_n675), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(KEYINPUT54), .B1(new_n674), .B2(new_n675), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n668), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n825), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(KEYINPUT117), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n673), .A2(new_n676), .A3(new_n826), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n665), .A2(KEYINPUT54), .A3(new_n828), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n834), .A2(new_n835), .A3(KEYINPUT55), .A4(new_n668), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n834), .A2(new_n668), .A3(new_n835), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT117), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n837), .A2(new_n838), .A3(new_n825), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n833), .A2(new_n670), .A3(new_n836), .A4(new_n839), .ZN(new_n840));
  OR3_X1    g639(.A1(new_n580), .A2(new_n581), .A3(new_n577), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n565), .B1(new_n563), .B2(new_n564), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n573), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n650), .A2(new_n588), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n588), .A2(new_n678), .A3(new_n844), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n847), .B1(new_n840), .B2(new_n721), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n846), .B1(new_n848), .B2(new_n707), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n824), .B1(new_n849), .B2(new_n722), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n474), .A2(new_n431), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n852), .A2(new_n464), .ZN(new_n853));
  AOI21_X1  g652(.A(G113gat), .B1(new_n853), .B2(new_n784), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n598), .A2(new_n310), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n854), .B1(new_n853), .B2(new_n855), .ZN(G1340gat));
  AOI21_X1  g655(.A(G120gat), .B1(new_n853), .B2(new_n678), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n719), .A2(new_n313), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n857), .B1(new_n853), .B2(new_n858), .ZN(G1341gat));
  NAND2_X1  g658(.A1(new_n853), .A2(new_n722), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(G127gat), .ZN(G1342gat));
  AND3_X1   g660(.A1(new_n852), .A2(new_n464), .A3(new_n650), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n317), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(KEYINPUT56), .ZN(new_n864));
  XOR2_X1   g663(.A(new_n864), .B(KEYINPUT118), .Z(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(KEYINPUT56), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n865), .B(new_n866), .C1(new_n317), .C2(new_n862), .ZN(G1343gat));
  INV_X1    g666(.A(KEYINPUT58), .ZN(new_n868));
  INV_X1    g667(.A(new_n824), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n848), .A2(new_n707), .ZN(new_n870));
  INV_X1    g669(.A(new_n846), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n869), .B1(new_n872), .B2(new_n618), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n690), .A2(new_n851), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n873), .A2(new_n266), .A3(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n598), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n875), .A2(new_n224), .A3(new_n876), .ZN(new_n877));
  XOR2_X1   g676(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n837), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(new_n670), .A3(new_n836), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(KEYINPUT120), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT120), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n880), .A2(new_n883), .A3(new_n670), .A4(new_n836), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n882), .B(new_n884), .C1(new_n596), .C2(new_n597), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n650), .B1(new_n885), .B2(new_n847), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n618), .B1(new_n886), .B2(new_n846), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n887), .A2(new_n824), .ZN(new_n888));
  OAI21_X1  g687(.A(KEYINPUT57), .B1(new_n888), .B2(new_n266), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n873), .A2(new_n266), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT57), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n874), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(KEYINPUT121), .A3(new_n876), .ZN(new_n895));
  INV_X1    g694(.A(new_n372), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(KEYINPUT121), .B1(new_n894), .B2(new_n876), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n868), .B(new_n877), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n896), .B1(new_n893), .B2(new_n721), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n900), .A2(new_n877), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n899), .B1(new_n868), .B2(new_n901), .ZN(G1344gat));
  NAND3_X1  g701(.A1(new_n875), .A2(new_n368), .A3(new_n678), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT59), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n266), .A2(KEYINPUT57), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n681), .A2(new_n598), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n906), .B1(new_n887), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n891), .B1(new_n850), .B2(new_n265), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n911), .A2(new_n679), .A3(new_n874), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n912), .A2(KEYINPUT122), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n368), .B1(new_n912), .B2(KEYINPUT122), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n904), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AOI211_X1 g714(.A(KEYINPUT59), .B(new_n368), .C1(new_n894), .C2(new_n678), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n903), .B1(new_n915), .B2(new_n916), .ZN(G1345gat));
  OAI21_X1  g716(.A(G155gat), .B1(new_n893), .B2(new_n618), .ZN(new_n918));
  INV_X1    g717(.A(new_n875), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n618), .A2(G155gat), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  XOR2_X1   g720(.A(new_n921), .B(KEYINPUT123), .Z(G1346gat));
  OAI21_X1  g721(.A(G162gat), .B1(new_n893), .B2(new_n707), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n707), .A2(G162gat), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n923), .B1(new_n919), .B2(new_n924), .ZN(G1347gat));
  NOR3_X1   g724(.A1(new_n354), .A2(new_n475), .A3(new_n488), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n850), .A2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(G169gat), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n927), .A2(new_n928), .A3(new_n598), .ZN(new_n929));
  INV_X1    g728(.A(new_n927), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n784), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n929), .B1(new_n928), .B2(new_n931), .ZN(G1348gat));
  OAI21_X1  g731(.A(G176gat), .B1(new_n927), .B2(new_n719), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n679), .A2(G176gat), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n933), .B1(new_n927), .B2(new_n934), .ZN(G1349gat));
  NOR2_X1   g734(.A1(new_n927), .A2(new_n618), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(new_n283), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n937), .B1(new_n292), .B2(new_n936), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT60), .ZN(G1350gat));
  NAND2_X1  g738(.A1(new_n930), .A2(new_n650), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(G190gat), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT61), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n942), .B1(G190gat), .B2(new_n940), .ZN(G1351gat));
  NOR2_X1   g742(.A1(new_n475), .A2(new_n488), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n690), .A2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n890), .A2(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(G197gat), .B1(new_n948), .B2(new_n784), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n911), .A2(new_n945), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n876), .A2(G197gat), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(G1352gat));
  NOR2_X1   g751(.A1(new_n679), .A2(G204gat), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n948), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(KEYINPUT124), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT62), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT124), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n948), .A2(new_n957), .A3(new_n953), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n955), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT125), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n959), .B(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n956), .B1(new_n955), .B2(new_n958), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n950), .A2(new_n720), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n962), .B1(G204gat), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n961), .A2(new_n964), .ZN(G1353gat));
  OR3_X1    g764(.A1(new_n947), .A2(new_n202), .A3(new_n618), .ZN(new_n966));
  INV_X1    g765(.A(G211gat), .ZN(new_n967));
  NOR4_X1   g766(.A1(new_n908), .A2(new_n909), .A3(new_n618), .A4(new_n945), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT126), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n887), .A2(new_n907), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(new_n905), .ZN(new_n972));
  OAI21_X1  g771(.A(KEYINPUT57), .B1(new_n873), .B2(new_n266), .ZN(new_n973));
  NAND4_X1  g772(.A1(new_n972), .A2(new_n722), .A3(new_n973), .A4(new_n946), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(KEYINPUT126), .ZN(new_n975));
  AOI21_X1  g774(.A(KEYINPUT63), .B1(new_n970), .B2(new_n975), .ZN(new_n976));
  NAND4_X1  g775(.A1(new_n910), .A2(new_n969), .A3(new_n722), .A4(new_n946), .ZN(new_n977));
  AND4_X1   g776(.A1(KEYINPUT63), .A2(new_n975), .A3(G211gat), .A4(new_n977), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n966), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(KEYINPUT127), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT127), .ZN(new_n981));
  OAI211_X1 g780(.A(new_n981), .B(new_n966), .C1(new_n976), .C2(new_n978), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n980), .A2(new_n982), .ZN(G1354gat));
  INV_X1    g782(.A(G218gat), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n948), .A2(new_n984), .A3(new_n650), .ZN(new_n985));
  NOR3_X1   g784(.A1(new_n911), .A2(new_n707), .A3(new_n945), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n985), .B1(new_n986), .B2(new_n984), .ZN(G1355gat));
endmodule


