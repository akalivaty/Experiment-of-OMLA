//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 0 1 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 0 0 1 1 1 0 0 0 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n551,
    new_n553, new_n554, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n563, new_n564, new_n565, new_n566, new_n568, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n607, new_n610, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1162, new_n1163, new_n1164, new_n1165;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  XNOR2_X1  g033(.A(KEYINPUT3), .B(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G125), .ZN(new_n460));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  AOI22_X1  g039(.A1(new_n462), .A2(G2105), .B1(G101), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  AND3_X1   g041(.A1(KEYINPUT64), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(KEYINPUT3), .B1(KEYINPUT64), .B2(G2104), .ZN(new_n468));
  OAI211_X1 g043(.A(G137), .B(new_n466), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT65), .ZN(new_n470));
  XNOR2_X1  g045(.A(new_n469), .B(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  NOR2_X1   g048(.A1(new_n467), .A2(new_n468), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(new_n466), .ZN(new_n476));
  INV_X1    g051(.A(G136), .ZN(new_n477));
  NOR2_X1   g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(new_n466), .B2(G112), .ZN(new_n479));
  OAI22_X1  g054(.A1(new_n476), .A2(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n475), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n480), .B1(G124), .B2(new_n482), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT66), .ZN(G162));
  INV_X1    g059(.A(KEYINPUT67), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(KEYINPUT4), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(KEYINPUT67), .ZN(new_n488));
  OAI21_X1  g063(.A(G138), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  AND2_X1   g064(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n490));
  NOR2_X1   g065(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n466), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(KEYINPUT68), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  OAI211_X1 g068(.A(G138), .B(new_n466), .C1(new_n467), .C2(new_n468), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n487), .A2(KEYINPUT67), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n485), .A2(KEYINPUT4), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT68), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n499), .A2(new_n500), .A3(new_n466), .A4(new_n459), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n493), .A2(new_n495), .A3(new_n501), .ZN(new_n502));
  AND2_X1   g077(.A1(new_n464), .A2(G102), .ZN(new_n503));
  NAND2_X1  g078(.A1(G114), .A2(G2104), .ZN(new_n504));
  INV_X1    g079(.A(G126), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n504), .B1(new_n474), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n503), .B1(new_n506), .B2(G2105), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(KEYINPUT69), .ZN(new_n510));
  AND3_X1   g085(.A1(new_n510), .A2(KEYINPUT6), .A3(G651), .ZN(new_n511));
  AOI21_X1  g086(.A(KEYINPUT6), .B1(new_n510), .B2(G651), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G50), .B1(G75), .B2(G651), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  OR2_X1    g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n511), .A2(new_n512), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n522), .A2(G88), .B1(G62), .B2(new_n524), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n516), .A2(new_n525), .ZN(G166));
  NOR2_X1   g101(.A1(new_n517), .A2(new_n515), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G51), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n522), .A2(G89), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n524), .A2(G63), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n528), .A2(new_n529), .A3(new_n530), .A4(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  AND2_X1   g109(.A1(new_n518), .A2(new_n520), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n535), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n523), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n537), .B1(G52), .B2(new_n527), .ZN(new_n538));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  INV_X1    g114(.A(new_n522), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  AOI22_X1  g117(.A1(G43), .A2(new_n527), .B1(new_n522), .B2(G81), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT70), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n535), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n523), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT71), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(G188));
  NAND2_X1  g130(.A1(new_n527), .A2(G53), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT9), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n521), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n522), .A2(G91), .B1(G651), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n557), .A2(new_n561), .ZN(G299));
  NAND2_X1  g137(.A1(G166), .A2(KEYINPUT72), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n516), .A2(new_n525), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT72), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n563), .A2(new_n566), .ZN(G303));
  NAND2_X1  g142(.A1(new_n527), .A2(G49), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n522), .A2(G87), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n535), .B2(G74), .ZN(new_n570));
  AND3_X1   g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(G288));
  NAND2_X1  g147(.A1(new_n522), .A2(G86), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT73), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n522), .A2(KEYINPUT73), .A3(G86), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n521), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G651), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n513), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G48), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n577), .A2(new_n585), .ZN(G305));
  AOI22_X1  g161(.A1(new_n535), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n587), .A2(new_n523), .ZN(new_n588));
  XOR2_X1   g163(.A(new_n588), .B(KEYINPUT74), .Z(new_n589));
  AOI22_X1  g164(.A1(G47), .A2(new_n527), .B1(new_n522), .B2(G85), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  XOR2_X1   g167(.A(new_n592), .B(KEYINPUT75), .Z(new_n593));
  INV_X1    g168(.A(G92), .ZN(new_n594));
  OR3_X1    g169(.A1(new_n540), .A2(KEYINPUT10), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G66), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n521), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n527), .A2(G54), .B1(G651), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(KEYINPUT10), .B1(new_n540), .B2(new_n594), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n595), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n593), .B1(G868), .B2(new_n602), .ZN(G284));
  OAI21_X1  g178(.A(new_n593), .B1(G868), .B2(new_n602), .ZN(G321));
  NAND2_X1  g179(.A1(G286), .A2(G868), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT76), .Z(new_n606));
  INV_X1    g181(.A(G299), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(G868), .B2(new_n607), .ZN(G297));
  OAI21_X1  g183(.A(new_n606), .B1(G868), .B2(new_n607), .ZN(G280));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n602), .B1(new_n610), .B2(G860), .ZN(G148));
  NAND2_X1  g186(.A1(new_n602), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(new_n548), .B2(G868), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n482), .A2(G123), .ZN(new_n616));
  INV_X1    g191(.A(new_n476), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G135), .ZN(new_n618));
  NOR2_X1   g193(.A1(G99), .A2(G2105), .ZN(new_n619));
  OAI21_X1  g194(.A(G2104), .B1(new_n466), .B2(G111), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n616), .B(new_n618), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(G2096), .Z(new_n622));
  NOR2_X1   g197(.A1(new_n492), .A2(new_n463), .ZN(new_n623));
  XOR2_X1   g198(.A(KEYINPUT77), .B(KEYINPUT12), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT13), .B(G2100), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n622), .A2(new_n627), .ZN(G156));
  XNOR2_X1  g203(.A(KEYINPUT15), .B(G2430), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2435), .ZN(new_n630));
  XOR2_X1   g205(.A(G2427), .B(G2438), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(KEYINPUT14), .ZN(new_n633));
  XOR2_X1   g208(.A(G2451), .B(G2454), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n633), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G1341), .B(G1348), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n638), .B(new_n639), .Z(new_n640));
  AND2_X1   g215(.A1(new_n640), .A2(G14), .ZN(G401));
  XNOR2_X1  g216(.A(G2072), .B(G2078), .ZN(new_n642));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT78), .ZN(new_n644));
  XOR2_X1   g219(.A(G2067), .B(G2678), .Z(new_n645));
  NOR2_X1   g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT79), .B(KEYINPUT18), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n642), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT80), .Z(new_n649));
  XNOR2_X1  g224(.A(G2096), .B(G2100), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n644), .A2(new_n645), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(KEYINPUT17), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n647), .B1(new_n653), .B2(new_n646), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n651), .B(new_n654), .ZN(G227));
  XOR2_X1   g230(.A(G1956), .B(G2474), .Z(new_n656));
  XOR2_X1   g231(.A(G1961), .B(G1966), .Z(new_n657));
  NOR2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1971), .B(G1976), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT19), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n656), .A2(new_n657), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT20), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n659), .A2(new_n661), .A3(new_n663), .ZN(new_n667));
  OAI211_X1 g242(.A(new_n666), .B(new_n667), .C1(new_n665), .C2(new_n664), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT21), .B(G1986), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G1991), .B(G1996), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT81), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n670), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT22), .B(G1981), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(G229));
  INV_X1    g250(.A(KEYINPUT94), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n676), .B1(G5), .B2(G16), .ZN(new_n677));
  OR3_X1    g252(.A1(new_n676), .A2(G5), .A3(G16), .ZN(new_n678));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  OAI211_X1 g254(.A(new_n677), .B(new_n678), .C1(G301), .C2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G1961), .ZN(new_n681));
  INV_X1    g256(.A(G29), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT24), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n682), .B1(new_n683), .B2(G34), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n684), .A2(KEYINPUT89), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(G34), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n684), .A2(KEYINPUT89), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(new_n472), .B2(new_n682), .ZN(new_n689));
  INV_X1    g264(.A(G2084), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(G164), .A2(G29), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(G27), .B2(G29), .ZN(new_n693));
  INV_X1    g268(.A(G2078), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n681), .A2(new_n691), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n679), .A2(G22), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G166), .B2(new_n679), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n698), .A2(G1971), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(G1971), .ZN(new_n700));
  NOR2_X1   g275(.A1(G16), .A2(G23), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(new_n571), .B2(G16), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT33), .B(G1976), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n699), .A2(new_n700), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n679), .A2(G6), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n584), .B1(new_n575), .B2(new_n576), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(new_n707), .B2(new_n679), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT32), .B(G1981), .Z(new_n709));
  XOR2_X1   g284(.A(new_n708), .B(new_n709), .Z(new_n710));
  INV_X1    g285(.A(KEYINPUT86), .ZN(new_n711));
  OAI22_X1  g286(.A1(new_n705), .A2(new_n710), .B1(new_n711), .B2(KEYINPUT34), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(KEYINPUT34), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  MUX2_X1   g290(.A(G24), .B(G290), .S(G16), .Z(new_n716));
  XOR2_X1   g291(.A(KEYINPUT84), .B(G1986), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT85), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n716), .B(new_n718), .Z(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n682), .A2(G25), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n482), .A2(G119), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n617), .A2(G131), .ZN(new_n723));
  NOR2_X1   g298(.A1(G95), .A2(G2105), .ZN(new_n724));
  OAI21_X1  g299(.A(G2104), .B1(new_n466), .B2(G107), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n722), .B(new_n723), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n726), .A2(KEYINPUT82), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(KEYINPUT82), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n721), .B1(new_n730), .B2(new_n682), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT35), .B(G1991), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT83), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n731), .B(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n720), .A2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT36), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n715), .B(new_n735), .C1(KEYINPUT87), .C2(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n736), .A2(KEYINPUT87), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n720), .A2(new_n734), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n738), .B1(new_n739), .B2(new_n714), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n696), .B1(new_n737), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n464), .A2(G103), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT25), .Z(new_n743));
  AOI22_X1  g318(.A1(new_n459), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n744));
  INV_X1    g319(.A(G139), .ZN(new_n745));
  OAI221_X1 g320(.A(new_n743), .B1(new_n744), .B2(new_n466), .C1(new_n476), .C2(new_n745), .ZN(new_n746));
  MUX2_X1   g321(.A(G33), .B(new_n746), .S(G29), .Z(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(G2072), .Z(new_n748));
  NAND2_X1  g323(.A1(new_n679), .A2(G4), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n602), .B2(new_n679), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G1348), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n750), .A2(G1348), .ZN(new_n752));
  NAND2_X1  g327(.A1(G168), .A2(G16), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G16), .B2(G21), .ZN(new_n754));
  INV_X1    g329(.A(G1966), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g331(.A1(new_n748), .A2(new_n751), .A3(new_n752), .A4(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n679), .A2(G20), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT95), .Z(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT23), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G299), .B2(G16), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT96), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(G1956), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n764), .A2(new_n765), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n741), .A2(new_n758), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n682), .A2(G26), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n482), .A2(G128), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n617), .A2(G140), .ZN(new_n772));
  OR2_X1    g347(.A1(G104), .A2(G2105), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n773), .B(G2104), .C1(G116), .C2(new_n466), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n771), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n770), .B1(new_n776), .B2(new_n682), .ZN(new_n777));
  MUX2_X1   g352(.A(new_n770), .B(new_n777), .S(KEYINPUT28), .Z(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT88), .B(G2067), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n694), .B2(new_n693), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n769), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(G29), .A2(G35), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G162), .B2(G29), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT29), .B(G2090), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n679), .A2(G19), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n548), .B2(new_n679), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(G1341), .Z(new_n789));
  OR2_X1    g364(.A1(new_n754), .A2(new_n755), .ZN(new_n790));
  OAI221_X1 g365(.A(new_n790), .B1(new_n690), .B2(new_n689), .C1(new_n778), .C2(new_n779), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n782), .A2(new_n786), .A3(new_n789), .A4(new_n792), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT30), .B(G28), .ZN(new_n794));
  OR2_X1    g369(.A1(KEYINPUT31), .A2(G11), .ZN(new_n795));
  NAND2_X1  g370(.A1(KEYINPUT31), .A2(G11), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n794), .A2(new_n682), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n621), .B2(new_n682), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT93), .Z(new_n799));
  NAND2_X1  g374(.A1(new_n682), .A2(G32), .ZN(new_n800));
  AOI22_X1  g375(.A1(G129), .A2(new_n482), .B1(new_n617), .B2(G141), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n464), .A2(G105), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT90), .B(KEYINPUT26), .ZN(new_n804));
  NAND3_X1  g379(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT91), .Z(new_n808));
  OAI21_X1  g383(.A(new_n800), .B1(new_n808), .B2(new_n682), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT27), .B(G1996), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT92), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n809), .B(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  NOR3_X1   g388(.A1(new_n793), .A2(new_n799), .A3(new_n813), .ZN(G311));
  AND3_X1   g389(.A1(new_n782), .A2(new_n789), .A3(new_n792), .ZN(new_n815));
  INV_X1    g390(.A(new_n799), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n815), .A2(new_n816), .A3(new_n812), .A4(new_n786), .ZN(G150));
  AOI22_X1  g392(.A1(G55), .A2(new_n527), .B1(new_n522), .B2(G93), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT97), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n535), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n523), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G860), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT98), .B(KEYINPUT37), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n548), .A2(new_n821), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n548), .A2(new_n821), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n601), .A2(new_n610), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n824), .B1(new_n831), .B2(G860), .ZN(G145));
  NAND2_X1  g407(.A1(new_n508), .A2(KEYINPUT99), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT99), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n502), .A2(new_n834), .A3(new_n507), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(new_n776), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT100), .ZN(new_n838));
  INV_X1    g413(.A(new_n807), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(new_n746), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n808), .B(new_n837), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n842), .A2(new_n746), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n482), .A2(KEYINPUT101), .A3(G130), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n617), .A2(G142), .ZN(new_n846));
  OR2_X1    g421(.A1(G106), .A2(G2105), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n847), .B(G2104), .C1(G118), .C2(new_n466), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT101), .ZN(new_n849));
  INV_X1    g424(.A(G130), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n849), .B1(new_n481), .B2(new_n850), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n845), .A2(new_n846), .A3(new_n848), .A4(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n729), .B(new_n852), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(new_n625), .Z(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n844), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT102), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n841), .A2(new_n843), .A3(new_n854), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n858), .A2(new_n857), .ZN(new_n860));
  XNOR2_X1  g435(.A(G162), .B(new_n472), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n621), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n859), .A2(new_n860), .A3(new_n863), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n864), .A2(KEYINPUT103), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n856), .A2(new_n858), .ZN(new_n866));
  AOI21_X1  g441(.A(G37), .B1(new_n866), .B2(new_n862), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n864), .A2(KEYINPUT103), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n865), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(KEYINPUT40), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT40), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n865), .A2(new_n871), .A3(new_n867), .A4(new_n868), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(G395));
  INV_X1    g448(.A(KEYINPUT104), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n827), .B(new_n612), .Z(new_n875));
  XNOR2_X1  g450(.A(new_n602), .B(G299), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT41), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n875), .A2(new_n876), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n874), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(KEYINPUT104), .B1(new_n875), .B2(new_n876), .ZN(new_n881));
  OR3_X1    g456(.A1(new_n880), .A2(new_n881), .A3(KEYINPUT42), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n564), .B(new_n707), .ZN(new_n883));
  XNOR2_X1  g458(.A(G290), .B(new_n571), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT105), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n885), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n886), .B(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(KEYINPUT42), .B1(new_n880), .B2(new_n881), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n882), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n888), .B1(new_n882), .B2(new_n889), .ZN(new_n891));
  OAI21_X1  g466(.A(G868), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(G868), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n821), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n894), .ZN(G295));
  NAND2_X1  g470(.A1(new_n892), .A2(new_n894), .ZN(G331));
  INV_X1    g471(.A(KEYINPUT108), .ZN(new_n897));
  INV_X1    g472(.A(new_n876), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT106), .ZN(new_n899));
  OAI21_X1  g474(.A(G301), .B1(new_n899), .B2(G168), .ZN(new_n900));
  NOR2_X1   g475(.A1(G286), .A2(KEYINPUT106), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n900), .B(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n902), .A2(new_n825), .A3(new_n826), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT107), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n902), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n827), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(new_n903), .ZN(new_n909));
  AOI211_X1 g484(.A(new_n898), .B(new_n906), .C1(new_n909), .C2(KEYINPUT107), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n877), .B1(new_n903), .B2(new_n908), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n897), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n906), .B1(new_n909), .B2(KEYINPUT107), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n911), .B1(new_n913), .B2(new_n876), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT108), .ZN(new_n915));
  INV_X1    g490(.A(new_n888), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n912), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(G37), .B1(new_n914), .B2(new_n888), .ZN(new_n918));
  AOI21_X1  g493(.A(KEYINPUT43), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n909), .A2(new_n898), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(KEYINPUT109), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n913), .A2(new_n877), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n916), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n918), .A2(new_n923), .A3(KEYINPUT43), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT44), .B1(new_n919), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT43), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n926), .B1(new_n917), .B2(new_n918), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n923), .A2(new_n926), .A3(new_n918), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n925), .B1(KEYINPUT44), .B2(new_n929), .ZN(G397));
  AND3_X1   g505(.A1(new_n465), .A2(new_n471), .A3(G40), .ZN(new_n931));
  AOI21_X1  g506(.A(G1384), .B1(new_n502), .B2(new_n507), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n931), .B1(new_n932), .B2(KEYINPUT45), .ZN(new_n933));
  INV_X1    g508(.A(G1384), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n502), .A2(new_n834), .A3(new_n507), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n834), .B1(new_n502), .B2(new_n507), .ZN(new_n936));
  OAI211_X1 g511(.A(KEYINPUT45), .B(new_n934), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT110), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT110), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n836), .A2(new_n939), .A3(KEYINPUT45), .A4(new_n934), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n933), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n932), .A2(KEYINPUT50), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n932), .A2(KEYINPUT50), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n931), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OAI22_X1  g520(.A1(new_n941), .A2(G1971), .B1(G2090), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT55), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n947), .B1(G303), .B2(G8), .ZN(new_n948));
  INV_X1    g523(.A(G8), .ZN(new_n949));
  AOI211_X1 g524(.A(KEYINPUT55), .B(new_n949), .C1(new_n563), .C2(new_n566), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n946), .A2(G8), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n951), .B1(new_n946), .B2(G8), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n931), .A2(new_n932), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(G8), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n955), .B(KEYINPUT111), .ZN(new_n956));
  INV_X1    g531(.A(G1976), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT52), .B1(G288), .B2(new_n957), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n956), .B(new_n958), .C1(new_n957), .C2(G288), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT111), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n955), .B(new_n960), .ZN(new_n961));
  NOR2_X1   g536(.A1(G288), .A2(new_n957), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT52), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n585), .A2(new_n573), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(G1981), .ZN(new_n965));
  INV_X1    g540(.A(G1981), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n707), .A2(KEYINPUT112), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT112), .B1(new_n707), .B2(new_n966), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n965), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g544(.A1(KEYINPUT113), .A2(KEYINPUT49), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI221_X1 g546(.A(new_n965), .B1(KEYINPUT113), .B2(KEYINPUT49), .C1(new_n967), .C2(new_n968), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(new_n956), .A3(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n959), .A2(new_n963), .A3(new_n973), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n952), .A2(new_n953), .A3(new_n974), .ZN(new_n975));
  XOR2_X1   g550(.A(KEYINPUT115), .B(G2084), .Z(new_n976));
  OAI211_X1 g551(.A(new_n931), .B(new_n976), .C1(new_n943), .C2(new_n944), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT114), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n508), .A2(new_n934), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n978), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n932), .A2(KEYINPUT114), .A3(KEYINPUT45), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n933), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n977), .B1(new_n983), .B2(G1966), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n984), .A2(G8), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n975), .A2(G168), .A3(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT63), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n975), .A2(KEYINPUT63), .A3(G168), .A4(new_n985), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n952), .A2(new_n963), .A3(new_n973), .A4(new_n959), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n973), .A2(new_n957), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n571), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n993), .B1(new_n968), .B2(new_n967), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n956), .ZN(new_n995));
  AND3_X1   g570(.A1(new_n990), .A2(new_n991), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT126), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT57), .ZN(new_n998));
  NAND2_X1  g573(.A1(G299), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n557), .A2(KEYINPUT57), .A3(new_n561), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(KEYINPUT56), .B(G2072), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n941), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n931), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n979), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1005), .B1(new_n1007), .B2(new_n942), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1008), .A2(G1956), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1002), .B1(new_n1004), .B2(new_n1010), .ZN(new_n1011));
  AOI211_X1 g586(.A(new_n1001), .B(new_n1009), .C1(new_n941), .C2(new_n1003), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1012), .A2(new_n601), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n954), .A2(KEYINPUT116), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT116), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n931), .A2(new_n1015), .A3(new_n932), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1017), .A2(G2067), .ZN(new_n1018));
  INV_X1    g593(.A(G1348), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1018), .B1(new_n1019), .B2(new_n945), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1011), .B1(new_n1013), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT119), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT61), .B1(new_n1012), .B2(new_n1011), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n938), .A2(new_n940), .ZN(new_n1026));
  INV_X1    g601(.A(new_n933), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n1026), .A2(new_n1027), .A3(new_n1003), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1001), .B1(new_n1028), .B2(new_n1009), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT61), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1004), .A2(new_n1002), .A3(new_n1010), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n1033));
  INV_X1    g608(.A(G1996), .ZN(new_n1034));
  AOI21_X1  g609(.A(G1384), .B1(new_n833), .B2(new_n835), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n939), .B1(new_n1035), .B2(KEYINPUT45), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n937), .A2(KEYINPUT110), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1034), .B(new_n1027), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  XOR2_X1   g613(.A(KEYINPUT58), .B(G1341), .Z(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1040), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n547), .B1(new_n1038), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT59), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1033), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1041), .B1(new_n941), .B2(new_n1034), .ZN(new_n1046));
  NOR4_X1   g621(.A1(new_n1046), .A2(KEYINPUT118), .A3(KEYINPUT59), .A4(new_n547), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT117), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT117), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1050), .B(KEYINPUT59), .C1(new_n1046), .C2(new_n547), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  AOI221_X4 g627(.A(new_n1024), .B1(new_n1025), .B2(new_n1032), .C1(new_n1048), .C2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1038), .A2(new_n1042), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1054), .A2(new_n1044), .A3(new_n548), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT118), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1043), .A2(new_n1033), .A3(new_n1044), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1052), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1025), .A2(new_n1032), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT119), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1053), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1020), .A2(KEYINPUT60), .ZN(new_n1062));
  XNOR2_X1  g637(.A(new_n1062), .B(new_n602), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1063), .B1(KEYINPUT60), .B2(new_n1020), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1023), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n1066));
  INV_X1    g641(.A(G1961), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n945), .A2(KEYINPUT122), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT122), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1069), .B1(new_n1008), .B2(G1961), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  OR2_X1    g646(.A1(new_n1035), .A2(KEYINPUT45), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1073), .A2(G2078), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1026), .A2(new_n1072), .A3(new_n931), .A4(new_n1074), .ZN(new_n1075));
  AOI211_X1 g650(.A(G2078), .B(new_n933), .C1(new_n938), .C2(new_n940), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1071), .B(new_n1075), .C1(new_n1076), .C2(KEYINPUT53), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1066), .B1(new_n1077), .B2(G171), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1026), .A2(new_n694), .A3(new_n1027), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n1073), .ZN(new_n1080));
  AOI22_X1  g655(.A1(new_n983), .A2(new_n1074), .B1(new_n945), .B2(new_n1067), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1080), .A2(G301), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT124), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT124), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1080), .A2(new_n1084), .A3(G301), .A4(new_n1081), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1078), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT125), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1078), .A2(new_n1083), .A3(KEYINPUT125), .A4(new_n1085), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1080), .A2(G301), .A3(new_n1075), .A4(new_n1071), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT53), .B1(new_n941), .B2(new_n694), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n983), .A2(new_n1074), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1093), .B1(G1961), .B2(new_n1008), .ZN(new_n1094));
  OAI21_X1  g669(.A(G171), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1091), .A2(KEYINPUT123), .A3(new_n1095), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1079), .A2(new_n1073), .B1(new_n1070), .B2(new_n1068), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT123), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1097), .A2(new_n1098), .A3(G301), .A4(new_n1075), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1096), .A2(new_n1066), .A3(new_n1099), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1100), .A2(new_n975), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT51), .B1(new_n985), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n1104));
  NOR2_X1   g679(.A1(G168), .A2(new_n949), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1102), .B1(new_n984), .B2(G8), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1103), .A2(new_n1104), .A3(new_n1106), .A4(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(KEYINPUT51), .B1(new_n985), .B2(new_n1105), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT51), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n984), .A2(G8), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1111), .B(new_n1106), .C1(new_n1112), .C2(KEYINPUT120), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT121), .B1(new_n1113), .B2(new_n1107), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1109), .A2(new_n1110), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n984), .A2(new_n1105), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1090), .A2(new_n1101), .A3(new_n1117), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n996), .B(new_n997), .C1(new_n1065), .C2(new_n1118), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1059), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(new_n1024), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1058), .A2(KEYINPUT119), .A3(new_n1059), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1123), .A2(new_n1124), .A3(new_n1064), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1118), .B1(new_n1125), .B2(new_n1022), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n990), .A2(new_n991), .A3(new_n995), .ZN(new_n1127));
  OAI21_X1  g702(.A(KEYINPUT126), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OR2_X1    g703(.A1(new_n1117), .A2(KEYINPUT62), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1117), .A2(KEYINPUT62), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1095), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1129), .A2(new_n1130), .A3(new_n975), .A4(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1119), .A2(new_n1128), .A3(new_n1132), .ZN(new_n1133));
  XOR2_X1   g708(.A(new_n775), .B(G2067), .Z(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1135), .B1(new_n808), .B2(new_n1034), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1136), .B1(new_n1034), .B2(new_n807), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n729), .B(new_n732), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  XOR2_X1   g714(.A(G290), .B(G1986), .Z(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1072), .A2(new_n1005), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1133), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT46), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1142), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1145), .B1(new_n1146), .B2(G1996), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1142), .B1(new_n839), .B2(new_n1135), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1142), .A2(KEYINPUT46), .A3(new_n1034), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  XOR2_X1   g725(.A(new_n1150), .B(KEYINPUT47), .Z(new_n1151));
  OR2_X1    g726(.A1(new_n729), .A2(new_n732), .ZN(new_n1152));
  OAI22_X1  g727(.A1(new_n1137), .A2(new_n1152), .B1(G2067), .B2(new_n775), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1153), .A2(new_n1142), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1139), .A2(new_n1146), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(KEYINPUT127), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n1146), .A2(G1986), .A3(G290), .ZN(new_n1157));
  XOR2_X1   g732(.A(new_n1157), .B(KEYINPUT48), .Z(new_n1158));
  AOI211_X1 g733(.A(new_n1151), .B(new_n1154), .C1(new_n1156), .C2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1144), .A2(new_n1159), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g735(.A(G227), .ZN(new_n1162));
  OAI211_X1 g736(.A(G319), .B(new_n1162), .C1(new_n927), .C2(new_n928), .ZN(new_n1163));
  INV_X1    g737(.A(new_n1163), .ZN(new_n1164));
  NOR2_X1   g738(.A1(G401), .A2(G229), .ZN(new_n1165));
  AND3_X1   g739(.A1(new_n1164), .A2(new_n869), .A3(new_n1165), .ZN(G308));
  NAND3_X1  g740(.A1(new_n1164), .A2(new_n869), .A3(new_n1165), .ZN(G225));
endmodule


