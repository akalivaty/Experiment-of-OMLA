//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 1 1 1 1 1 1 0 1 1 0 1 1 1 0 1 1 0 0 0 1 0 0 1 0 1 0 0 1 1 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n835,
    new_n836, new_n837, new_n838, new_n840, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959;
  INV_X1    g000(.A(KEYINPUT94), .ZN(new_n202));
  INV_X1    g001(.A(G43gat), .ZN(new_n203));
  OR2_X1    g002(.A1(new_n203), .A2(G50gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(G50gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n204), .A2(KEYINPUT15), .A3(new_n205), .ZN(new_n206));
  OR2_X1    g005(.A1(KEYINPUT90), .A2(G50gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(KEYINPUT90), .A2(G50gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n207), .A2(new_n203), .A3(new_n208), .ZN(new_n209));
  AOI21_X1  g008(.A(KEYINPUT15), .B1(new_n209), .B2(new_n204), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n206), .B1(new_n210), .B2(KEYINPUT91), .ZN(new_n211));
  INV_X1    g010(.A(G29gat), .ZN(new_n212));
  INV_X1    g011(.A(G36gat), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT14), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AND3_X1   g013(.A1(new_n212), .A2(new_n213), .A3(KEYINPUT14), .ZN(new_n215));
  XNOR2_X1  g014(.A(KEYINPUT89), .B(G36gat), .ZN(new_n216));
  AOI211_X1 g015(.A(new_n214), .B(new_n215), .C1(G29gat), .C2(new_n216), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n211), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n206), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n210), .A2(KEYINPUT91), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n219), .B1(new_n220), .B2(new_n217), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G15gat), .B(G22gat), .ZN(new_n223));
  OR2_X1    g022(.A1(new_n223), .A2(G1gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT16), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n223), .B1(new_n225), .B2(G1gat), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n223), .A2(G1gat), .ZN(new_n228));
  OAI21_X1  g027(.A(G8gat), .B1(new_n228), .B2(KEYINPUT92), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n227), .B(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n202), .B1(new_n222), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n220), .A2(new_n217), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(new_n206), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n211), .A2(new_n217), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n224), .A2(new_n226), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(new_n229), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n235), .A2(KEYINPUT94), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n230), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n231), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G229gat), .A2(G233gat), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n241), .B(KEYINPUT13), .Z(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT95), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT17), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n246), .B1(new_n218), .B2(new_n221), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n233), .A2(KEYINPUT17), .A3(new_n234), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n230), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n241), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n235), .A2(new_n237), .ZN(new_n251));
  NOR3_X1   g050(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT18), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n240), .A2(KEYINPUT95), .A3(new_n242), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n245), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n252), .A2(KEYINPUT18), .ZN(new_n256));
  XNOR2_X1  g055(.A(G113gat), .B(G141gat), .ZN(new_n257));
  INV_X1    g056(.A(G197gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(KEYINPUT11), .B(G169gat), .ZN(new_n260));
  XOR2_X1   g059(.A(new_n259), .B(new_n260), .Z(new_n261));
  XNOR2_X1  g060(.A(new_n261), .B(KEYINPUT12), .ZN(new_n262));
  NOR3_X1   g061(.A1(new_n255), .A2(new_n256), .A3(new_n262), .ZN(new_n263));
  AND3_X1   g062(.A1(new_n240), .A2(KEYINPUT95), .A3(new_n242), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT95), .B1(new_n240), .B2(new_n242), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n249), .A2(new_n251), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(new_n241), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT18), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n268), .A2(KEYINPUT93), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT93), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n271), .B1(new_n252), .B2(KEYINPUT18), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n266), .A2(new_n253), .A3(new_n270), .A4(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(new_n262), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT96), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT96), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n270), .A2(new_n272), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n276), .B(new_n262), .C1(new_n277), .C2(new_n255), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n263), .B1(new_n275), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G230gat), .A2(G233gat), .ZN(new_n280));
  XOR2_X1   g079(.A(KEYINPUT97), .B(G57gat), .Z(new_n281));
  INV_X1    g080(.A(G64gat), .ZN(new_n282));
  OR3_X1    g081(.A1(new_n281), .A2(KEYINPUT98), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G71gat), .A2(G78gat), .ZN(new_n284));
  OR2_X1    g083(.A1(G71gat), .A2(G78gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT9), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n281), .A2(new_n282), .ZN(new_n288));
  INV_X1    g087(.A(G57gat), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT98), .B1(new_n289), .B2(G64gat), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n283), .B(new_n287), .C1(new_n288), .C2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G57gat), .B(G64gat), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n284), .B(new_n285), .C1(new_n292), .C2(new_n286), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(G85gat), .A2(G92gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n295), .B(KEYINPUT7), .ZN(new_n296));
  INV_X1    g095(.A(G99gat), .ZN(new_n297));
  INV_X1    g096(.A(G106gat), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT8), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n296), .B(new_n299), .C1(G85gat), .C2(G92gat), .ZN(new_n300));
  XOR2_X1   g099(.A(G99gat), .B(G106gat), .Z(new_n301));
  XNOR2_X1  g100(.A(new_n300), .B(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT102), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n294), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n302), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n291), .A2(new_n293), .A3(new_n304), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT10), .B1(new_n305), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n291), .A2(new_n293), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT10), .ZN(new_n311));
  NOR3_X1   g110(.A1(new_n310), .A2(new_n302), .A3(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n280), .B1(new_n309), .B2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G176gat), .B(G204gat), .ZN(new_n314));
  INV_X1    g113(.A(G148gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n314), .B(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(KEYINPUT103), .B(G120gat), .ZN(new_n317));
  XOR2_X1   g116(.A(new_n316), .B(new_n317), .Z(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n305), .A2(G230gat), .A3(G233gat), .A4(new_n308), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n313), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n318), .A2(KEYINPUT104), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n280), .B(KEYINPUT105), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n323), .B1(new_n309), .B2(new_n312), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n322), .B1(new_n324), .B2(new_n320), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n318), .A2(KEYINPUT104), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n327), .A2(KEYINPUT106), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(KEYINPUT106), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n321), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n279), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G113gat), .B(G120gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n333), .A2(KEYINPUT1), .ZN(new_n334));
  XNOR2_X1  g133(.A(G127gat), .B(G134gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(KEYINPUT27), .B(G183gat), .ZN(new_n337));
  INV_X1    g136(.A(G190gat), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(KEYINPUT28), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(G183gat), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT27), .B1(new_n341), .B2(KEYINPUT69), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT69), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT27), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n343), .A2(new_n344), .A3(G183gat), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n342), .A2(new_n345), .A3(new_n338), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT70), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT28), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n342), .A2(new_n345), .A3(KEYINPUT70), .A4(new_n338), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT71), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n348), .A2(KEYINPUT71), .A3(new_n349), .A4(new_n350), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n340), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G183gat), .A2(G190gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(G169gat), .A2(G176gat), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT26), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(G169gat), .A2(G176gat), .ZN(new_n361));
  OAI21_X1  g160(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NOR3_X1   g163(.A1(new_n355), .A2(new_n357), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n366), .B(KEYINPUT66), .ZN(new_n367));
  NAND3_X1  g166(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n368), .B(KEYINPUT67), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n341), .A2(new_n338), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n367), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT68), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT25), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n358), .A2(KEYINPUT23), .ZN(new_n376));
  AND2_X1   g175(.A1(new_n361), .A2(KEYINPUT23), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n376), .B1(new_n377), .B2(new_n358), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n378), .B1(new_n371), .B2(new_n372), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT65), .ZN(new_n380));
  OR2_X1    g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n366), .B1(new_n341), .B2(new_n338), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n368), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n378), .A2(new_n380), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n381), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  AOI22_X1  g184(.A1(new_n375), .A2(new_n379), .B1(new_n374), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n336), .B1(new_n365), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n353), .A2(new_n354), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(new_n339), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n389), .A2(new_n356), .A3(new_n363), .ZN(new_n390));
  INV_X1    g189(.A(new_n336), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n379), .B(KEYINPUT25), .C1(new_n372), .C2(new_n371), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n385), .A2(new_n374), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n390), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(G227gat), .A2(G233gat), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n387), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT34), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT72), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n397), .A2(KEYINPUT72), .A3(KEYINPUT34), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AND2_X1   g201(.A1(new_n387), .A2(new_n395), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n396), .B(KEYINPUT64), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT32), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT34), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n403), .A2(KEYINPUT73), .A3(new_n406), .A4(new_n404), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n387), .A2(new_n395), .A3(new_n406), .A4(new_n404), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT73), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  AND3_X1   g210(.A1(new_n402), .A2(new_n405), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n405), .B1(new_n402), .B2(new_n411), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n403), .A2(new_n404), .ZN(new_n414));
  OR2_X1    g213(.A1(new_n414), .A2(KEYINPUT33), .ZN(new_n415));
  XNOR2_X1  g214(.A(G15gat), .B(G43gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n416), .B(G71gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(new_n297), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  NOR3_X1   g218(.A1(new_n412), .A2(new_n413), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n405), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n397), .A2(KEYINPUT72), .A3(KEYINPUT34), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT72), .B1(new_n397), .B2(KEYINPUT34), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n408), .B(KEYINPUT73), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n421), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n402), .A2(new_n411), .A3(new_n405), .ZN(new_n427));
  AOI22_X1  g226(.A1(new_n426), .A2(new_n427), .B1(new_n415), .B2(new_n418), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT36), .ZN(new_n429));
  OAI22_X1  g228(.A1(new_n420), .A2(new_n428), .B1(KEYINPUT74), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n419), .B1(new_n412), .B2(new_n413), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n426), .A2(new_n415), .A3(new_n427), .A4(new_n418), .ZN(new_n432));
  XNOR2_X1  g231(.A(KEYINPUT74), .B(KEYINPUT36), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n431), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(G78gat), .B(G106gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n436), .B(G22gat), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(G228gat), .ZN(new_n439));
  INV_X1    g238(.A(G233gat), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(G155gat), .A2(G162gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n442), .B(KEYINPUT78), .ZN(new_n443));
  INV_X1    g242(.A(G155gat), .ZN(new_n444));
  INV_X1    g243(.A(G162gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n442), .A2(KEYINPUT2), .ZN(new_n447));
  XNOR2_X1  g246(.A(G141gat), .B(G148gat), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n443), .B(new_n446), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT79), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n450), .B1(new_n315), .B2(G141gat), .ZN(new_n451));
  INV_X1    g250(.A(G141gat), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n452), .A2(KEYINPUT79), .A3(G148gat), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n451), .B(new_n453), .C1(new_n452), .C2(G148gat), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n442), .B1(new_n446), .B2(KEYINPUT2), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n449), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT80), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT80), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n449), .A2(new_n459), .A3(new_n456), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(G211gat), .A2(G218gat), .ZN(new_n463));
  INV_X1    g262(.A(G211gat), .ZN(new_n464));
  INV_X1    g263(.A(G218gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT22), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(G197gat), .B(G204gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  XOR2_X1   g269(.A(new_n470), .B(KEYINPUT75), .Z(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(KEYINPUT22), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n472), .A2(new_n463), .A3(new_n466), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT29), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT3), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OR2_X1    g275(.A1(new_n457), .A2(KEYINPUT3), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n475), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n478), .B(KEYINPUT84), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n474), .B(KEYINPUT76), .ZN(new_n480));
  OAI221_X1 g279(.A(new_n441), .B1(new_n462), .B2(new_n476), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(KEYINPUT31), .B(G50gat), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n476), .B1(new_n456), .B2(new_n449), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n474), .B1(new_n475), .B2(new_n477), .ZN(new_n485));
  OAI22_X1  g284(.A1(new_n484), .A2(new_n485), .B1(new_n439), .B2(new_n440), .ZN(new_n486));
  AND3_X1   g285(.A1(new_n481), .A2(new_n483), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n483), .B1(new_n481), .B2(new_n486), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n438), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n481), .A2(new_n486), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(new_n482), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n481), .A2(new_n483), .A3(new_n486), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n437), .A3(new_n492), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(G1gat), .B(G29gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(G85gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(KEYINPUT0), .B(G57gat), .ZN(new_n497));
  XOR2_X1   g296(.A(new_n496), .B(new_n497), .Z(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(G225gat), .A2(G233gat), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n391), .B1(new_n458), .B2(new_n460), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n336), .A2(new_n457), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n504), .A2(KEYINPUT82), .A3(KEYINPUT5), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT82), .ZN(new_n506));
  INV_X1    g305(.A(new_n460), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n459), .B1(new_n449), .B2(new_n456), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n336), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n503), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n500), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT5), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n506), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT4), .ZN(new_n514));
  NOR3_X1   g313(.A1(new_n503), .A2(KEYINPUT81), .A3(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n457), .A2(KEYINPUT3), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n516), .B1(new_n461), .B2(KEYINPUT3), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n515), .B1(new_n517), .B2(new_n336), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n510), .A2(KEYINPUT4), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT81), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n520), .B1(new_n503), .B2(new_n514), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n501), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  AOI22_X1  g321(.A1(new_n505), .A2(new_n513), .B1(new_n518), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n517), .A2(new_n336), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n503), .B(new_n514), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n524), .A2(new_n512), .A3(new_n500), .A4(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n499), .B1(new_n523), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n518), .A2(new_n522), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT82), .B1(new_n504), .B2(KEYINPUT5), .ZN(new_n530));
  NOR3_X1   g329(.A1(new_n511), .A2(new_n506), .A3(new_n512), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n532), .A2(new_n498), .A3(new_n526), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT6), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n528), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT83), .ZN(new_n536));
  OAI211_X1 g335(.A(KEYINPUT6), .B(new_n499), .C1(new_n523), .C2(new_n527), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT83), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n528), .A2(new_n533), .A3(new_n538), .A4(new_n534), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G8gat), .B(G36gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(G64gat), .B(G92gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(G226gat), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n544), .A2(new_n440), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n545), .A2(KEYINPUT29), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n547), .B1(new_n365), .B2(new_n386), .ZN(new_n548));
  INV_X1    g347(.A(new_n545), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n390), .A2(new_n549), .A3(new_n394), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n548), .A2(new_n550), .A3(new_n474), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n480), .B1(new_n548), .B2(new_n550), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n543), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n480), .ZN(new_n554));
  NOR3_X1   g353(.A1(new_n365), .A2(new_n386), .A3(new_n545), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n546), .B1(new_n390), .B2(new_n394), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n548), .A2(new_n550), .A3(new_n474), .ZN(new_n558));
  INV_X1    g357(.A(new_n543), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n557), .A2(new_n558), .A3(KEYINPUT30), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n553), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT77), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n557), .A2(new_n559), .A3(new_n558), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT30), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n540), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n430), .A2(new_n435), .B1(new_n494), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT37), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n568), .B1(new_n557), .B2(new_n558), .ZN(new_n569));
  OAI21_X1  g368(.A(KEYINPUT86), .B1(new_n569), .B2(new_n559), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n557), .A2(new_n568), .A3(new_n558), .ZN(new_n571));
  OAI21_X1  g370(.A(KEYINPUT37), .B1(new_n551), .B2(new_n552), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT86), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n572), .A2(new_n573), .A3(new_n543), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n570), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  XOR2_X1   g374(.A(KEYINPUT85), .B(KEYINPUT38), .Z(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT87), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n474), .B1(new_n555), .B2(new_n556), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n554), .A2(new_n548), .A3(new_n550), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n580), .A2(new_n581), .A3(KEYINPUT37), .ZN(new_n582));
  INV_X1    g381(.A(new_n576), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n582), .A2(new_n571), .A3(new_n543), .A4(new_n583), .ZN(new_n584));
  AND4_X1   g383(.A1(new_n537), .A2(new_n535), .A3(new_n563), .A4(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n575), .A2(KEYINPUT87), .A3(new_n576), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n579), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT88), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n524), .A2(KEYINPUT39), .A3(new_n525), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT39), .B1(new_n524), .B2(new_n525), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n501), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  OAI211_X1 g390(.A(KEYINPUT39), .B(new_n500), .C1(new_n502), .C2(new_n503), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n591), .A2(new_n498), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT40), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n528), .B1(new_n593), .B2(new_n594), .ZN(new_n596));
  INV_X1    g395(.A(new_n561), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n596), .B1(new_n565), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n494), .B1(new_n595), .B2(new_n598), .ZN(new_n599));
  AND3_X1   g398(.A1(new_n587), .A2(new_n588), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n588), .B1(new_n587), .B2(new_n599), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n567), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n489), .A2(new_n493), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n431), .A2(new_n603), .A3(new_n432), .ZN(new_n604));
  OAI21_X1  g403(.A(KEYINPUT35), .B1(new_n604), .B2(new_n566), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n535), .A2(new_n537), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n597), .A2(new_n565), .ZN(new_n607));
  NOR3_X1   g406(.A1(new_n606), .A2(new_n607), .A3(KEYINPUT35), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n608), .A2(new_n603), .A3(new_n432), .A4(new_n431), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n332), .B1(new_n602), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT21), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n237), .B1(new_n310), .B2(new_n612), .ZN(new_n613));
  OR2_X1    g412(.A1(new_n613), .A2(G183gat), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(G183gat), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n294), .A2(KEYINPUT21), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n616), .B1(new_n614), .B2(new_n615), .ZN(new_n618));
  XNOR2_X1  g417(.A(G127gat), .B(G155gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(G211gat), .ZN(new_n620));
  OR3_X1    g419(.A1(new_n617), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT99), .ZN(new_n623));
  NAND2_X1  g422(.A1(G231gat), .A2(G233gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n620), .B1(new_n617), .B2(new_n618), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n621), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n625), .B1(new_n621), .B2(new_n626), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n247), .A2(new_n248), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(new_n302), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n222), .A2(new_n306), .ZN(new_n633));
  NAND3_X1  g432(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G190gat), .B(G218gat), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n636), .B(KEYINPUT100), .Z(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n635), .B(new_n638), .ZN(new_n639));
  OR2_X1    g438(.A1(new_n639), .A2(KEYINPUT101), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(KEYINPUT101), .ZN(new_n641));
  XNOR2_X1  g440(.A(G134gat), .B(G162gat), .ZN(new_n642));
  AOI21_X1  g441(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n640), .A2(new_n641), .A3(new_n644), .ZN(new_n645));
  OR2_X1    g444(.A1(new_n641), .A2(new_n644), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n611), .A2(new_n630), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n540), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(G1gat), .ZN(G1324gat));
  INV_X1    g451(.A(new_n607), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n655));
  INV_X1    g454(.A(G8gat), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n225), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n654), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT42), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  OAI211_X1 g460(.A(new_n660), .B(new_n661), .C1(new_n656), .C2(new_n654), .ZN(G1325gat));
  INV_X1    g461(.A(new_n435), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n429), .A2(KEYINPUT74), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n664), .B1(new_n431), .B2(new_n432), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  AND3_X1   g465(.A1(new_n649), .A2(G15gat), .A3(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n420), .A2(new_n428), .ZN(new_n668));
  AOI21_X1  g467(.A(G15gat), .B1(new_n649), .B2(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n667), .A2(new_n669), .ZN(G1326gat));
  NOR2_X1   g469(.A1(new_n648), .A2(new_n603), .ZN(new_n671));
  XOR2_X1   g470(.A(KEYINPUT43), .B(G22gat), .Z(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(G1327gat));
  NAND2_X1  g472(.A1(new_n566), .A2(new_n494), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n674), .B1(new_n663), .B2(new_n665), .ZN(new_n675));
  INV_X1    g474(.A(new_n601), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n587), .A2(new_n599), .A3(new_n588), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n675), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n610), .ZN(new_n679));
  OAI211_X1 g478(.A(new_n629), .B(new_n331), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  NOR4_X1   g479(.A1(new_n680), .A2(G29gat), .A3(new_n540), .A4(new_n647), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n681), .B(KEYINPUT45), .Z(new_n682));
  INV_X1    g481(.A(new_n647), .ZN(new_n683));
  OAI211_X1 g482(.A(KEYINPUT44), .B(new_n683), .C1(new_n678), .C2(new_n679), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n629), .B(KEYINPUT107), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n332), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT108), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n610), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n605), .A2(KEYINPUT108), .A3(new_n609), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n647), .B1(new_n690), .B2(new_n602), .ZN(new_n691));
  OAI211_X1 g490(.A(new_n684), .B(new_n686), .C1(new_n691), .C2(KEYINPUT44), .ZN(new_n692));
  OR3_X1    g491(.A1(new_n692), .A2(KEYINPUT109), .A3(new_n540), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT109), .B1(new_n692), .B2(new_n540), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n693), .A2(G29gat), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n682), .A2(new_n695), .ZN(G1328gat));
  NOR4_X1   g495(.A1(new_n680), .A2(new_n216), .A3(new_n647), .A4(new_n653), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT46), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n216), .B1(new_n692), .B2(new_n653), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(G1329gat));
  INV_X1    g499(.A(new_n666), .ZN(new_n701));
  OAI21_X1  g500(.A(G43gat), .B1(new_n692), .B2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT47), .ZN(new_n703));
  INV_X1    g502(.A(new_n668), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n680), .A2(new_n647), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n703), .B1(new_n705), .B2(new_n203), .ZN(new_n706));
  AND3_X1   g505(.A1(new_n702), .A2(new_n706), .A3(KEYINPUT111), .ZN(new_n707));
  AOI21_X1  g506(.A(KEYINPUT111), .B1(new_n702), .B2(new_n706), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT110), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n709), .B1(new_n705), .B2(new_n203), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n702), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n703), .B1(new_n702), .B2(KEYINPUT110), .ZN(new_n712));
  OAI22_X1  g511(.A1(new_n707), .A2(new_n708), .B1(new_n711), .B2(new_n712), .ZN(G1330gat));
  OAI21_X1  g512(.A(KEYINPUT112), .B1(new_n680), .B2(new_n647), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT112), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n611), .A2(new_n715), .A3(new_n629), .A4(new_n683), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n207), .A2(new_n208), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n717), .A2(new_n718), .A3(new_n494), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT48), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n207), .B(new_n208), .C1(new_n692), .C2(new_n603), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n720), .B1(new_n719), .B2(new_n721), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n722), .A2(new_n723), .ZN(G1331gat));
  NAND3_X1  g523(.A1(new_n279), .A2(new_n630), .A3(new_n647), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n725), .B1(new_n690), .B2(new_n602), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n330), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n650), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(new_n281), .ZN(G1332gat));
  NOR2_X1   g529(.A1(new_n727), .A2(new_n653), .ZN(new_n731));
  NOR2_X1   g530(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n732));
  AND2_X1   g531(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n734), .B1(new_n731), .B2(new_n732), .ZN(G1333gat));
  OAI21_X1  g534(.A(G71gat), .B1(new_n727), .B2(new_n701), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n727), .A2(G71gat), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n736), .B1(new_n737), .B2(new_n704), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT50), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(G1334gat));
  NAND2_X1  g539(.A1(new_n728), .A2(new_n494), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(G78gat), .ZN(G1335gat));
  INV_X1    g541(.A(new_n263), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n276), .B1(new_n273), .B2(new_n262), .ZN(new_n744));
  INV_X1    g543(.A(new_n278), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n746), .A2(new_n630), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n330), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n684), .B(new_n749), .C1(new_n691), .C2(KEYINPUT44), .ZN(new_n750));
  INV_X1    g549(.A(G85gat), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n750), .A2(new_n751), .A3(new_n540), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n605), .A2(KEYINPUT108), .A3(new_n609), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT108), .B1(new_n605), .B2(new_n609), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n683), .B(new_n747), .C1(new_n755), .C2(new_n678), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT51), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n602), .B1(new_n754), .B2(new_n753), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n758), .A2(new_n759), .A3(new_n683), .A4(new_n747), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n757), .A2(new_n650), .A3(new_n330), .A4(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n752), .B1(new_n751), .B2(new_n761), .ZN(G1336gat));
  OAI21_X1  g561(.A(G92gat), .B1(new_n750), .B2(new_n653), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT113), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n653), .A2(G92gat), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n757), .A2(new_n330), .A3(new_n760), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n765), .A2(new_n768), .A3(KEYINPUT52), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n763), .B(new_n767), .C1(new_n764), .C2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(G1337gat));
  XOR2_X1   g571(.A(KEYINPUT114), .B(G99gat), .Z(new_n773));
  OAI21_X1  g572(.A(new_n773), .B1(new_n750), .B2(new_n701), .ZN(new_n774));
  INV_X1    g573(.A(new_n773), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n757), .A2(new_n330), .A3(new_n760), .A4(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n774), .B1(new_n704), .B2(new_n776), .ZN(G1338gat));
  NOR2_X1   g576(.A1(KEYINPUT115), .A2(KEYINPUT53), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT44), .B1(new_n758), .B2(new_n683), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT44), .ZN(new_n780));
  AOI211_X1 g579(.A(new_n780), .B(new_n647), .C1(new_n602), .C2(new_n610), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n779), .A2(new_n781), .A3(new_n748), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n603), .A2(new_n298), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n778), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n757), .A2(new_n494), .A3(new_n330), .A4(new_n760), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n298), .ZN(new_n786));
  NAND2_X1  g585(.A1(KEYINPUT115), .A2(KEYINPUT53), .ZN(new_n787));
  AND3_X1   g586(.A1(new_n784), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n787), .B1(new_n784), .B2(new_n786), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n788), .A2(new_n789), .ZN(G1339gat));
  NOR2_X1   g589(.A1(new_n725), .A2(new_n330), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n793), .B(new_n323), .C1(new_n309), .C2(new_n312), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n794), .A2(new_n318), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n305), .A2(new_n308), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n311), .ZN(new_n797));
  INV_X1    g596(.A(new_n312), .ZN(new_n798));
  INV_X1    g597(.A(new_n323), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n800), .A2(KEYINPUT54), .A3(new_n313), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n795), .A2(KEYINPUT55), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n321), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT116), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n795), .A2(new_n801), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n802), .A2(KEYINPUT116), .A3(new_n321), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n805), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n261), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n267), .A2(new_n241), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n240), .A2(new_n242), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n811), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n743), .A2(new_n814), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n810), .A2(new_n647), .A3(new_n815), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n743), .A2(new_n814), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n330), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n818), .B1(new_n279), .B2(new_n810), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n816), .B1(new_n819), .B2(new_n647), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n792), .B1(new_n820), .B2(new_n685), .ZN(new_n821));
  INV_X1    g620(.A(new_n604), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n540), .A2(new_n607), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT117), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(G113gat), .B1(new_n827), .B2(new_n279), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n279), .A2(G113gat), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n828), .B1(new_n825), .B2(new_n829), .ZN(G1340gat));
  INV_X1    g629(.A(new_n330), .ZN(new_n831));
  OAI21_X1  g630(.A(G120gat), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  OR2_X1    g631(.A1(new_n831), .A2(G120gat), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n832), .B1(new_n825), .B2(new_n833), .ZN(G1341gat));
  INV_X1    g633(.A(new_n685), .ZN(new_n835));
  INV_X1    g634(.A(G127gat), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n823), .A2(new_n630), .A3(new_n824), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n826), .A2(new_n837), .B1(new_n836), .B2(new_n838), .ZN(G1342gat));
  OAI21_X1  g638(.A(G134gat), .B1(new_n827), .B2(new_n647), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n825), .A2(G134gat), .A3(new_n647), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(KEYINPUT56), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(G1343gat));
  NOR2_X1   g642(.A1(new_n666), .A2(new_n540), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n821), .A2(new_n494), .A3(new_n844), .ZN(new_n845));
  OR2_X1    g644(.A1(new_n845), .A2(KEYINPUT119), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n279), .A2(G141gat), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(KEYINPUT119), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n846), .A2(new_n653), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n821), .A2(new_n850), .A3(new_n494), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n844), .A2(new_n653), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n803), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n746), .A2(new_n808), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n683), .B1(new_n855), .B2(new_n818), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n629), .B1(new_n856), .B2(new_n816), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n603), .B1(new_n857), .B2(new_n792), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n851), .B(new_n853), .C1(new_n850), .C2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(G141gat), .B1(new_n859), .B2(new_n279), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT58), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n849), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n821), .A2(new_n494), .ZN(new_n863));
  NOR4_X1   g662(.A1(new_n863), .A2(new_n852), .A3(G141gat), .A4(new_n279), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n857), .A2(new_n792), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n494), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n852), .B1(new_n866), .B2(KEYINPUT57), .ZN(new_n867));
  AOI21_X1  g666(.A(KEYINPUT118), .B1(new_n867), .B2(new_n851), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n859), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n746), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n864), .B1(new_n871), .B2(G141gat), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n862), .B1(new_n872), .B2(new_n861), .ZN(G1344gat));
  NAND4_X1  g672(.A1(new_n846), .A2(new_n653), .A3(new_n330), .A4(new_n848), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n874), .A2(KEYINPUT59), .A3(new_n315), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n867), .A2(KEYINPUT118), .A3(new_n851), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n859), .A2(new_n869), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n831), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n856), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT120), .ZN(new_n880));
  OR3_X1    g679(.A1(new_n810), .A2(new_n647), .A3(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n880), .B1(new_n810), .B2(new_n647), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n881), .A2(new_n817), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n630), .B1(new_n879), .B2(new_n883), .ZN(new_n884));
  OR3_X1    g683(.A1(new_n884), .A2(KEYINPUT121), .A3(new_n791), .ZN(new_n885));
  OAI21_X1  g684(.A(KEYINPUT121), .B1(new_n884), .B2(new_n791), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n885), .A2(new_n850), .A3(new_n494), .A4(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n863), .A2(KEYINPUT57), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n887), .A2(new_n330), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n853), .A2(KEYINPUT59), .ZN(new_n890));
  OAI22_X1  g689(.A1(new_n878), .A2(KEYINPUT59), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n875), .B1(new_n891), .B2(G148gat), .ZN(G1345gat));
  NAND4_X1  g691(.A1(new_n846), .A2(new_n630), .A3(new_n653), .A4(new_n848), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n893), .A2(new_n444), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n868), .A2(new_n870), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n895), .A2(new_n835), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n894), .B1(new_n896), .B2(G155gat), .ZN(G1346gat));
  NAND4_X1  g696(.A1(new_n846), .A2(new_n683), .A3(new_n653), .A4(new_n848), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n898), .A2(new_n445), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n895), .A2(new_n647), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g700(.A1(new_n650), .A2(new_n653), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n821), .A2(new_n822), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n746), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n330), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(G176gat), .ZN(G1349gat));
  INV_X1    g706(.A(KEYINPUT60), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n903), .A2(new_n685), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(G183gat), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n821), .A2(new_n902), .A3(new_n337), .A4(new_n822), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n911), .A2(new_n629), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n912), .A2(KEYINPUT122), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT122), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n911), .A2(new_n914), .A3(new_n629), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n910), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n908), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n912), .B(KEYINPUT122), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT123), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n920), .A2(new_n908), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n919), .A2(KEYINPUT124), .A3(new_n910), .A4(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n916), .A2(new_n920), .ZN(new_n923));
  AND3_X1   g722(.A1(new_n918), .A2(new_n922), .A3(new_n923), .ZN(G1350gat));
  NAND2_X1  g723(.A1(new_n903), .A2(new_n683), .ZN(new_n925));
  XOR2_X1   g724(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n338), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(KEYINPUT126), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT126), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n925), .A2(new_n931), .A3(new_n928), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n927), .A2(new_n338), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n933), .B(new_n935), .ZN(G1351gat));
  INV_X1    g735(.A(new_n902), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n863), .A2(new_n666), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n938), .A2(new_n258), .A3(new_n746), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n666), .A2(new_n937), .ZN(new_n940));
  AND4_X1   g739(.A1(new_n746), .A2(new_n887), .A3(new_n888), .A4(new_n940), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n939), .B1(new_n941), .B2(new_n258), .ZN(G1352gat));
  INV_X1    g741(.A(G204gat), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n938), .A2(new_n943), .A3(new_n330), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(KEYINPUT62), .ZN(new_n945));
  OR2_X1    g744(.A1(new_n944), .A2(KEYINPUT62), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n889), .A2(new_n666), .A3(new_n937), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n945), .B(new_n946), .C1(new_n947), .C2(new_n943), .ZN(G1353gat));
  NAND4_X1  g747(.A1(new_n887), .A2(new_n630), .A3(new_n888), .A4(new_n940), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(G211gat), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n950), .A2(new_n951), .A3(KEYINPUT63), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n938), .A2(new_n464), .A3(new_n630), .ZN(new_n953));
  OR2_X1    g752(.A1(new_n951), .A2(KEYINPUT63), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n951), .A2(KEYINPUT63), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n949), .A2(G211gat), .A3(new_n954), .A4(new_n955), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n952), .A2(new_n953), .A3(new_n956), .ZN(G1354gat));
  NAND3_X1  g756(.A1(new_n938), .A2(new_n465), .A3(new_n683), .ZN(new_n958));
  AND4_X1   g757(.A1(new_n683), .A2(new_n887), .A3(new_n888), .A4(new_n940), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n958), .B1(new_n959), .B2(new_n465), .ZN(G1355gat));
endmodule


