//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 0 0 1 1 0 1 0 1 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 0 1 1 1 0 1 0 1 1 1 0 0 0 1 1 0 1 1 0 0 0 0 0 0 1 1 0 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n456, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n559, new_n561, new_n562, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n577, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n879, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  AOI22_X1  g029(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n452), .ZN(G319));
  NAND2_X1  g030(.A1(G113), .A2(G2104), .ZN(new_n456));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2104), .ZN(new_n458));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G125), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n456), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT65), .A2(G2105), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT65), .A2(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT66), .B(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n463), .A2(new_n467), .B1(new_n469), .B2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n459), .A2(KEYINPUT66), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT66), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n471), .A2(new_n473), .A3(KEYINPUT3), .ZN(new_n474));
  NAND4_X1  g049(.A1(new_n474), .A2(G137), .A3(new_n466), .A4(new_n458), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  NAND2_X1  g052(.A1(new_n474), .A2(new_n458), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n478), .A2(new_n466), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OAI221_X1 g057(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n466), .C2(G112), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n480), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  NOR3_X1   g061(.A1(new_n464), .A2(new_n465), .A3(new_n486), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n487), .A2(KEYINPUT4), .A3(new_n474), .A4(new_n458), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  OR2_X1    g064(.A1(KEYINPUT65), .A2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(KEYINPUT65), .A2(G2105), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n490), .A2(G138), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n489), .B1(new_n492), .B2(new_n461), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g069(.A1(G126), .A2(G2105), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n474), .A2(new_n458), .A3(new_n495), .ZN(new_n496));
  OR2_X1    g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(G2105), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n497), .B(G2104), .C1(G114), .C2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT67), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT67), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n496), .A2(new_n502), .A3(new_n499), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n494), .B1(new_n501), .B2(new_n503), .ZN(G164));
  NAND2_X1  g079(.A1(G75), .A2(G543), .ZN(new_n505));
  AND3_X1   g080(.A1(KEYINPUT68), .A2(KEYINPUT5), .A3(G543), .ZN(new_n506));
  AOI21_X1  g081(.A(G543), .B1(KEYINPUT68), .B2(KEYINPUT5), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G62), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n505), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n510), .A2(G651), .B1(G50), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT69), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n517), .B1(new_n508), .B2(new_n513), .ZN(new_n518));
  OAI221_X1 g093(.A(KEYINPUT69), .B1(new_n511), .B2(new_n512), .C1(new_n506), .C2(new_n507), .ZN(new_n519));
  XOR2_X1   g094(.A(KEYINPUT70), .B(G88), .Z(new_n520));
  NAND3_X1  g095(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n516), .A2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  NAND2_X1  g098(.A1(KEYINPUT68), .A2(KEYINPUT5), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(new_n514), .ZN(new_n525));
  NAND3_X1  g100(.A1(KEYINPUT68), .A2(KEYINPUT5), .A3(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(G63), .A2(G651), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n515), .A2(G51), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n518), .A2(new_n519), .ZN(new_n531));
  XOR2_X1   g106(.A(KEYINPUT71), .B(G89), .Z(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  AOI21_X1  g110(.A(KEYINPUT72), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n533), .A2(KEYINPUT72), .A3(new_n535), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n530), .B1(new_n537), .B2(new_n538), .ZN(G168));
  AOI22_X1  g114(.A1(new_n527), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(KEYINPUT73), .ZN(new_n541));
  INV_X1    g116(.A(G77), .ZN(new_n542));
  INV_X1    g117(.A(G64), .ZN(new_n543));
  OAI221_X1 g118(.A(KEYINPUT73), .B1(new_n542), .B2(new_n514), .C1(new_n508), .C2(new_n543), .ZN(new_n544));
  AND3_X1   g119(.A1(new_n541), .A2(G651), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n515), .A2(G52), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n518), .A2(new_n519), .ZN(new_n547));
  INV_X1    g122(.A(G90), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n545), .A2(new_n549), .ZN(G171));
  NAND2_X1  g125(.A1(new_n531), .A2(G81), .ZN(new_n551));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G56), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n508), .B2(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n554), .A2(G651), .B1(G43), .B2(new_n515), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  AND3_X1   g133(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G36), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(G188));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n564), .B1(new_n525), .B2(new_n526), .ZN(new_n565));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT74), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT74), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n569), .B(new_n566), .C1(new_n508), .C2(new_n564), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n570), .A3(G651), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n518), .A2(new_n519), .A3(G91), .ZN(new_n572));
  OAI211_X1 g147(.A(G53), .B(G543), .C1(new_n511), .C2(new_n512), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT9), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n571), .A2(new_n572), .A3(new_n574), .ZN(G299));
  INV_X1    g150(.A(G171), .ZN(G301));
  AND3_X1   g151(.A1(new_n533), .A2(KEYINPUT72), .A3(new_n535), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n529), .B1(new_n577), .B2(new_n536), .ZN(G286));
  INV_X1    g153(.A(G74), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n508), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(G651), .A2(new_n580), .B1(new_n515), .B2(G49), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n518), .A2(new_n519), .A3(G87), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G288));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n584), .B1(new_n525), .B2(new_n526), .ZN(new_n585));
  AND2_X1   g160(.A1(G73), .A2(G543), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT75), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n518), .A2(new_n519), .A3(G86), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n515), .A2(G48), .ZN(new_n591));
  OAI211_X1 g166(.A(KEYINPUT75), .B(G651), .C1(new_n585), .C2(new_n586), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n589), .A2(new_n590), .A3(new_n591), .A4(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(KEYINPUT76), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n593), .A2(KEYINPUT76), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n595), .A2(new_n596), .ZN(G305));
  NAND2_X1  g172(.A1(G72), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G60), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n508), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(G651), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT77), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n601), .B(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n515), .A2(G47), .ZN(new_n604));
  INV_X1    g179(.A(G85), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n547), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(G290));
  NAND3_X1  g183(.A1(new_n531), .A2(KEYINPUT10), .A3(G92), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  INV_X1    g185(.A(G92), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n547), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(G79), .A2(G543), .ZN(new_n614));
  INV_X1    g189(.A(G66), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n508), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G651), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n515), .A2(G54), .ZN(new_n618));
  AND2_X1   g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n613), .A2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(G868), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(new_n621), .B2(G171), .ZN(G284));
  OAI21_X1  g198(.A(new_n622), .B1(new_n621), .B2(G171), .ZN(G321));
  NAND2_X1  g199(.A1(G299), .A2(new_n621), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G168), .B2(new_n621), .ZN(G297));
  OAI21_X1  g201(.A(new_n625), .B1(G168), .B2(new_n621), .ZN(G280));
  INV_X1    g202(.A(new_n620), .ZN(new_n628));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(G860), .ZN(G148));
  OAI21_X1  g205(.A(KEYINPUT78), .B1(new_n557), .B2(G868), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n628), .A2(new_n629), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G868), .ZN(new_n633));
  MUX2_X1   g208(.A(KEYINPUT78), .B(new_n631), .S(new_n633), .Z(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g210(.A(KEYINPUT3), .B(G2104), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n469), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT12), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT13), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2100), .ZN(new_n640));
  OAI221_X1 g215(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n466), .C2(G111), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n481), .A2(G123), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n479), .A2(G135), .ZN(new_n643));
  AND2_X1   g218(.A1(new_n643), .A2(KEYINPUT79), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n643), .A2(KEYINPUT79), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n641), .B(new_n642), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n646), .A2(G2096), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(G2096), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n640), .A2(new_n647), .A3(new_n648), .ZN(G156));
  XNOR2_X1  g224(.A(KEYINPUT15), .B(G2435), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT81), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2427), .B(G2430), .Z(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(KEYINPUT14), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2443), .B(G2446), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n656), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2451), .B(G2454), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n661), .B(new_n662), .Z(new_n663));
  OR2_X1    g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n660), .A2(new_n663), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n664), .A2(G14), .A3(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(G401));
  XNOR2_X1  g242(.A(G2072), .B(G2078), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT17), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2067), .B(G2678), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2084), .B(G2090), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT82), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n669), .A2(new_n670), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n674), .B(new_n671), .C1(new_n668), .C2(new_n670), .ZN(new_n675));
  INV_X1    g250(.A(new_n671), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n676), .A2(new_n668), .A3(new_n670), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT18), .Z(new_n678));
  NAND3_X1  g253(.A1(new_n673), .A2(new_n675), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2096), .B(G2100), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n681), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(G227));
  XNOR2_X1  g259(.A(G1981), .B(G1986), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1956), .B(G2474), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1961), .B(G1966), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n688), .A2(KEYINPUT83), .ZN(new_n689));
  XOR2_X1   g264(.A(G1971), .B(G1976), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT19), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n688), .A2(KEYINPUT83), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n689), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT84), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT20), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n694), .A2(new_n695), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n686), .A2(new_n687), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n691), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT85), .Z(new_n700));
  NOR3_X1   g275(.A1(new_n691), .A2(new_n688), .A3(new_n698), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n696), .A2(new_n697), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g281(.A1(new_n696), .A2(new_n697), .A3(new_n702), .A4(new_n704), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(G1991), .B(G1996), .Z(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n709), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n706), .A2(new_n711), .A3(new_n707), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n685), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n710), .A2(new_n685), .A3(new_n712), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(G229));
  INV_X1    g292(.A(G16), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G20), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT23), .Z(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G299), .B2(G16), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(G1956), .ZN(new_n722));
  INV_X1    g297(.A(G29), .ZN(new_n723));
  INV_X1    g298(.A(G2084), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT24), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n725), .A2(G34), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(G34), .ZN(new_n727));
  AOI21_X1  g302(.A(G29), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n476), .B2(G29), .ZN(new_n729));
  OAI22_X1  g304(.A1(new_n646), .A2(new_n723), .B1(new_n724), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n724), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT31), .B(G11), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT30), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n733), .A2(G28), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n723), .B1(new_n733), .B2(G28), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n731), .B(new_n732), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n730), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n723), .A2(G27), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G164), .B2(new_n723), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(G2078), .Z(new_n740));
  XOR2_X1   g315(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT93), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n723), .A2(G26), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(new_n458), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n468), .B2(KEYINPUT3), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n746), .A2(G140), .A3(new_n498), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n746), .A2(G128), .A3(new_n467), .ZN(new_n748));
  OAI221_X1 g323(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n466), .C2(G116), .ZN(new_n749));
  AND3_X1   g324(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n744), .B1(new_n723), .B2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G2067), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n737), .A2(new_n740), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n723), .A2(G33), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n746), .A2(new_n498), .ZN(new_n756));
  INV_X1    g331(.A(G139), .ZN(new_n757));
  OAI21_X1  g332(.A(KEYINPUT94), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT94), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n479), .A2(new_n759), .A3(G139), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT95), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT25), .ZN(new_n763));
  NAND2_X1  g338(.A1(G103), .A2(G2104), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n467), .B2(new_n764), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n466), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n766));
  NAND2_X1  g341(.A1(G115), .A2(G2104), .ZN(new_n767));
  INV_X1    g342(.A(G127), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(new_n461), .B2(new_n768), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n765), .A2(new_n766), .B1(new_n769), .B2(new_n467), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n761), .A2(new_n762), .A3(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n762), .B1(new_n761), .B2(new_n770), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n755), .B1(new_n774), .B2(new_n723), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n754), .B1(G2072), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n718), .A2(G19), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n557), .B2(new_n718), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G1341), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n723), .A2(G32), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n481), .A2(G129), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n469), .A2(KEYINPUT97), .A3(G105), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(KEYINPUT97), .B1(new_n469), .B2(G105), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n781), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n479), .A2(G141), .ZN(new_n786));
  NAND3_X1  g361(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT26), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n780), .B1(new_n790), .B2(new_n723), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT27), .B(G1996), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n779), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n723), .A2(G35), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G162), .B2(new_n723), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT29), .Z(new_n797));
  INV_X1    g372(.A(G2090), .ZN(new_n798));
  NOR2_X1   g373(.A1(G4), .A2(G16), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(new_n628), .B2(G16), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n797), .A2(new_n798), .B1(G1348), .B2(new_n800), .ZN(new_n801));
  AND4_X1   g376(.A1(new_n722), .A2(new_n776), .A3(new_n794), .A4(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT99), .B(G1966), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(G168), .A2(G16), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n805), .A2(KEYINPUT98), .ZN(new_n806));
  OAI21_X1  g381(.A(KEYINPUT98), .B1(G16), .B2(G21), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G168), .B2(G16), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n804), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT100), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n775), .A2(G2072), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT96), .Z(new_n812));
  NOR3_X1   g387(.A1(new_n806), .A2(new_n804), .A3(new_n808), .ZN(new_n813));
  OAI22_X1  g388(.A1(new_n797), .A2(new_n798), .B1(G1348), .B2(new_n800), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n718), .A2(G5), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G171), .B2(new_n718), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G1961), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n813), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n802), .A2(new_n810), .A3(new_n812), .A4(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n718), .B1(new_n516), .B2(new_n521), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n718), .A2(G22), .ZN(new_n821));
  OR3_X1    g396(.A1(new_n820), .A2(KEYINPUT90), .A3(new_n821), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT89), .B(G1971), .Z(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(KEYINPUT90), .B1(new_n820), .B2(new_n821), .ZN(new_n825));
  AND3_X1   g400(.A1(new_n822), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n824), .B1(new_n822), .B2(new_n825), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n718), .B1(new_n581), .B2(new_n582), .ZN(new_n829));
  AND2_X1   g404(.A1(new_n718), .A2(G23), .ZN(new_n830));
  OR3_X1    g405(.A1(new_n829), .A2(KEYINPUT88), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(KEYINPUT88), .B1(new_n829), .B2(new_n830), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT33), .B(G1976), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n834), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n831), .A2(new_n836), .A3(new_n832), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  XOR2_X1   g413(.A(KEYINPUT32), .B(G1981), .Z(new_n839));
  INV_X1    g414(.A(new_n596), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n718), .B1(new_n840), .B2(new_n594), .ZN(new_n841));
  NOR2_X1   g416(.A1(G6), .A2(G16), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n839), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n839), .ZN(new_n844));
  INV_X1    g419(.A(new_n842), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n844), .B(new_n845), .C1(G305), .C2(new_n718), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n828), .A2(new_n838), .A3(new_n843), .A4(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(KEYINPUT34), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n607), .A2(new_n718), .ZN(new_n849));
  INV_X1    g424(.A(G1986), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n718), .A2(G24), .ZN(new_n851));
  OR3_X1    g426(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n850), .B1(new_n849), .B2(new_n851), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n723), .A2(G25), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT86), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n479), .A2(G131), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n481), .A2(G119), .ZN(new_n857));
  OAI221_X1 g432(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n466), .C2(G107), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT87), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n855), .B1(new_n860), .B2(new_n723), .ZN(new_n861));
  XOR2_X1   g436(.A(KEYINPUT35), .B(G1991), .Z(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n862), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n864), .B(new_n855), .C1(new_n860), .C2(new_n723), .ZN(new_n865));
  AOI22_X1  g440(.A1(new_n852), .A2(new_n853), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT91), .ZN(new_n867));
  OAI211_X1 g442(.A(new_n866), .B(new_n867), .C1(new_n847), .C2(KEYINPUT34), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n843), .A2(new_n846), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT34), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n870), .A2(new_n871), .A3(new_n838), .A4(new_n828), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n867), .B1(new_n872), .B2(new_n866), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n848), .B1(new_n869), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(KEYINPUT36), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT36), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n876), .B(new_n848), .C1(new_n869), .C2(new_n873), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n819), .B1(new_n875), .B2(new_n877), .ZN(G311));
  INV_X1    g453(.A(KEYINPUT101), .ZN(new_n879));
  XNOR2_X1  g454(.A(G311), .B(new_n879), .ZN(G150));
  NAND2_X1  g455(.A1(new_n515), .A2(G55), .ZN(new_n881));
  INV_X1    g456(.A(G651), .ZN(new_n882));
  AOI22_X1  g457(.A1(new_n527), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n883));
  INV_X1    g458(.A(G93), .ZN(new_n884));
  OAI221_X1 g459(.A(new_n881), .B1(new_n882), .B2(new_n883), .C1(new_n547), .C2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(G860), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT104), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT37), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n620), .A2(new_n629), .ZN(new_n889));
  XOR2_X1   g464(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n890));
  XNOR2_X1  g465(.A(new_n889), .B(new_n890), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n556), .B(new_n885), .Z(new_n892));
  XNOR2_X1  g467(.A(new_n891), .B(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(KEYINPUT39), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT103), .ZN(new_n895));
  INV_X1    g470(.A(G860), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n896), .B1(new_n893), .B2(KEYINPUT39), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n888), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT105), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n898), .B(new_n899), .ZN(G145));
  XNOR2_X1  g475(.A(new_n484), .B(new_n476), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n646), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n488), .A2(new_n493), .A3(new_n496), .A4(new_n499), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n750), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n904), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n790), .A2(new_n905), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n784), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(new_n782), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n911), .A2(new_n786), .A3(new_n788), .A4(new_n781), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n750), .A2(new_n904), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n906), .A2(new_n907), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT106), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n761), .A2(new_n770), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n909), .A2(new_n915), .A3(new_n916), .A4(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n909), .A2(new_n915), .A3(new_n917), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT106), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n917), .A2(KEYINPUT95), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n771), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n922), .B1(new_n909), .B2(new_n915), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n918), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n924), .A2(new_n860), .ZN(new_n925));
  INV_X1    g500(.A(new_n860), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n909), .A2(new_n915), .ZN(new_n927));
  OAI211_X1 g502(.A(KEYINPUT106), .B(new_n919), .C1(new_n927), .C2(new_n922), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n926), .B1(new_n928), .B2(new_n918), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n479), .A2(G142), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n481), .A2(G130), .ZN(new_n931));
  OAI221_X1 g506(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n466), .C2(G118), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n933), .B(new_n638), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NOR3_X1   g510(.A1(new_n925), .A2(new_n929), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n924), .A2(new_n860), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n928), .A2(new_n926), .A3(new_n918), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n934), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n903), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(G37), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n935), .B1(new_n925), .B2(new_n929), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n937), .A2(new_n934), .A3(new_n938), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n942), .A2(new_n902), .A3(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n940), .A2(new_n941), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT107), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT107), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n940), .A2(new_n947), .A3(new_n941), .A4(new_n944), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n946), .A2(new_n948), .A3(KEYINPUT40), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT40), .B1(new_n946), .B2(new_n948), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n949), .A2(new_n950), .ZN(G395));
  NAND2_X1  g526(.A1(new_n885), .A2(new_n621), .ZN(new_n952));
  INV_X1    g527(.A(G288), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n607), .B(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(G305), .A2(G303), .ZN(new_n955));
  OAI21_X1  g530(.A(G166), .B1(new_n595), .B2(new_n596), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n959), .B(KEYINPUT42), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n892), .B(new_n632), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n620), .B(G299), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT41), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n620), .A2(G299), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n620), .A2(G299), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n968), .A2(KEYINPUT41), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n966), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n964), .B1(new_n961), .B2(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n960), .B(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n952), .B1(new_n973), .B2(new_n621), .ZN(G295));
  OAI21_X1  g549(.A(new_n952), .B1(new_n973), .B2(new_n621), .ZN(G331));
  INV_X1    g550(.A(KEYINPUT44), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT109), .ZN(new_n977));
  NAND2_X1  g552(.A1(G286), .A2(G301), .ZN(new_n978));
  OAI211_X1 g553(.A(G171), .B(new_n529), .C1(new_n536), .C2(new_n577), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n978), .A2(new_n892), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n892), .B1(new_n978), .B2(new_n979), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n977), .B1(new_n982), .B2(new_n971), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n978), .A2(new_n892), .A3(new_n979), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT108), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n978), .A2(new_n979), .ZN(new_n986));
  INV_X1    g561(.A(new_n892), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT108), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n978), .A2(new_n892), .A3(new_n989), .A4(new_n979), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n985), .A2(new_n988), .A3(new_n963), .A4(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n988), .A2(new_n984), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT41), .B1(new_n968), .B2(new_n969), .ZN(new_n993));
  INV_X1    g568(.A(new_n969), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n994), .A2(new_n967), .A3(new_n965), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n992), .A2(new_n996), .A3(KEYINPUT109), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n983), .A2(new_n991), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n959), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n985), .A2(new_n990), .A3(new_n988), .ZN(new_n1001));
  AOI22_X1  g576(.A1(new_n1001), .A2(new_n996), .B1(new_n982), .B2(new_n963), .ZN(new_n1002));
  AOI21_X1  g577(.A(G37), .B1(new_n1002), .B2(new_n959), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n976), .B1(new_n1004), .B2(KEYINPUT43), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1003), .B1(new_n959), .B2(new_n1002), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1005), .B1(KEYINPUT43), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT110), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1001), .A2(new_n996), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n982), .A2(new_n963), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(new_n959), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n941), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1002), .A2(new_n959), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT43), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT43), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1000), .A2(new_n1003), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1008), .B1(new_n1017), .B2(new_n976), .ZN(new_n1018));
  AOI211_X1 g593(.A(KEYINPUT110), .B(KEYINPUT44), .C1(new_n1014), .C2(new_n1016), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1007), .B1(new_n1018), .B2(new_n1019), .ZN(G397));
  XNOR2_X1  g595(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G1384), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n904), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1022), .B1(new_n1024), .B2(KEYINPUT111), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n492), .A2(new_n489), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n466), .A2(new_n636), .A3(G138), .ZN(new_n1027));
  AOI22_X1  g602(.A1(new_n1026), .A2(new_n746), .B1(new_n1027), .B2(new_n489), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n496), .A2(new_n499), .ZN(new_n1029));
  AOI21_X1  g604(.A(G1384), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT111), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1025), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n463), .A2(new_n467), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n469), .A2(G101), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1034), .A2(G40), .A3(new_n1035), .A4(new_n475), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n907), .B(G2067), .ZN(new_n1039));
  XNOR2_X1  g614(.A(new_n1039), .B(KEYINPUT113), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1038), .B1(new_n1040), .B2(new_n790), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n1041), .B(KEYINPUT125), .ZN(new_n1042));
  INV_X1    g617(.A(G1996), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1037), .A2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g619(.A(new_n1044), .B(KEYINPUT46), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1042), .A2(new_n1045), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n1046), .B(KEYINPUT47), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n607), .A2(new_n850), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1038), .A2(new_n1048), .ZN(new_n1049));
  XOR2_X1   g624(.A(new_n1049), .B(KEYINPUT48), .Z(new_n1050));
  NAND2_X1  g625(.A1(new_n926), .A2(new_n864), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n912), .B(new_n1043), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n860), .A2(new_n862), .ZN(new_n1053));
  AND4_X1   g628(.A1(new_n1040), .A2(new_n1051), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1050), .B1(new_n1054), .B2(new_n1038), .ZN(new_n1055));
  AND4_X1   g630(.A1(new_n862), .A2(new_n1040), .A3(new_n860), .A4(new_n1052), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n907), .A2(G2067), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1037), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1047), .A2(new_n1055), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT124), .ZN(new_n1060));
  NAND2_X1  g635(.A1(G290), .A2(G1986), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1054), .A2(new_n1048), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n1037), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT63), .ZN(new_n1064));
  OAI21_X1  g639(.A(G8), .B1(new_n1024), .B2(new_n1036), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n590), .A2(new_n591), .A3(new_n587), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(G1981), .ZN(new_n1067));
  XOR2_X1   g642(.A(KEYINPUT115), .B(G1981), .Z(new_n1068));
  OAI21_X1  g643(.A(new_n1067), .B1(new_n593), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT49), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1065), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1067), .B(KEYINPUT49), .C1(new_n593), .C2(new_n1068), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT116), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1071), .A2(KEYINPUT116), .A3(new_n1072), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  XOR2_X1   g652(.A(KEYINPUT114), .B(G1971), .Z(new_n1078));
  OAI21_X1  g653(.A(new_n1021), .B1(G164), .B2(G1384), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1036), .B1(new_n1030), .B2(KEYINPUT45), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1078), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n496), .A2(new_n502), .A3(new_n499), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n502), .B1(new_n496), .B2(new_n499), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1028), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT50), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1084), .A2(new_n1085), .A3(new_n1023), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1036), .B1(new_n1024), .B2(KEYINPUT50), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1086), .A2(new_n1087), .A3(new_n798), .ZN(new_n1088));
  OAI21_X1  g663(.A(G8), .B1(new_n1081), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(G303), .A2(G8), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT55), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n1090), .B(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1089), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1085), .B1(new_n1084), .B2(new_n1023), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n904), .A2(new_n1085), .A3(new_n1023), .ZN(new_n1096));
  AND4_X1   g671(.A1(G40), .A2(new_n1034), .A3(new_n475), .A4(new_n1035), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n1095), .A2(G2090), .A3(new_n1098), .ZN(new_n1099));
  OAI211_X1 g674(.A(G8), .B(new_n1092), .C1(new_n1099), .C2(new_n1081), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1065), .ZN(new_n1101));
  INV_X1    g676(.A(G1976), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT52), .B1(G288), .B2(new_n1102), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1101), .B(new_n1103), .C1(new_n1102), .C2(G288), .ZN(new_n1104));
  NOR2_X1   g679(.A1(G288), .A2(new_n1102), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT52), .B1(new_n1065), .B2(new_n1105), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1077), .A2(new_n1094), .A3(new_n1100), .A4(new_n1107), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n1095), .A2(G2084), .A3(new_n1098), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1084), .A2(new_n1023), .A3(new_n1022), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT45), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1036), .B1(new_n1024), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n804), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g688(.A(G168), .B(G8), .C1(new_n1109), .C2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1064), .B1(new_n1108), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT118), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1114), .A2(new_n1064), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1078), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1022), .B1(new_n1084), .B2(new_n1023), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1097), .B1(new_n1024), .B2(new_n1111), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1118), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1036), .B1(new_n1030), .B2(new_n1085), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1122), .A2(new_n1123), .A3(new_n798), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1121), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(G8), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(new_n1093), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1117), .A2(new_n1127), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1071), .A2(KEYINPUT116), .A3(new_n1072), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT116), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1107), .B(new_n1100), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1116), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n803), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1122), .A2(new_n1123), .A3(new_n724), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1136), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1092), .B1(new_n1125), .B2(G8), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1140), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1139), .A2(new_n1141), .A3(KEYINPUT118), .A4(new_n1100), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1115), .A2(new_n1132), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1100), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n593), .A2(new_n1068), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1146), .B(KEYINPUT117), .ZN(new_n1147));
  NOR2_X1   g722(.A1(G288), .A2(G1976), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1147), .B1(new_n1077), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1145), .B1(new_n1149), .B2(new_n1065), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT53), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1152), .A2(G2078), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1033), .A2(new_n1080), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(G1961), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1155), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n1119), .A2(new_n1120), .A3(G2078), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1154), .B(new_n1156), .C1(new_n1157), .C2(KEYINPUT53), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(G171), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1152), .B1(new_n1160), .B2(G2078), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1110), .A2(new_n1112), .A3(new_n1153), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1161), .A2(G301), .A3(new_n1156), .A4(new_n1162), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1159), .A2(new_n1163), .A3(KEYINPUT54), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1164), .A2(new_n1108), .ZN(new_n1165));
  NAND2_X1  g740(.A1(G286), .A2(G8), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(new_n1136), .ZN(new_n1168));
  OAI21_X1  g743(.A(G8), .B1(new_n1109), .B2(new_n1113), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n1166), .ZN(new_n1170));
  AOI21_X1  g745(.A(KEYINPUT51), .B1(new_n1170), .B2(KEYINPUT122), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT122), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT51), .ZN(new_n1173));
  AOI211_X1 g748(.A(new_n1172), .B(new_n1173), .C1(new_n1169), .C2(new_n1166), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1168), .B1(new_n1171), .B2(new_n1174), .ZN(new_n1175));
  OAI211_X1 g750(.A(new_n1156), .B(new_n1162), .C1(new_n1157), .C2(KEYINPUT53), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(G171), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1161), .A2(G301), .A3(new_n1156), .A4(new_n1154), .ZN(new_n1178));
  AOI21_X1  g753(.A(KEYINPUT54), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1165), .A2(new_n1175), .A3(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT57), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(KEYINPUT119), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n571), .A2(new_n572), .A3(new_n574), .A4(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1182), .A2(KEYINPUT119), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n1184), .B(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g761(.A(KEYINPUT56), .B(G2072), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1187), .ZN(new_n1188));
  NOR3_X1   g763(.A1(new_n1119), .A2(new_n1120), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g764(.A(G1956), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1186), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NOR3_X1   g766(.A1(new_n1189), .A2(new_n1190), .A3(new_n1186), .ZN(new_n1192));
  AOI21_X1  g767(.A(G1348), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1030), .A2(new_n1097), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1194), .A2(G2067), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n628), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1191), .B1(new_n1192), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1197), .A2(KEYINPUT120), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT120), .ZN(new_n1199));
  OAI211_X1 g774(.A(new_n1199), .B(new_n1191), .C1(new_n1192), .C2(new_n1196), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT61), .ZN(new_n1202));
  INV_X1    g777(.A(new_n1185), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n1184), .B(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1205));
  INV_X1    g780(.A(G1956), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1079), .A2(new_n1080), .A3(new_n1187), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1204), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1202), .B1(new_n1192), .B2(new_n1209), .ZN(new_n1210));
  NOR3_X1   g785(.A1(new_n1193), .A2(new_n628), .A3(new_n1195), .ZN(new_n1211));
  INV_X1    g786(.A(G1348), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1212), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1213));
  INV_X1    g788(.A(new_n1195), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n620), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g790(.A(KEYINPUT60), .B1(new_n1211), .B2(new_n1215), .ZN(new_n1216));
  NOR2_X1   g791(.A1(new_n620), .A2(KEYINPUT60), .ZN(new_n1217));
  NAND3_X1  g792(.A1(new_n1213), .A2(new_n1217), .A3(new_n1214), .ZN(new_n1218));
  NAND3_X1  g793(.A1(new_n1207), .A2(new_n1204), .A3(new_n1208), .ZN(new_n1219));
  NAND3_X1  g794(.A1(new_n1191), .A2(new_n1219), .A3(KEYINPUT61), .ZN(new_n1220));
  AND4_X1   g795(.A1(new_n1210), .A2(new_n1216), .A3(new_n1218), .A4(new_n1220), .ZN(new_n1221));
  NAND3_X1  g796(.A1(new_n1079), .A2(new_n1080), .A3(new_n1043), .ZN(new_n1222));
  INV_X1    g797(.A(KEYINPUT121), .ZN(new_n1223));
  XOR2_X1   g798(.A(KEYINPUT58), .B(G1341), .Z(new_n1224));
  AOI22_X1  g799(.A1(new_n1222), .A2(new_n1223), .B1(new_n1194), .B2(new_n1224), .ZN(new_n1225));
  NAND4_X1  g800(.A1(new_n1079), .A2(new_n1080), .A3(KEYINPUT121), .A4(new_n1043), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1227), .A2(new_n557), .ZN(new_n1228));
  NAND2_X1  g803(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1229));
  INV_X1    g804(.A(KEYINPUT59), .ZN(new_n1230));
  NAND3_X1  g805(.A1(new_n1227), .A2(new_n1230), .A3(new_n557), .ZN(new_n1231));
  NAND2_X1  g806(.A1(new_n1229), .A2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g807(.A(new_n1201), .B1(new_n1221), .B2(new_n1232), .ZN(new_n1233));
  OAI211_X1 g808(.A(new_n1143), .B(new_n1151), .C1(new_n1181), .C2(new_n1233), .ZN(new_n1234));
  INV_X1    g809(.A(KEYINPUT123), .ZN(new_n1235));
  INV_X1    g810(.A(new_n1168), .ZN(new_n1236));
  OAI211_X1 g811(.A(KEYINPUT122), .B(G8), .C1(new_n1136), .C2(G286), .ZN(new_n1237));
  NAND2_X1  g812(.A1(new_n1237), .A2(new_n1173), .ZN(new_n1238));
  INV_X1    g813(.A(G8), .ZN(new_n1239));
  AOI21_X1  g814(.A(new_n1239), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1240));
  OAI211_X1 g815(.A(KEYINPUT122), .B(KEYINPUT51), .C1(new_n1240), .C2(new_n1167), .ZN(new_n1241));
  AOI21_X1  g816(.A(new_n1236), .B1(new_n1238), .B2(new_n1241), .ZN(new_n1242));
  INV_X1    g817(.A(KEYINPUT62), .ZN(new_n1243));
  OAI21_X1  g818(.A(new_n1235), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  AND2_X1   g819(.A1(new_n1176), .A2(G171), .ZN(new_n1245));
  NAND4_X1  g820(.A1(new_n1141), .A2(new_n1245), .A3(new_n1094), .A4(new_n1100), .ZN(new_n1246));
  AOI21_X1  g821(.A(new_n1246), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1247));
  NAND3_X1  g822(.A1(new_n1175), .A2(KEYINPUT123), .A3(KEYINPUT62), .ZN(new_n1248));
  AND3_X1   g823(.A1(new_n1244), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  OAI211_X1 g824(.A(new_n1060), .B(new_n1063), .C1(new_n1234), .C2(new_n1249), .ZN(new_n1250));
  INV_X1    g825(.A(new_n1250), .ZN(new_n1251));
  AND2_X1   g826(.A1(new_n1132), .A2(new_n1142), .ZN(new_n1252));
  AOI21_X1  g827(.A(new_n1150), .B1(new_n1252), .B2(new_n1115), .ZN(new_n1253));
  NOR3_X1   g828(.A1(new_n1164), .A2(new_n1108), .A3(new_n1179), .ZN(new_n1254));
  NAND4_X1  g829(.A1(new_n1210), .A2(new_n1216), .A3(new_n1220), .A4(new_n1218), .ZN(new_n1255));
  AOI21_X1  g830(.A(new_n1255), .B1(new_n1229), .B2(new_n1231), .ZN(new_n1256));
  OAI211_X1 g831(.A(new_n1254), .B(new_n1175), .C1(new_n1256), .C2(new_n1201), .ZN(new_n1257));
  NAND3_X1  g832(.A1(new_n1244), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1258));
  NAND3_X1  g833(.A1(new_n1253), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1259));
  AOI21_X1  g834(.A(new_n1060), .B1(new_n1259), .B2(new_n1063), .ZN(new_n1260));
  OAI21_X1  g835(.A(new_n1059), .B1(new_n1251), .B2(new_n1260), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g836(.A1(new_n946), .A2(new_n948), .ZN(new_n1263));
  NAND3_X1  g837(.A1(new_n682), .A2(G319), .A3(new_n683), .ZN(new_n1264));
  INV_X1    g838(.A(KEYINPUT126), .ZN(new_n1265));
  OAI21_X1  g839(.A(new_n666), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g840(.A(new_n1266), .B1(new_n1265), .B2(new_n1264), .ZN(new_n1267));
  INV_X1    g841(.A(new_n715), .ZN(new_n1268));
  OAI21_X1  g842(.A(new_n1267), .B1(new_n1268), .B2(new_n713), .ZN(new_n1269));
  INV_X1    g843(.A(KEYINPUT127), .ZN(new_n1270));
  NAND2_X1  g844(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g845(.A1(new_n716), .A2(KEYINPUT127), .A3(new_n1267), .ZN(new_n1272));
  NAND2_X1  g846(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g847(.A1(new_n1263), .A2(new_n1017), .A3(new_n1273), .ZN(G225));
  INV_X1    g848(.A(G225), .ZN(G308));
endmodule


