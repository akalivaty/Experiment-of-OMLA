//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 1 1 0 0 0 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT22), .ZN(new_n203));
  INV_X1    g002(.A(G211gat), .ZN(new_n204));
  INV_X1    g003(.A(G218gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n202), .A2(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(G211gat), .B(G218gat), .Z(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT71), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n207), .A2(KEYINPUT71), .A3(new_n208), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n207), .A2(new_n208), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT72), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n213), .A2(KEYINPUT72), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n211), .B(new_n212), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220));
  OAI221_X1 g019(.A(new_n218), .B1(new_n219), .B2(KEYINPUT24), .C1(new_n220), .C2(KEYINPUT23), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(KEYINPUT24), .ZN(new_n222));
  INV_X1    g021(.A(G183gat), .ZN(new_n223));
  INV_X1    g022(.A(G190gat), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n221), .A2(new_n225), .ZN(new_n226));
  XOR2_X1   g025(.A(KEYINPUT64), .B(G169gat), .Z(new_n227));
  XOR2_X1   g026(.A(KEYINPUT65), .B(G176gat), .Z(new_n228));
  NAND3_X1  g027(.A1(new_n227), .A2(new_n228), .A3(KEYINPUT23), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT25), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n220), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT23), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT25), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NOR3_X1   g032(.A1(new_n221), .A2(new_n225), .A3(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT27), .B(G183gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(new_n224), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT28), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n235), .A2(KEYINPUT28), .A3(new_n224), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT26), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n231), .A2(new_n241), .A3(new_n218), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n219), .B1(new_n231), .B2(new_n241), .ZN(new_n243));
  OR2_X1    g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  OAI22_X1  g043(.A1(new_n230), .A2(new_n234), .B1(new_n240), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(G226gat), .A2(G233gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(KEYINPUT73), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT29), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n245), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n246), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n217), .B(new_n248), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(G8gat), .B(G36gat), .Z(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(KEYINPUT74), .ZN(new_n255));
  XNOR2_X1  g054(.A(G64gat), .B(G92gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n247), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n250), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n245), .A2(new_n252), .ZN(new_n260));
  AND2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n253), .B(new_n257), .C1(new_n261), .C2(new_n217), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT75), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT30), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT30), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n262), .A2(new_n263), .A3(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n257), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n261), .A2(new_n217), .ZN(new_n269));
  INV_X1    g068(.A(new_n253), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n265), .A2(new_n267), .A3(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G113gat), .B(G120gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n273), .A2(KEYINPUT1), .ZN(new_n274));
  INV_X1    g073(.A(G127gat), .ZN(new_n275));
  INV_X1    g074(.A(G134gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(G127gat), .A2(G134gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  AND2_X1   g080(.A1(G155gat), .A2(G162gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(G155gat), .A2(G162gat), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT2), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G141gat), .B(G148gat), .ZN(new_n287));
  OR3_X1    g086(.A1(new_n284), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n284), .B1(new_n286), .B2(new_n287), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT66), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n273), .B(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT67), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n277), .A2(KEYINPUT67), .A3(new_n278), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT1), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT68), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n293), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n298), .B1(new_n293), .B2(new_n297), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n281), .B(new_n291), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT4), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT80), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n301), .ZN(new_n305));
  XOR2_X1   g104(.A(KEYINPUT76), .B(KEYINPUT4), .Z(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n301), .A2(KEYINPUT80), .A3(KEYINPUT4), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n304), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT5), .ZN(new_n310));
  NAND2_X1  g109(.A1(G225gat), .A2(G233gat), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n290), .A2(KEYINPUT3), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT3), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n314), .B1(new_n288), .B2(new_n289), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n281), .B1(new_n299), .B2(new_n300), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n312), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n309), .A2(new_n310), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n293), .A2(new_n297), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT68), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n293), .A2(new_n297), .A3(new_n298), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n280), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n323), .A2(KEYINPUT4), .A3(new_n291), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n301), .A2(new_n306), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n318), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n326), .B(KEYINPUT77), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n323), .A2(new_n291), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n312), .B1(new_n328), .B2(new_n305), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT78), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT78), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n331), .B(new_n312), .C1(new_n328), .C2(new_n305), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n330), .A2(KEYINPUT5), .A3(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n319), .B1(new_n327), .B2(new_n333), .ZN(new_n334));
  XOR2_X1   g133(.A(G1gat), .B(G29gat), .Z(new_n335));
  XNOR2_X1  g134(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n335), .B(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G57gat), .B(G85gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n337), .B(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n334), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT6), .ZN(new_n341));
  INV_X1    g140(.A(new_n339), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n342), .B(new_n319), .C1(new_n327), .C2(new_n333), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n340), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n334), .A2(KEYINPUT6), .A3(new_n339), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n272), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G78gat), .B(G106gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT31), .B(G50gat), .ZN(new_n348));
  XOR2_X1   g147(.A(new_n347), .B(new_n348), .Z(new_n349));
  XOR2_X1   g148(.A(new_n349), .B(KEYINPUT81), .Z(new_n350));
  INV_X1    g149(.A(new_n217), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n351), .B1(KEYINPUT29), .B2(new_n313), .ZN(new_n352));
  OAI21_X1  g151(.A(KEYINPUT82), .B1(new_n215), .B2(new_n216), .ZN(new_n353));
  OR2_X1    g152(.A1(new_n207), .A2(new_n208), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT72), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT82), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n356), .A2(new_n357), .A3(new_n214), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n353), .A2(new_n209), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT3), .B1(new_n359), .B2(new_n249), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n352), .B1(new_n360), .B2(new_n291), .ZN(new_n361));
  INV_X1    g160(.A(G228gat), .ZN(new_n362));
  INV_X1    g161(.A(G233gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT83), .B(G22gat), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n314), .B1(new_n351), .B2(KEYINPUT29), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(new_n290), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n369), .A2(new_n364), .A3(new_n352), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n366), .A2(new_n367), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n367), .B1(new_n366), .B2(new_n370), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n350), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n366), .A2(new_n370), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(G22gat), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n366), .A2(new_n367), .A3(new_n370), .ZN(new_n376));
  INV_X1    g175(.A(new_n349), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n230), .ZN(new_n380));
  INV_X1    g179(.A(new_n234), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OR2_X1    g181(.A1(new_n240), .A2(new_n244), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n317), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n323), .A2(new_n245), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT34), .ZN(new_n387));
  INV_X1    g186(.A(G227gat), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n386), .B(new_n387), .C1(new_n388), .C2(new_n363), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n388), .A2(new_n363), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT69), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n390), .B1(new_n386), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n384), .A2(new_n385), .A3(KEYINPUT69), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT70), .B1(new_n394), .B2(KEYINPUT34), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT70), .ZN(new_n396));
  AOI211_X1 g195(.A(new_n396), .B(new_n387), .C1(new_n392), .C2(new_n393), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n389), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G15gat), .B(G43gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(G71gat), .B(G99gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n399), .B(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n385), .A3(new_n390), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT33), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(KEYINPUT32), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n402), .B(KEYINPUT32), .C1(new_n403), .C2(new_n401), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n398), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n408), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n410), .B(new_n389), .C1(new_n395), .C2(new_n397), .ZN(new_n411));
  AND3_X1   g210(.A1(new_n409), .A2(KEYINPUT36), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT36), .B1(new_n409), .B2(new_n411), .ZN(new_n413));
  OAI22_X1  g212(.A1(new_n346), .A2(new_n379), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT38), .ZN(new_n415));
  XOR2_X1   g214(.A(KEYINPUT85), .B(KEYINPUT37), .Z(new_n416));
  OAI211_X1 g215(.A(new_n253), .B(new_n416), .C1(new_n261), .C2(new_n217), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n417), .A2(new_n268), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT37), .B1(new_n269), .B2(new_n270), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n415), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n261), .A2(new_n351), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n248), .B1(new_n251), .B2(new_n252), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT37), .B1(new_n422), .B2(new_n217), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n415), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n417), .A2(new_n268), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n262), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n420), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n344), .A2(new_n427), .A3(new_n345), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n316), .A2(new_n317), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n311), .B1(new_n309), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT39), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n339), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n317), .A2(new_n290), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n433), .A2(new_n311), .A3(new_n301), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT39), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT84), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n435), .B(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n432), .B1(new_n430), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT40), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n432), .B(KEYINPUT40), .C1(new_n430), .C2(new_n437), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n440), .A2(new_n441), .A3(new_n340), .A4(new_n272), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n428), .A2(new_n442), .A3(new_n379), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT86), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT86), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n428), .A2(new_n442), .A3(new_n445), .A4(new_n379), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n414), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n379), .A2(new_n409), .A3(new_n411), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT35), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n448), .A2(new_n346), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n449), .B1(new_n448), .B2(new_n346), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n447), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g252(.A(G15gat), .B(G22gat), .Z(new_n454));
  INV_X1    g253(.A(G1gat), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(G8gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(G15gat), .B(G22gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n455), .A2(KEYINPUT16), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n456), .A2(new_n457), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n457), .B1(new_n456), .B2(new_n460), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(G29gat), .ZN(new_n464));
  INV_X1    g263(.A(G36gat), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT90), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT90), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n467), .B1(G29gat), .B2(G36gat), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT14), .ZN(new_n469));
  INV_X1    g268(.A(G43gat), .ZN(new_n470));
  INV_X1    g269(.A(G50gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT15), .ZN(new_n473));
  NAND2_X1  g272(.A1(G43gat), .A2(G50gat), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(G29gat), .A2(G36gat), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT14), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n467), .B(new_n477), .C1(G29gat), .C2(G36gat), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n469), .A2(new_n475), .A3(new_n476), .A4(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n474), .ZN(new_n480));
  NOR2_X1   g279(.A1(G43gat), .A2(G50gat), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT89), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT89), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n472), .A2(new_n483), .A3(new_n474), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n482), .A2(KEYINPUT15), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n479), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n472), .A2(new_n474), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n473), .B1(new_n487), .B2(KEYINPUT89), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n478), .A2(new_n476), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n488), .A2(new_n489), .A3(new_n484), .A4(new_n469), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT17), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n486), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n463), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n486), .A2(new_n490), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT91), .B1(new_n494), .B2(KEYINPUT17), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT91), .ZN(new_n496));
  AOI211_X1 g295(.A(new_n496), .B(new_n491), .C1(new_n486), .C2(new_n490), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n493), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n463), .A2(new_n494), .ZN(new_n499));
  NAND2_X1  g298(.A1(G229gat), .A2(G233gat), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n498), .A2(KEYINPUT18), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT92), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n463), .B(new_n494), .ZN(new_n505));
  XOR2_X1   g304(.A(new_n500), .B(KEYINPUT13), .Z(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n503), .A2(new_n504), .A3(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(G113gat), .B(G141gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(KEYINPUT87), .B(G197gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n509), .B(new_n510), .ZN(new_n511));
  XOR2_X1   g310(.A(KEYINPUT11), .B(G169gat), .Z(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  XOR2_X1   g312(.A(KEYINPUT88), .B(KEYINPUT12), .Z(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n508), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n503), .A2(new_n507), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT18), .B1(new_n498), .B2(new_n502), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n508), .B(new_n515), .C1(new_n517), .C2(new_n518), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n453), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT93), .ZN(new_n525));
  NOR2_X1   g324(.A1(G71gat), .A2(G78gat), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(G71gat), .A2(G78gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(G57gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(G64gat), .ZN(new_n531));
  INV_X1    g330(.A(G64gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(G57gat), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n528), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n535), .A2(KEYINPUT9), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n525), .B(new_n529), .C1(new_n534), .C2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT9), .ZN(new_n538));
  AOI22_X1  g337(.A1(new_n531), .A2(new_n533), .B1(new_n538), .B2(new_n528), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n527), .A2(KEYINPUT93), .A3(new_n528), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n525), .B1(new_n535), .B2(new_n526), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  XOR2_X1   g342(.A(KEYINPUT94), .B(KEYINPUT21), .Z(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G231gat), .A2(G233gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(G127gat), .B(G155gat), .Z(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT20), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n547), .B(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(G183gat), .B(G211gat), .Z(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n543), .ZN(new_n553));
  AOI211_X1 g352(.A(new_n462), .B(new_n461), .C1(KEYINPUT21), .C2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n552), .B(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT10), .ZN(new_n558));
  NAND2_X1  g357(.A1(G85gat), .A2(G92gat), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT7), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT8), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n562), .B1(G99gat), .B2(G106gat), .ZN(new_n563));
  NOR2_X1   g362(.A1(G85gat), .A2(G92gat), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT97), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G99gat), .A2(G106gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT8), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT97), .ZN(new_n568));
  INV_X1    g367(.A(G85gat), .ZN(new_n569));
  INV_X1    g368(.A(G92gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n567), .A2(new_n568), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n561), .B1(new_n565), .B2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G99gat), .B(G106gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n559), .B(KEYINPUT7), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n567), .A2(new_n568), .A3(new_n571), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n568), .B1(new_n567), .B2(new_n571), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n574), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n575), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(new_n543), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT98), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g384(.A(KEYINPUT98), .B(new_n576), .C1(new_n577), .C2(new_n578), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT99), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n574), .B(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  AOI22_X1  g388(.A1(new_n573), .A2(new_n574), .B1(new_n537), .B2(new_n542), .ZN(new_n590));
  AND3_X1   g389(.A1(new_n589), .A2(KEYINPUT100), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(KEYINPUT100), .B1(new_n589), .B2(new_n590), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n558), .B(new_n583), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  NOR3_X1   g392(.A1(new_n582), .A2(new_n558), .A3(new_n543), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(G230gat), .A2(G233gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G120gat), .B(G148gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(G176gat), .B(G204gat), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n599), .B(new_n600), .Z(new_n601));
  INV_X1    g400(.A(new_n583), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n588), .B1(new_n573), .B2(KEYINPUT98), .ZN(new_n603));
  INV_X1    g402(.A(new_n586), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n590), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT100), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n589), .A2(KEYINPUT100), .A3(new_n590), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n602), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI211_X1 g408(.A(new_n598), .B(new_n601), .C1(new_n609), .C2(new_n597), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT101), .ZN(new_n611));
  INV_X1    g410(.A(new_n601), .ZN(new_n612));
  INV_X1    g411(.A(new_n597), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n613), .B1(new_n593), .B2(new_n595), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n609), .A2(new_n597), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n612), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n610), .A2(new_n611), .A3(new_n616), .ZN(new_n617));
  OAI211_X1 g416(.A(KEYINPUT101), .B(new_n612), .C1(new_n614), .C2(new_n615), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G232gat), .A2(G233gat), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n621), .A2(KEYINPUT41), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT96), .ZN(new_n623));
  XNOR2_X1  g422(.A(G134gat), .B(G162gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n582), .A2(new_n492), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n494), .A2(KEYINPUT17), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n496), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n494), .A2(KEYINPUT91), .A3(KEYINPUT17), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n627), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(G190gat), .B(G218gat), .Z(new_n632));
  NAND2_X1  g431(.A1(new_n621), .A2(KEYINPUT41), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n633), .B1(new_n582), .B2(new_n494), .ZN(new_n634));
  NOR3_X1   g433(.A1(new_n631), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n632), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n492), .B(new_n582), .C1(new_n495), .C2(new_n497), .ZN(new_n637));
  INV_X1    g436(.A(new_n634), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n626), .B1(new_n635), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n632), .B1(new_n631), .B2(new_n634), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n637), .A2(new_n636), .A3(new_n638), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n641), .A2(new_n625), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n557), .A2(new_n619), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n524), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n344), .A2(new_n345), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT102), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n344), .A2(KEYINPUT102), .A3(new_n345), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n647), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(new_n455), .ZN(G1324gat));
  INV_X1    g454(.A(new_n272), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n647), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(KEYINPUT16), .B(G8gat), .Z(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT42), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n657), .A2(new_n457), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n661), .A2(KEYINPUT103), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(KEYINPUT103), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n660), .A2(new_n662), .A3(new_n663), .ZN(G1325gat));
  NOR2_X1   g463(.A1(new_n412), .A2(new_n413), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(G15gat), .B1(new_n647), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n409), .A2(new_n411), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n668), .A2(G15gat), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n667), .B1(new_n647), .B2(new_n669), .ZN(G1326gat));
  INV_X1    g469(.A(new_n379), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n524), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(new_n646), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT43), .B(G22gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(G1327gat));
  OAI21_X1  g475(.A(new_n645), .B1(new_n447), .B2(new_n452), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n557), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n680), .A2(new_n523), .A3(new_n619), .ZN(new_n681));
  OAI211_X1 g480(.A(KEYINPUT44), .B(new_n645), .C1(new_n447), .C2(new_n452), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n679), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(G29gat), .B1(new_n683), .B2(new_n653), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT45), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n444), .A2(new_n446), .ZN(new_n686));
  INV_X1    g485(.A(new_n414), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n452), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n690), .A2(new_n645), .A3(new_n681), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n652), .A2(new_n464), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n685), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OR3_X1    g492(.A1(new_n691), .A2(new_n685), .A3(new_n692), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n684), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT104), .Z(G1328gat));
  NOR3_X1   g495(.A1(new_n691), .A2(G36gat), .A3(new_n656), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT46), .ZN(new_n698));
  OAI21_X1  g497(.A(G36gat), .B1(new_n683), .B2(new_n656), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(G1329gat));
  OAI21_X1  g499(.A(new_n470), .B1(new_n691), .B2(new_n668), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n665), .A2(G43gat), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n701), .B1(new_n683), .B2(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g503(.A(G50gat), .B1(new_n683), .B2(new_n379), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT48), .B1(new_n705), .B2(KEYINPUT105), .ZN(new_n706));
  INV_X1    g505(.A(new_n619), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n557), .A2(new_n471), .A3(new_n645), .A4(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n705), .B1(new_n672), .B2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n706), .B(new_n709), .ZN(G1331gat));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n680), .A2(new_n523), .A3(new_n644), .A4(new_n619), .ZN(new_n712));
  OR3_X1    g511(.A1(new_n453), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n711), .B1(new_n453), .B2(new_n712), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n715), .A2(new_n653), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(new_n530), .ZN(G1332gat));
  NOR2_X1   g516(.A1(new_n715), .A2(new_n656), .ZN(new_n718));
  NOR2_X1   g517(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n719));
  AND2_X1   g518(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n721), .B1(new_n718), .B2(new_n719), .ZN(G1333gat));
  INV_X1    g521(.A(G71gat), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n666), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n713), .A2(new_n714), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(KEYINPUT107), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n713), .A2(new_n727), .A3(new_n714), .A4(new_n724), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n723), .B1(new_n715), .B2(new_n668), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT50), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT50), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n729), .A2(new_n733), .A3(new_n730), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(G1334gat));
  NOR2_X1   g534(.A1(new_n715), .A2(new_n379), .ZN(new_n736));
  XNOR2_X1  g535(.A(KEYINPUT108), .B(G78gat), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1335gat));
  NOR3_X1   g537(.A1(new_n680), .A2(new_n707), .A3(new_n522), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n679), .A2(new_n682), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT109), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT109), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n679), .A2(new_n742), .A3(new_n682), .A4(new_n739), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n741), .A2(new_n652), .A3(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n680), .A2(new_n522), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n690), .A2(KEYINPUT51), .A3(new_n645), .A4(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT110), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n645), .B(new_n745), .C1(new_n447), .C2(new_n452), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT51), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n746), .A2(new_n747), .A3(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n748), .A2(KEYINPUT110), .A3(new_n749), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n652), .A2(new_n569), .A3(new_n619), .ZN(new_n754));
  OAI22_X1  g553(.A1(new_n744), .A2(new_n569), .B1(new_n753), .B2(new_n754), .ZN(G1336gat));
  INV_X1    g554(.A(KEYINPUT52), .ZN(new_n756));
  OAI21_X1  g555(.A(G92gat), .B1(new_n740), .B2(new_n656), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n707), .A2(G92gat), .A3(new_n656), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n756), .B(new_n757), .C1(new_n753), .C2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n761));
  AOI211_X1 g560(.A(new_n761), .B(new_n759), .C1(new_n746), .C2(new_n750), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n750), .ZN(new_n763));
  AOI21_X1  g562(.A(KEYINPUT111), .B1(new_n763), .B2(new_n758), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n741), .A2(new_n272), .A3(new_n743), .ZN(new_n765));
  AOI211_X1 g564(.A(new_n762), .B(new_n764), .C1(new_n765), .C2(G92gat), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n760), .B1(new_n766), .B2(new_n756), .ZN(G1337gat));
  NAND3_X1  g566(.A1(new_n741), .A2(new_n665), .A3(new_n743), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(G99gat), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n668), .A2(new_n707), .A3(G99gat), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(KEYINPUT112), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n753), .B2(new_n771), .ZN(G1338gat));
  NOR3_X1   g571(.A1(new_n707), .A2(G106gat), .A3(new_n379), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n751), .A2(new_n752), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(KEYINPUT113), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT53), .ZN(new_n776));
  INV_X1    g575(.A(G106gat), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n740), .A2(new_n379), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n775), .B(new_n776), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n774), .A2(KEYINPUT113), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n741), .A2(new_n671), .A3(new_n743), .ZN(new_n781));
  AOI22_X1  g580(.A1(new_n781), .A2(G106gat), .B1(new_n763), .B2(new_n773), .ZN(new_n782));
  OAI22_X1  g581(.A1(new_n779), .A2(new_n780), .B1(new_n782), .B2(new_n776), .ZN(G1339gat));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n601), .B1(new_n614), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n594), .A2(new_n597), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n784), .B1(new_n593), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n594), .B1(new_n609), .B2(new_n558), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n787), .B1(new_n788), .B2(new_n613), .ZN(new_n789));
  AND4_X1   g588(.A1(KEYINPUT114), .A2(new_n785), .A3(KEYINPUT55), .A4(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT55), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n791), .B1(new_n598), .B2(new_n787), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT114), .B1(new_n792), .B2(new_n785), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n596), .A2(new_n784), .A3(new_n597), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n593), .A2(new_n786), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(KEYINPUT54), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n795), .B(new_n612), .C1(new_n797), .C2(new_n614), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n791), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n517), .A2(new_n518), .A3(new_n515), .ZN(new_n800));
  INV_X1    g599(.A(new_n499), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n498), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n501), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT115), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n802), .A2(KEYINPUT115), .A3(new_n501), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n505), .A2(new_n506), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n800), .B1(new_n808), .B2(new_n513), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n614), .A2(new_n615), .A3(new_n612), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n644), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n799), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n794), .A2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n617), .A2(new_n809), .A3(new_n618), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n799), .A2(new_n522), .A3(new_n610), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n816), .B1(new_n794), .B2(new_n817), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n818), .A2(new_n644), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n557), .B1(new_n815), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n646), .A2(new_n523), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n671), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n653), .A2(new_n668), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT117), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n272), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n822), .A2(KEYINPUT117), .A3(new_n823), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(G113gat), .B1(new_n828), .B2(new_n522), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n824), .A2(new_n272), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n522), .A2(G113gat), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(G1340gat));
  AOI21_X1  g631(.A(G120gat), .B1(new_n828), .B2(new_n619), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n619), .A2(G120gat), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n833), .B1(new_n830), .B2(new_n834), .ZN(G1341gat));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n828), .A2(new_n836), .A3(new_n680), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n837), .A2(new_n275), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n828), .A2(new_n680), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(KEYINPUT118), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n557), .A2(new_n275), .ZN(new_n841));
  AOI22_X1  g640(.A1(new_n838), .A2(new_n840), .B1(new_n830), .B2(new_n841), .ZN(G1342gat));
  NAND3_X1  g641(.A1(new_n828), .A2(new_n276), .A3(new_n645), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n843), .A2(KEYINPUT56), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n656), .A2(new_n645), .ZN(new_n845));
  OAI21_X1  g644(.A(G134gat), .B1(new_n824), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n843), .A2(KEYINPUT56), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n844), .A2(new_n846), .A3(new_n847), .ZN(G1343gat));
  NAND3_X1  g647(.A1(new_n666), .A2(new_n656), .A3(new_n652), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n820), .A2(new_n821), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n671), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n850), .A2(KEYINPUT57), .A3(new_n671), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n849), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n522), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(G141gat), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT120), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n851), .A2(new_n849), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n523), .A2(G141gat), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n861), .B(KEYINPUT119), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n857), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n859), .A2(new_n864), .A3(KEYINPUT58), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT58), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n857), .B(new_n863), .C1(new_n858), .C2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(G1344gat));
  OR4_X1    g667(.A1(G148gat), .A2(new_n851), .A3(new_n707), .A4(new_n849), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n849), .A2(new_n707), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n813), .B1(new_n818), .B2(new_n644), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n821), .B1(new_n872), .B2(new_n680), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n379), .B1(new_n873), .B2(KEYINPUT121), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT121), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n821), .B(new_n875), .C1(new_n872), .C2(new_n680), .ZN(new_n876));
  AOI21_X1  g675(.A(KEYINPUT57), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n854), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AOI211_X1 g678(.A(KEYINPUT122), .B(KEYINPUT57), .C1(new_n874), .C2(new_n876), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n871), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n870), .B1(new_n881), .B2(G148gat), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n870), .A2(G148gat), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n883), .B1(new_n855), .B2(new_n619), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n869), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT123), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI211_X1 g686(.A(KEYINPUT123), .B(new_n869), .C1(new_n882), .C2(new_n884), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(G1345gat));
  AOI21_X1  g688(.A(G155gat), .B1(new_n860), .B2(new_n680), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n680), .A2(G155gat), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n890), .B1(new_n855), .B2(new_n891), .ZN(G1346gat));
  INV_X1    g691(.A(G162gat), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n860), .A2(new_n893), .A3(new_n645), .ZN(new_n894));
  XOR2_X1   g693(.A(new_n894), .B(KEYINPUT124), .Z(new_n895));
  AND2_X1   g694(.A1(new_n855), .A2(new_n645), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n893), .B2(new_n896), .ZN(G1347gat));
  NAND2_X1  g696(.A1(new_n653), .A2(new_n272), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n898), .A2(new_n668), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n822), .A2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(G169gat), .B1(new_n901), .B2(new_n523), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n652), .B1(new_n820), .B2(new_n821), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n903), .A2(new_n272), .A3(new_n448), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(new_n522), .A3(new_n227), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n902), .A2(new_n905), .ZN(G1348gat));
  AOI21_X1  g705(.A(G176gat), .B1(new_n904), .B2(new_n619), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n707), .A2(new_n228), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n900), .B2(new_n908), .ZN(G1349gat));
  AOI21_X1  g708(.A(new_n223), .B1(new_n900), .B2(new_n680), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n680), .A2(new_n235), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n910), .B1(new_n904), .B2(new_n911), .ZN(new_n912));
  XOR2_X1   g711(.A(new_n912), .B(KEYINPUT60), .Z(G1350gat));
  AOI21_X1  g712(.A(new_n224), .B1(new_n900), .B2(new_n645), .ZN(new_n914));
  XOR2_X1   g713(.A(new_n914), .B(KEYINPUT61), .Z(new_n915));
  NAND3_X1  g714(.A1(new_n904), .A2(new_n224), .A3(new_n645), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(G1351gat));
  XNOR2_X1  g716(.A(KEYINPUT125), .B(G197gat), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n879), .A2(new_n880), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n898), .A2(new_n665), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(KEYINPUT126), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n918), .B1(new_n922), .B2(new_n522), .ZN(new_n923));
  AND4_X1   g722(.A1(new_n272), .A2(new_n903), .A3(new_n671), .A4(new_n666), .ZN(new_n924));
  AND3_X1   g723(.A1(new_n924), .A2(new_n522), .A3(new_n918), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n923), .A2(new_n925), .ZN(G1352gat));
  INV_X1    g725(.A(G204gat), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n927), .B1(new_n922), .B2(new_n619), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n924), .A2(new_n927), .A3(new_n619), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT62), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n928), .A2(new_n930), .ZN(G1353gat));
  NAND3_X1  g730(.A1(new_n924), .A2(new_n204), .A3(new_n680), .ZN(new_n932));
  OR2_X1    g731(.A1(new_n879), .A2(new_n880), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n898), .A2(new_n665), .A3(new_n557), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n204), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n935), .A2(KEYINPUT63), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n935), .A2(KEYINPUT63), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n932), .B1(new_n936), .B2(new_n937), .ZN(G1354gat));
  INV_X1    g737(.A(KEYINPUT127), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n645), .B1(new_n922), .B2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(new_n921), .ZN(new_n941));
  OAI211_X1 g740(.A(new_n941), .B(new_n939), .C1(new_n880), .C2(new_n879), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  OAI21_X1  g742(.A(G218gat), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n924), .A2(new_n205), .A3(new_n645), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1355gat));
endmodule


