//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 0 1 1 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 0 1 0 1 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n873, new_n874, new_n876, new_n877, new_n878,
    new_n879, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n985, new_n986;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(G169gat), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n205), .A2(G197gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(G197gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT81), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT81), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n206), .A2(new_n210), .A3(new_n207), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(KEYINPUT12), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT12), .ZN(new_n213));
  INV_X1    g012(.A(new_n211), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n210), .B1(new_n206), .B2(new_n207), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(G229gat), .A2(G233gat), .ZN(new_n217));
  XOR2_X1   g016(.A(new_n217), .B(KEYINPUT13), .Z(new_n218));
  XNOR2_X1  g017(.A(G15gat), .B(G22gat), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n219), .A2(KEYINPUT85), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n219), .A2(KEYINPUT85), .ZN(new_n221));
  OR3_X1    g020(.A1(new_n220), .A2(new_n221), .A3(G1gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT86), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n224));
  OAI22_X1  g023(.A1(new_n220), .A2(new_n221), .B1(new_n224), .B2(G1gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n222), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G8gat), .ZN(new_n227));
  INV_X1    g026(.A(G8gat), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n222), .A2(new_n223), .A3(new_n228), .A4(new_n225), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(G29gat), .A2(G36gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT14), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT83), .B(G36gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G29gat), .ZN(new_n235));
  INV_X1    g034(.A(G43gat), .ZN(new_n236));
  INV_X1    g035(.A(G50gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT15), .ZN(new_n239));
  NAND2_X1  g038(.A1(G43gat), .A2(G50gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n233), .A2(new_n235), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n238), .A2(new_n240), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT82), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n238), .A2(KEYINPUT82), .A3(new_n240), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(KEYINPUT15), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n242), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n239), .B1(new_n243), .B2(new_n244), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n249), .A2(new_n233), .A3(new_n246), .A4(new_n235), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n230), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n248), .A2(new_n250), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n252), .B1(new_n227), .B2(new_n229), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n218), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n230), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT17), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n256), .B1(new_n252), .B2(KEYINPUT84), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT84), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n248), .A2(new_n258), .A3(KEYINPUT17), .A4(new_n250), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n255), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n253), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT87), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n263), .A2(KEYINPUT18), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n261), .A2(new_n217), .A3(new_n262), .A4(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n254), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n253), .B1(new_n255), .B2(new_n260), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n265), .B1(new_n268), .B2(new_n217), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n212), .B(new_n216), .C1(new_n267), .C2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n269), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n216), .A2(new_n212), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n271), .A2(new_n272), .A3(new_n254), .A4(new_n266), .ZN(new_n273));
  AND2_X1   g072(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  AND2_X1   g073(.A1(G71gat), .A2(G78gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(G71gat), .A2(G78gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G57gat), .B(G64gat), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G57gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(G64gat), .ZN(new_n282));
  INV_X1    g081(.A(G64gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(G57gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G71gat), .B(G78gat), .ZN(new_n286));
  INV_X1    g085(.A(new_n279), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  AND3_X1   g087(.A1(new_n280), .A2(new_n288), .A3(KEYINPUT89), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT89), .B1(new_n280), .B2(new_n288), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT21), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n255), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G183gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n288), .ZN(new_n296));
  XOR2_X1   g095(.A(KEYINPUT88), .B(KEYINPUT21), .Z(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n299));
  XOR2_X1   g098(.A(new_n298), .B(new_n299), .Z(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n295), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n295), .A2(new_n301), .ZN(new_n303));
  XNOR2_X1  g102(.A(G127gat), .B(G155gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(G231gat), .A2(G233gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n304), .B(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G211gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n306), .B(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  OR3_X1    g108(.A1(new_n302), .A2(new_n303), .A3(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n309), .B1(new_n302), .B2(new_n303), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G134gat), .B(G162gat), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n314));
  XOR2_X1   g113(.A(new_n313), .B(new_n314), .Z(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(G85gat), .A2(G92gat), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT90), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(KEYINPUT90), .A2(G85gat), .A3(G92gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n319), .A2(KEYINPUT7), .A3(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(G99gat), .B(G106gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT7), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n317), .A2(new_n318), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G99gat), .A2(G106gat), .ZN(new_n325));
  INV_X1    g124(.A(G85gat), .ZN(new_n326));
  INV_X1    g125(.A(G92gat), .ZN(new_n327));
  AOI22_X1  g126(.A1(KEYINPUT8), .A2(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n321), .A2(new_n322), .A3(new_n324), .A4(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n322), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n319), .A2(KEYINPUT7), .A3(new_n320), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n325), .A2(KEYINPUT8), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n326), .A2(new_n327), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n324), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n330), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n248), .A2(new_n250), .A3(new_n329), .A4(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n337));
  AND3_X1   g136(.A1(new_n336), .A2(KEYINPUT91), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT91), .B1(new_n336), .B2(new_n337), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n335), .A2(new_n329), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n341), .B1(new_n257), .B2(new_n259), .ZN(new_n342));
  OAI21_X1  g141(.A(G190gat), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n342), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n336), .A2(new_n337), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT91), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n336), .A2(KEYINPUT91), .A3(new_n337), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(G190gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n344), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  AND3_X1   g150(.A1(new_n343), .A2(new_n351), .A3(G218gat), .ZN(new_n352));
  AOI21_X1  g151(.A(G218gat), .B1(new_n343), .B2(new_n351), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n316), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT93), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI211_X1 g155(.A(KEYINPUT93), .B(new_n316), .C1(new_n352), .C2(new_n353), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n343), .A2(new_n351), .ZN(new_n358));
  INV_X1    g157(.A(G218gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n343), .A2(new_n351), .A3(G218gat), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n360), .A2(new_n315), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT92), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n360), .A2(KEYINPUT92), .A3(new_n315), .A4(new_n361), .ZN(new_n365));
  AOI22_X1  g164(.A1(new_n356), .A2(new_n357), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT94), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT89), .ZN(new_n368));
  AND3_X1   g167(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n286), .B1(new_n287), .B2(new_n285), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n280), .A2(new_n288), .A3(KEYINPUT89), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n371), .A2(KEYINPUT10), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n335), .A2(new_n329), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n367), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n291), .A2(KEYINPUT94), .A3(KEYINPUT10), .A4(new_n341), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n296), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n335), .A2(new_n280), .A3(new_n288), .A4(new_n329), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n375), .A2(new_n376), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(G230gat), .A2(G233gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n377), .A2(new_n379), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n383), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(G120gat), .B(G148gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n386), .B(G176gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(G204gat), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n385), .A2(new_n388), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n312), .A2(new_n366), .A3(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(G78gat), .B(G106gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n395), .B(G22gat), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  AND2_X1   g196(.A1(G228gat), .A2(G233gat), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT29), .ZN(new_n399));
  NAND2_X1  g198(.A1(G211gat), .A2(G218gat), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT22), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT72), .B(G197gat), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n403), .A2(G204gat), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(G204gat), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n402), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n307), .A2(new_n359), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n400), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT73), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n407), .A2(KEYINPUT73), .A3(new_n400), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n406), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n403), .B(G204gat), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n412), .B1(new_n415), .B2(new_n402), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n399), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT3), .ZN(new_n418));
  XNOR2_X1  g217(.A(G141gat), .B(G148gat), .ZN(new_n419));
  OR2_X1    g218(.A1(new_n419), .A2(KEYINPUT77), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(KEYINPUT77), .ZN(new_n421));
  NAND2_X1  g220(.A1(G155gat), .A2(G162gat), .ZN(new_n422));
  INV_X1    g221(.A(G155gat), .ZN(new_n423));
  INV_X1    g222(.A(G162gat), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n422), .B1(new_n425), .B2(KEYINPUT2), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n420), .A2(new_n421), .A3(new_n426), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n425), .A2(new_n422), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n428), .B1(KEYINPUT2), .B2(new_n419), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT76), .ZN(new_n430));
  XOR2_X1   g229(.A(G141gat), .B(G148gat), .Z(new_n431));
  INV_X1    g230(.A(KEYINPUT2), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT76), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n433), .A2(new_n434), .A3(new_n428), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n430), .A2(new_n435), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n417), .A2(new_n418), .B1(new_n427), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n406), .A2(new_n413), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n415), .A2(new_n412), .A3(new_n402), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n429), .A2(KEYINPUT76), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n434), .B1(new_n433), .B2(new_n428), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n418), .B(new_n427), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n440), .B1(new_n399), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n398), .B1(new_n437), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n443), .A2(new_n399), .ZN(new_n446));
  INV_X1    g245(.A(new_n440), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n398), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT80), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT29), .B1(new_n416), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n438), .A2(KEYINPUT80), .A3(new_n439), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT3), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT78), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n453), .B(new_n427), .C1(new_n441), .C2(new_n442), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n453), .B1(new_n436), .B2(new_n427), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n448), .B1(new_n452), .B2(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(G50gat), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n445), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n461), .B1(new_n445), .B2(new_n458), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n397), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n445), .A2(new_n458), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(new_n460), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n445), .A2(new_n458), .A3(new_n461), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(new_n396), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(KEYINPUT27), .B(G183gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n350), .ZN(new_n471));
  AOI22_X1  g270(.A1(new_n471), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(G169gat), .A2(G176gat), .ZN(new_n473));
  OAI21_X1  g272(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n474));
  NOR4_X1   g273(.A1(KEYINPUT66), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT66), .ZN(new_n476));
  NOR2_X1   g275(.A1(G169gat), .A2(G176gat), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT26), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n473), .B(new_n474), .C1(new_n475), .C2(new_n479), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n472), .B(new_n480), .C1(KEYINPUT28), .C2(new_n471), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n482), .B1(new_n294), .B2(new_n350), .ZN(new_n483));
  NAND3_X1  g282(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT65), .ZN(new_n485));
  OR2_X1    g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n485), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n483), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n477), .A2(KEYINPUT23), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT23), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n490), .B1(G169gat), .B2(G176gat), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n489), .A2(new_n473), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT25), .B1(new_n488), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT64), .ZN(new_n494));
  OR2_X1    g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n492), .A2(new_n494), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT25), .B1(new_n483), .B2(new_n484), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n481), .A2(new_n493), .A3(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(G113gat), .B(G120gat), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT67), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT1), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n502), .B1(new_n501), .B2(new_n500), .ZN(new_n503));
  XOR2_X1   g302(.A(G127gat), .B(G134gat), .Z(new_n504));
  XOR2_X1   g303(.A(KEYINPUT68), .B(KEYINPUT1), .Z(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n500), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n503), .A2(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n499), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(G227gat), .ZN(new_n509));
  INV_X1    g308(.A(G233gat), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n503), .A2(new_n504), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n506), .A2(new_n505), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n514), .A2(new_n481), .A3(new_n493), .A4(new_n498), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n508), .A2(new_n511), .A3(new_n515), .ZN(new_n516));
  XOR2_X1   g315(.A(G71gat), .B(G99gat), .Z(new_n517));
  XNOR2_X1  g316(.A(G15gat), .B(G43gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT69), .B(KEYINPUT33), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n516), .A2(KEYINPUT32), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT70), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT70), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n516), .A2(new_n525), .A3(KEYINPUT32), .A4(new_n522), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n516), .A2(KEYINPUT32), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n516), .A2(new_n520), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(new_n529), .A3(new_n519), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n511), .B1(new_n508), .B2(new_n515), .ZN(new_n532));
  OR2_X1    g331(.A1(new_n532), .A2(KEYINPUT34), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(KEYINPUT34), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n527), .A2(new_n535), .A3(new_n530), .ZN(new_n538));
  AND3_X1   g337(.A1(new_n469), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(G226gat), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n540), .A2(new_n510), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n541), .A2(KEYINPUT29), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT74), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n499), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n481), .A2(new_n493), .A3(KEYINPUT74), .A4(new_n498), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n543), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NOR3_X1   g346(.A1(new_n499), .A2(new_n540), .A3(new_n510), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n440), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G8gat), .B(G36gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(G92gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(KEYINPUT75), .B(G64gat), .ZN(new_n552));
  XOR2_X1   g351(.A(new_n551), .B(new_n552), .Z(new_n553));
  NAND3_X1  g352(.A1(new_n545), .A2(new_n546), .A3(new_n541), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n499), .A2(new_n542), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n554), .A2(new_n447), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n549), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT30), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n553), .ZN(new_n560));
  INV_X1    g359(.A(new_n549), .ZN(new_n561));
  INV_X1    g360(.A(new_n556), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n549), .A2(KEYINPUT30), .A3(new_n553), .A4(new_n556), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n559), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n427), .B1(new_n441), .B2(new_n442), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT78), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n567), .A2(KEYINPUT4), .A3(new_n507), .A4(new_n454), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(KEYINPUT3), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n569), .A2(new_n443), .A3(new_n514), .ZN(new_n570));
  NAND2_X1  g369(.A1(G225gat), .A2(G233gat), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n507), .A2(new_n427), .A3(new_n436), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT4), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n568), .A2(new_n570), .A3(new_n571), .A4(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT5), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n514), .A2(new_n566), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(new_n572), .ZN(new_n578));
  INV_X1    g377(.A(new_n571), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n576), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n567), .A2(new_n573), .A3(new_n507), .A4(new_n454), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n572), .A2(KEYINPUT4), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n507), .B1(new_n566), .B2(KEYINPUT3), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n579), .B1(new_n585), .B2(new_n443), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n584), .A2(new_n576), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G1gat), .B(G29gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT0), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(G57gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(new_n326), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n588), .A2(KEYINPUT6), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n588), .A2(new_n593), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT6), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n581), .A2(new_n592), .A3(new_n587), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n565), .B1(new_n594), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(KEYINPUT35), .B1(new_n539), .B2(new_n599), .ZN(new_n600));
  AND3_X1   g399(.A1(new_n559), .A2(new_n563), .A3(new_n564), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n533), .A2(KEYINPUT71), .A3(new_n534), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n531), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n527), .A2(new_n602), .A3(new_n530), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n601), .A2(new_n469), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n598), .A2(new_n594), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(KEYINPUT35), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n600), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n607), .A2(new_n601), .ZN(new_n611));
  INV_X1    g410(.A(new_n469), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT36), .ZN(new_n613));
  INV_X1    g412(.A(new_n538), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n535), .B1(new_n527), .B2(new_n530), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n604), .A2(KEYINPUT36), .A3(new_n605), .ZN(new_n617));
  AOI22_X1  g416(.A1(new_n611), .A2(new_n612), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n577), .A2(new_n572), .A3(new_n571), .ZN(new_n619));
  AOI22_X1  g418(.A1(new_n582), .A2(new_n583), .B1(new_n443), .B2(new_n585), .ZN(new_n620));
  OAI211_X1 g419(.A(KEYINPUT39), .B(new_n619), .C1(new_n620), .C2(new_n571), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n584), .A2(new_n570), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT39), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n622), .A2(new_n623), .A3(new_n579), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n621), .A2(new_n624), .A3(new_n592), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT40), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n621), .A2(new_n624), .A3(KEYINPUT40), .A4(new_n592), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n565), .A2(new_n595), .A3(new_n627), .A4(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(KEYINPUT37), .B1(new_n561), .B2(new_n562), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT37), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n549), .A2(new_n631), .A3(new_n556), .ZN(new_n632));
  AND2_X1   g431(.A1(new_n632), .A2(KEYINPUT38), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n447), .B1(new_n547), .B2(new_n548), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n554), .A2(new_n440), .A3(new_n555), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n634), .A2(KEYINPUT37), .A3(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n632), .A2(new_n636), .A3(new_n560), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT38), .ZN(new_n638));
  AOI22_X1  g437(.A1(new_n630), .A2(new_n633), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n638), .B1(new_n561), .B2(new_n562), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(new_n553), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n598), .A2(new_n641), .A3(new_n594), .ZN(new_n642));
  OAI211_X1 g441(.A(new_n629), .B(new_n469), .C1(new_n639), .C2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n618), .A2(new_n643), .ZN(new_n644));
  AOI211_X1 g443(.A(new_n274), .B(new_n394), .C1(new_n610), .C2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n607), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g447(.A1(new_n645), .A2(new_n565), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n649), .A2(new_n228), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT42), .ZN(new_n651));
  XOR2_X1   g450(.A(KEYINPUT16), .B(G8gat), .Z(new_n652));
  NAND2_X1  g451(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n650), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n654), .B1(new_n651), .B2(new_n653), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT95), .ZN(G1325gat));
  NAND2_X1  g455(.A1(new_n616), .A2(new_n617), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n645), .A2(new_n658), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n614), .A2(G15gat), .A3(new_n615), .ZN(new_n660));
  AOI22_X1  g459(.A1(new_n659), .A2(G15gat), .B1(new_n645), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT96), .ZN(G1326gat));
  NAND2_X1  g461(.A1(new_n645), .A2(new_n612), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT43), .B(G22gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(G1327gat));
  AOI21_X1  g464(.A(new_n366), .B1(new_n610), .B2(new_n644), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n312), .A2(new_n274), .A3(new_n392), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(G29gat), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n668), .A2(new_n669), .A3(new_n646), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT97), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT45), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n356), .A2(new_n357), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n364), .A2(new_n365), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n618), .A2(new_n643), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT35), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n469), .A2(new_n537), .A3(new_n538), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n678), .B1(new_n611), .B2(new_n679), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n604), .A2(new_n605), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n678), .B1(new_n598), .B2(new_n594), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n681), .A2(new_n682), .A3(new_n601), .A4(new_n469), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n676), .B1(new_n677), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n685), .A2(KEYINPUT98), .A3(KEYINPUT44), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT98), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n687), .B1(new_n666), .B2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT99), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n690), .B1(new_n600), .B2(new_n609), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n680), .A2(KEYINPUT99), .A3(new_n683), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(new_n644), .A3(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n693), .A2(new_n688), .A3(new_n676), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n686), .A2(new_n689), .A3(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n695), .A2(new_n646), .A3(new_n667), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT100), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n669), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n698), .B1(new_n697), .B2(new_n696), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n671), .A2(new_n672), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n673), .A2(new_n699), .A3(new_n700), .ZN(G1328gat));
  NAND2_X1  g500(.A1(new_n695), .A2(new_n667), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n234), .B1(new_n702), .B2(new_n601), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n234), .B1(KEYINPUT101), .B2(KEYINPUT46), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n668), .A2(new_n565), .A3(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(KEYINPUT101), .A2(KEYINPUT46), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n703), .A2(new_n707), .ZN(G1329gat));
  OAI21_X1  g507(.A(G43gat), .B1(new_n702), .B2(new_n657), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n614), .A2(new_n615), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n668), .A2(new_n236), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n712), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g512(.A(G50gat), .B1(new_n702), .B2(new_n469), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n668), .A2(new_n237), .A3(new_n612), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT103), .ZN(new_n716));
  OR2_X1    g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n716), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n714), .A2(KEYINPUT48), .A3(new_n717), .A4(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(KEYINPUT48), .B1(new_n714), .B2(new_n715), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT102), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI211_X1 g521(.A(KEYINPUT102), .B(KEYINPUT48), .C1(new_n714), .C2(new_n715), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n719), .B1(new_n722), .B2(new_n723), .ZN(G1331gat));
  INV_X1    g523(.A(new_n312), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n270), .A2(new_n273), .ZN(new_n726));
  NOR4_X1   g525(.A1(new_n725), .A2(new_n726), .A3(new_n676), .A4(new_n393), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n693), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n728), .A2(new_n607), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(new_n281), .ZN(G1332gat));
  INV_X1    g529(.A(KEYINPUT104), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n693), .A2(KEYINPUT104), .A3(new_n727), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n565), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n735), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n736));
  XOR2_X1   g535(.A(KEYINPUT49), .B(G64gat), .Z(new_n737));
  OAI21_X1  g536(.A(new_n736), .B1(new_n735), .B2(new_n737), .ZN(G1333gat));
  NAND3_X1  g537(.A1(new_n732), .A2(new_n658), .A3(new_n733), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(G71gat), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT105), .ZN(new_n741));
  OR4_X1    g540(.A1(G71gat), .A2(new_n728), .A3(new_n615), .A4(new_n614), .ZN(new_n742));
  AND3_X1   g541(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n741), .B1(new_n740), .B2(new_n742), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT50), .ZN(new_n745));
  OR3_X1    g544(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n743), .B2(new_n744), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(G1334gat));
  NAND2_X1  g547(.A1(new_n734), .A2(new_n612), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g549(.A1(new_n312), .A2(new_n726), .A3(new_n393), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n695), .A2(new_n646), .A3(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT106), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n326), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n753), .B2(new_n752), .ZN(new_n755));
  AOI22_X1  g554(.A1(new_n684), .A2(new_n690), .B1(new_n643), .B2(new_n618), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n366), .B1(new_n756), .B2(new_n692), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT107), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n312), .A2(new_n726), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n757), .A2(new_n758), .A3(KEYINPUT51), .A4(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n693), .A2(KEYINPUT51), .A3(new_n676), .A4(new_n759), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT107), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n693), .A2(new_n676), .A3(new_n759), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n763), .B1(KEYINPUT51), .B2(new_n765), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n766), .A2(new_n326), .A3(new_n646), .A4(new_n392), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n755), .A2(new_n767), .ZN(G1336gat));
  XOR2_X1   g567(.A(KEYINPUT108), .B(KEYINPUT51), .Z(new_n769));
  NAND2_X1  g568(.A1(new_n764), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT109), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n764), .A2(KEYINPUT109), .A3(new_n769), .ZN(new_n773));
  AOI22_X1  g572(.A1(new_n772), .A2(new_n773), .B1(new_n762), .B2(new_n760), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n601), .A2(G92gat), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n392), .ZN(new_n776));
  OAI21_X1  g575(.A(KEYINPUT110), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n778));
  INV_X1    g577(.A(new_n776), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n764), .A2(KEYINPUT109), .A3(new_n769), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT109), .B1(new_n764), .B2(new_n769), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n761), .B(new_n758), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n778), .B(new_n779), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n695), .A2(new_n751), .ZN(new_n785));
  OAI21_X1  g584(.A(G92gat), .B1(new_n785), .B2(new_n601), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n777), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT52), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n766), .A2(new_n392), .A3(new_n775), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT111), .ZN(new_n790));
  OR2_X1    g589(.A1(new_n790), .A2(KEYINPUT52), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(KEYINPUT52), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n789), .A2(new_n786), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n788), .A2(new_n793), .ZN(G1337gat));
  INV_X1    g593(.A(G99gat), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n785), .A2(new_n795), .A3(new_n657), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n766), .A2(new_n710), .A3(new_n392), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n796), .B1(new_n797), .B2(new_n795), .ZN(G1338gat));
  NOR3_X1   g597(.A1(new_n393), .A2(new_n469), .A3(G106gat), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT53), .B1(new_n766), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n695), .A2(new_n612), .A3(new_n751), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n802), .A2(KEYINPUT114), .ZN(new_n803));
  XNOR2_X1  g602(.A(KEYINPUT112), .B(G106gat), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n804), .B1(new_n802), .B2(KEYINPUT114), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n800), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT113), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n799), .B1(new_n782), .B2(new_n783), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n801), .A2(new_n804), .ZN(new_n810));
  AOI211_X1 g609(.A(new_n807), .B(new_n808), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n799), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n810), .B1(new_n774), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT113), .B1(new_n813), .B2(KEYINPUT53), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n806), .B1(new_n811), .B2(new_n814), .ZN(G1339gat));
  INV_X1    g614(.A(new_n382), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n375), .A2(new_n376), .A3(new_n380), .A4(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n383), .A2(KEYINPUT54), .A3(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n821), .B1(new_n381), .B2(new_n382), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n822), .A2(KEYINPUT115), .A3(new_n817), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g623(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n381), .A2(new_n382), .A3(new_n825), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n826), .A2(KEYINPUT55), .A3(new_n388), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n389), .B1(new_n824), .B2(new_n827), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n826), .A2(new_n388), .ZN(new_n829));
  AND4_X1   g628(.A1(KEYINPUT115), .A2(new_n383), .A3(KEYINPUT54), .A4(new_n817), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT115), .B1(new_n822), .B2(new_n817), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT55), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n828), .A2(new_n834), .A3(KEYINPUT117), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT117), .B1(new_n828), .B2(new_n834), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n726), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT118), .B1(new_n268), .B2(new_n217), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n251), .A2(new_n253), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n838), .B1(new_n839), .B2(new_n218), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n268), .A2(KEYINPUT118), .A3(new_n217), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n208), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n273), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n392), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n676), .B1(new_n837), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT117), .ZN(new_n847));
  AOI21_X1  g646(.A(KEYINPUT55), .B1(new_n824), .B2(new_n829), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n827), .B1(new_n830), .B2(new_n831), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n390), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n847), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n828), .A2(new_n834), .A3(KEYINPUT117), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AND3_X1   g652(.A1(new_n676), .A2(new_n853), .A3(new_n844), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n725), .B1(new_n846), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n394), .A2(new_n726), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n607), .A2(new_n565), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n858), .A2(new_n539), .A3(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(G113gat), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n860), .A2(new_n861), .A3(new_n274), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n607), .B1(new_n855), .B2(new_n857), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n681), .A2(new_n469), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n863), .A2(new_n601), .A3(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n726), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n862), .B1(new_n867), .B2(new_n861), .ZN(G1340gat));
  INV_X1    g667(.A(G120gat), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n860), .A2(new_n869), .A3(new_n393), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n866), .A2(new_n392), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n870), .B1(new_n871), .B2(new_n869), .ZN(G1341gat));
  OAI21_X1  g671(.A(G127gat), .B1(new_n860), .B2(new_n725), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n725), .A2(G127gat), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n873), .B1(new_n865), .B2(new_n874), .ZN(G1342gat));
  INV_X1    g674(.A(G134gat), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n866), .A2(new_n876), .A3(new_n676), .ZN(new_n877));
  OR2_X1    g676(.A1(new_n860), .A2(new_n366), .ZN(new_n878));
  AOI22_X1  g677(.A1(new_n877), .A2(KEYINPUT56), .B1(G134gat), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n879), .B1(KEYINPUT56), .B2(new_n877), .ZN(G1343gat));
  NAND2_X1  g679(.A1(new_n828), .A2(new_n834), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n274), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n843), .A2(new_n393), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n366), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n676), .A2(new_n853), .A3(new_n844), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n312), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n612), .B1(new_n886), .B2(new_n856), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(KEYINPUT57), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n274), .B1(new_n851), .B2(new_n852), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n366), .B1(new_n890), .B2(new_n883), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n312), .B1(new_n891), .B2(new_n885), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n889), .B(new_n612), .C1(new_n892), .C2(new_n856), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n657), .A2(new_n859), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n888), .A2(new_n893), .A3(new_n726), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(G141gat), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n658), .A2(new_n565), .A3(new_n469), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n274), .A2(G141gat), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n863), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(KEYINPUT119), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT119), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n896), .A2(new_n899), .A3(new_n902), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n901), .A2(KEYINPUT58), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT58), .B1(new_n901), .B2(new_n903), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n904), .A2(new_n905), .ZN(G1344gat));
  INV_X1    g705(.A(G148gat), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n863), .A2(new_n907), .A3(new_n392), .A4(new_n897), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT59), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n889), .B1(new_n858), .B2(new_n612), .ZN(new_n910));
  OR3_X1    g709(.A1(new_n366), .A2(KEYINPUT120), .A3(new_n881), .ZN(new_n911));
  OAI21_X1  g710(.A(KEYINPUT120), .B1(new_n366), .B2(new_n881), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n911), .A2(new_n844), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n312), .B1(new_n913), .B2(new_n884), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n914), .A2(new_n856), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n469), .A2(KEYINPUT57), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n910), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n917), .A2(new_n392), .A3(new_n894), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n909), .B1(new_n918), .B2(G148gat), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n888), .A2(new_n893), .A3(new_n894), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n920), .A2(new_n393), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n921), .A2(KEYINPUT59), .A3(new_n907), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n908), .B1(new_n919), .B2(new_n922), .ZN(G1345gat));
  OAI21_X1  g722(.A(G155gat), .B1(new_n920), .B2(new_n725), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n863), .A2(new_n423), .A3(new_n312), .A4(new_n897), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1346gat));
  OAI21_X1  g725(.A(G162gat), .B1(new_n920), .B2(new_n366), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n863), .A2(new_n424), .A3(new_n676), .A4(new_n897), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(G1347gat));
  NAND2_X1  g728(.A1(new_n864), .A2(new_n565), .ZN(new_n930));
  XOR2_X1   g729(.A(new_n930), .B(KEYINPUT121), .Z(new_n931));
  NAND3_X1  g730(.A1(new_n858), .A2(new_n607), .A3(new_n931), .ZN(new_n932));
  OR3_X1    g731(.A1(new_n932), .A2(G169gat), .A3(new_n274), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n646), .A2(new_n601), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n539), .B(new_n934), .C1(new_n892), .C2(new_n856), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT122), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n858), .A2(KEYINPUT122), .A3(new_n539), .A4(new_n934), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g738(.A(G169gat), .B1(new_n939), .B2(new_n274), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT123), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n933), .B1(new_n942), .B2(new_n943), .ZN(G1348gat));
  OAI21_X1  g743(.A(G176gat), .B1(new_n939), .B2(new_n393), .ZN(new_n945));
  OR2_X1    g744(.A1(new_n393), .A2(G176gat), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n945), .B1(new_n932), .B2(new_n946), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT124), .ZN(G1349gat));
  NAND2_X1  g747(.A1(new_n312), .A2(new_n470), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n932), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n937), .A2(new_n938), .A3(new_n312), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n950), .B1(new_n951), .B2(G183gat), .ZN(new_n952));
  AOI211_X1 g751(.A(KEYINPUT125), .B(KEYINPUT60), .C1(new_n952), .C2(KEYINPUT126), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(KEYINPUT126), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT125), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT60), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n957), .B1(new_n952), .B2(KEYINPUT125), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n953), .B1(new_n956), .B2(new_n958), .ZN(G1350gat));
  OAI21_X1  g758(.A(G190gat), .B1(new_n939), .B2(new_n366), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n960), .A2(KEYINPUT61), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n960), .A2(KEYINPUT61), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n676), .A2(new_n350), .ZN(new_n963));
  OAI22_X1  g762(.A1(new_n961), .A2(new_n962), .B1(new_n932), .B2(new_n963), .ZN(G1351gat));
  NAND2_X1  g763(.A1(new_n934), .A2(new_n657), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n917), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g766(.A(G197gat), .B1(new_n967), .B2(new_n274), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n658), .A2(new_n601), .A3(new_n469), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n858), .A2(new_n607), .A3(new_n969), .ZN(new_n970));
  XOR2_X1   g769(.A(new_n970), .B(KEYINPUT127), .Z(new_n971));
  INV_X1    g770(.A(G197gat), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n971), .A2(new_n972), .A3(new_n726), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n968), .A2(new_n973), .ZN(G1352gat));
  NAND3_X1  g773(.A1(new_n917), .A2(new_n392), .A3(new_n966), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(G204gat), .ZN(new_n976));
  NOR3_X1   g775(.A1(new_n970), .A2(G204gat), .A3(new_n393), .ZN(new_n977));
  XNOR2_X1  g776(.A(new_n977), .B(KEYINPUT62), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n976), .A2(new_n978), .ZN(G1353gat));
  NAND3_X1  g778(.A1(new_n971), .A2(new_n307), .A3(new_n312), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n917), .A2(new_n312), .A3(new_n966), .ZN(new_n981));
  AND3_X1   g780(.A1(new_n981), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n982));
  AOI21_X1  g781(.A(KEYINPUT63), .B1(new_n981), .B2(G211gat), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(G1354gat));
  OAI21_X1  g783(.A(G218gat), .B1(new_n967), .B2(new_n366), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n971), .A2(new_n359), .A3(new_n676), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(G1355gat));
endmodule


