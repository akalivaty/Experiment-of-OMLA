//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 0 0 1 0 1 1 0 0 0 0 1 0 0 0 1 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n785,
    new_n787, new_n788, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n868, new_n869, new_n870,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT3), .ZN(new_n203));
  XNOR2_X1  g002(.A(G211gat), .B(G218gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT73), .ZN(new_n205));
  INV_X1    g004(.A(G197gat), .ZN(new_n206));
  INV_X1    g005(.A(G204gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G197gat), .A2(G204gat), .ZN(new_n209));
  AND2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n211));
  OR2_X1    g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n205), .B(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n203), .B1(new_n213), .B2(KEYINPUT29), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT76), .ZN(new_n215));
  INV_X1    g014(.A(G148gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n215), .B1(new_n216), .B2(G141gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT77), .ZN(new_n218));
  INV_X1    g017(.A(G141gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n218), .B1(new_n219), .B2(G148gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(KEYINPUT76), .A3(G148gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n216), .A2(KEYINPUT77), .A3(G141gat), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n217), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT2), .ZN(new_n224));
  INV_X1    g023(.A(G155gat), .ZN(new_n225));
  INV_X1    g024(.A(G162gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(new_n225), .B2(new_n226), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n223), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n216), .A2(G141gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n219), .A2(G148gat), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n224), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  XOR2_X1   g031(.A(G155gat), .B(G162gat), .Z(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n229), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n214), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n202), .B1(new_n236), .B2(KEYINPUT85), .ZN(new_n237));
  INV_X1    g036(.A(G22gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n229), .A2(new_n234), .A3(new_n203), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT29), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n213), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n236), .A2(new_n238), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n238), .B1(new_n236), .B2(new_n242), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n237), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n245), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n236), .A2(KEYINPUT85), .ZN(new_n248));
  AND2_X1   g047(.A1(G228gat), .A2(G233gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n247), .A2(new_n250), .A3(new_n243), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n246), .A2(new_n251), .ZN(new_n252));
  XOR2_X1   g051(.A(G78gat), .B(G106gat), .Z(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(KEYINPUT84), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT31), .B(G50gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n246), .A2(new_n251), .A3(new_n256), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G8gat), .B(G36gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(G64gat), .B(G92gat), .ZN(new_n262));
  XOR2_X1   g061(.A(new_n261), .B(new_n262), .Z(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(G169gat), .ZN(new_n265));
  INV_X1    g064(.A(G176gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(new_n266), .A3(KEYINPUT65), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G183gat), .A2(G190gat), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n265), .A2(new_n266), .A3(KEYINPUT65), .A4(KEYINPUT26), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT66), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT66), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n269), .A2(new_n274), .A3(new_n270), .A4(new_n271), .ZN(new_n275));
  INV_X1    g074(.A(G183gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT27), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT27), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(G183gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT64), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(G190gat), .B1(new_n277), .B2(KEYINPUT64), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT28), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT28), .ZN(new_n285));
  NOR3_X1   g084(.A1(new_n280), .A2(new_n285), .A3(G190gat), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n273), .B(new_n275), .C1(new_n284), .C2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT25), .ZN(new_n288));
  OAI21_X1  g087(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(new_n270), .ZN(new_n290));
  NAND3_X1  g089(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  NOR3_X1   g094(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n296));
  OAI22_X1  g095(.A1(new_n295), .A2(new_n296), .B1(new_n265), .B2(new_n266), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n288), .B1(new_n293), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n296), .ZN(new_n299));
  AOI22_X1  g098(.A1(new_n299), .A2(new_n294), .B1(G169gat), .B2(G176gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n300), .A2(KEYINPUT25), .A3(new_n292), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT74), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(G226gat), .ZN(new_n306));
  INV_X1    g105(.A(G233gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n308), .A2(KEYINPUT29), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT74), .B1(new_n287), .B2(new_n302), .ZN(new_n311));
  NOR3_X1   g110(.A1(new_n305), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n308), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n303), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n213), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n211), .B1(new_n208), .B2(new_n209), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n205), .B(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n303), .A2(new_n309), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n305), .A2(new_n311), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n317), .B(new_n318), .C1(new_n319), .C2(new_n313), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n264), .B1(new_n315), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n315), .A2(new_n320), .ZN(new_n322));
  XOR2_X1   g121(.A(new_n263), .B(KEYINPUT75), .Z(new_n323));
  OAI22_X1  g122(.A1(new_n321), .A2(KEYINPUT30), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n321), .A2(KEYINPUT30), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT35), .ZN(new_n327));
  AND2_X1   g126(.A1(G113gat), .A2(G120gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(G113gat), .A2(G120gat), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT67), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(G113gat), .ZN(new_n331));
  INV_X1    g130(.A(G120gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT67), .ZN(new_n334));
  NAND2_X1  g133(.A1(G113gat), .A2(G120gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT1), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n330), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G127gat), .B(G134gat), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT68), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT68), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n338), .A2(new_n343), .A3(new_n340), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n339), .A2(new_n337), .A3(new_n333), .A4(new_n335), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n303), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AND3_X1   g146(.A1(new_n338), .A2(new_n343), .A3(new_n340), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n343), .B1(new_n338), .B2(new_n340), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n346), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n350), .A2(new_n302), .A3(new_n287), .ZN(new_n351));
  AND2_X1   g150(.A1(G227gat), .A2(G233gat), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n347), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT32), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT33), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  XOR2_X1   g155(.A(G15gat), .B(G43gat), .Z(new_n357));
  XNOR2_X1  g156(.A(G71gat), .B(G99gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n357), .B(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n354), .A2(new_n356), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n359), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n353), .B(KEYINPUT32), .C1(new_n355), .C2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT69), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT34), .ZN(new_n365));
  XOR2_X1   g164(.A(new_n365), .B(KEYINPUT70), .Z(new_n366));
  NOR2_X1   g165(.A1(new_n364), .A2(KEYINPUT34), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n347), .A2(new_n351), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n366), .B(new_n368), .C1(new_n369), .C2(new_n352), .ZN(new_n370));
  INV_X1    g169(.A(new_n366), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n352), .B1(new_n347), .B2(new_n351), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n371), .B1(new_n372), .B2(new_n367), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n363), .A2(new_n374), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n360), .A2(new_n362), .A3(new_n370), .A4(new_n373), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n260), .A2(new_n326), .A3(new_n327), .A4(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(G1gat), .B(G29gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n380), .B(KEYINPUT0), .ZN(new_n381));
  XNOR2_X1  g180(.A(G57gat), .B(G85gat), .ZN(new_n382));
  XOR2_X1   g181(.A(new_n381), .B(new_n382), .Z(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n239), .A2(KEYINPUT78), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n235), .A2(KEYINPUT3), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n235), .A2(KEYINPUT78), .A3(KEYINPUT3), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(new_n388), .A3(new_n350), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT5), .ZN(new_n390));
  NAND2_X1  g189(.A1(G225gat), .A2(G233gat), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n391), .B(KEYINPUT79), .Z(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n389), .A2(new_n390), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT4), .ZN(new_n395));
  AND3_X1   g194(.A1(new_n229), .A2(new_n346), .A3(new_n234), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n396), .B1(new_n348), .B2(new_n349), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT80), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n345), .A2(KEYINPUT80), .A3(new_n396), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n395), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n397), .A2(new_n395), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(KEYINPUT81), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n229), .A2(new_n234), .A3(new_n346), .ZN(new_n405));
  AOI211_X1 g204(.A(new_n398), .B(new_n405), .C1(new_n342), .C2(new_n344), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT80), .B1(new_n345), .B2(new_n396), .ZN(new_n407));
  OAI21_X1  g206(.A(KEYINPUT4), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT81), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(new_n409), .A3(new_n402), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n394), .B1(new_n404), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n350), .A2(new_n235), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n399), .A2(new_n412), .A3(new_n400), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n392), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT5), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n399), .A2(new_n395), .A3(new_n400), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n345), .A2(KEYINPUT4), .A3(new_n396), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n389), .A2(new_n393), .A3(new_n417), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n384), .B1(new_n411), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT6), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT82), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n383), .B1(new_n415), .B2(new_n419), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n424), .B1(new_n425), .B2(new_n411), .ZN(new_n426));
  INV_X1    g225(.A(new_n394), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n409), .B1(new_n408), .B2(new_n402), .ZN(new_n428));
  NOR3_X1   g227(.A1(new_n401), .A2(KEYINPUT81), .A3(new_n403), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n390), .B1(new_n413), .B2(new_n392), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n399), .A2(new_n395), .A3(new_n400), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n432), .A2(new_n393), .A3(new_n389), .A4(new_n417), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n384), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n430), .A2(KEYINPUT82), .A3(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT6), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n426), .A2(new_n421), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n379), .B1(new_n423), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT88), .ZN(new_n439));
  INV_X1    g238(.A(new_n326), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT71), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n375), .A2(new_n441), .A3(new_n376), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n363), .A2(KEYINPUT71), .A3(new_n374), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n260), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n426), .A2(new_n435), .A3(new_n436), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT83), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n426), .A2(new_n435), .A3(KEYINPUT83), .A4(new_n436), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n421), .A3(new_n449), .ZN(new_n450));
  AOI211_X1 g249(.A(new_n440), .B(new_n445), .C1(new_n450), .C2(new_n423), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n439), .B1(new_n451), .B2(new_n327), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n450), .A2(new_n423), .ZN(new_n453));
  INV_X1    g252(.A(new_n445), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n453), .A2(new_n326), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n455), .A2(KEYINPUT88), .A3(KEYINPUT35), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n438), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n378), .A2(KEYINPUT72), .A3(KEYINPUT36), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT36), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n459), .B1(new_n442), .B2(new_n443), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT72), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n461), .B1(new_n377), .B2(new_n459), .ZN(new_n462));
  NOR3_X1   g261(.A1(new_n458), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(KEYINPUT86), .B(KEYINPUT37), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n464), .B1(new_n315), .B2(new_n320), .ZN(new_n465));
  OR2_X1    g264(.A1(new_n323), .A2(KEYINPUT38), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OR3_X1    g266(.A1(new_n312), .A2(new_n314), .A3(new_n213), .ZN(new_n468));
  INV_X1    g267(.A(new_n319), .ZN(new_n469));
  AOI22_X1  g268(.A1(new_n469), .A2(new_n308), .B1(new_n309), .B2(new_n303), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n468), .B(KEYINPUT37), .C1(new_n470), .C2(new_n317), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n321), .B1(new_n467), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n423), .A2(new_n437), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT87), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n423), .A2(new_n437), .A3(KEYINPUT87), .A4(new_n472), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT37), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n264), .B1(new_n322), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT38), .B1(new_n478), .B2(new_n465), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n475), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n260), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n421), .B1(new_n324), .B2(new_n325), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT40), .ZN(new_n483));
  OR2_X1    g282(.A1(new_n413), .A2(new_n392), .ZN(new_n484));
  INV_X1    g283(.A(new_n389), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n485), .B1(new_n404), .B2(new_n410), .ZN(new_n486));
  OAI211_X1 g285(.A(KEYINPUT39), .B(new_n484), .C1(new_n486), .C2(new_n393), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n389), .B1(new_n428), .B2(new_n429), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(new_n392), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n487), .B(new_n383), .C1(KEYINPUT39), .C2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n482), .B1(new_n483), .B2(new_n490), .ZN(new_n491));
  OR2_X1    g290(.A1(new_n490), .A2(new_n483), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n481), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n463), .B1(new_n480), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n422), .B1(new_n446), .B2(new_n447), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n495), .A2(new_n449), .B1(KEYINPUT6), .B2(new_n422), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n481), .B1(new_n496), .B2(new_n440), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  OR2_X1    g297(.A1(new_n457), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(G15gat), .B(G22gat), .ZN(new_n500));
  INV_X1    g299(.A(G1gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT16), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n503), .B1(G1gat), .B2(new_n500), .ZN(new_n504));
  INV_X1    g303(.A(G8gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n504), .B(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(KEYINPUT92), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n504), .B(G8gat), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT92), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(G36gat), .ZN(new_n512));
  AND2_X1   g311(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n513));
  NOR2_X1   g312(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(G29gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n516), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(G43gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(G50gat), .ZN(new_n520));
  INV_X1    g319(.A(G50gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(G43gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n520), .A2(new_n522), .A3(KEYINPUT15), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n521), .A2(KEYINPUT90), .A3(G43gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT15), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT90), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n520), .A2(new_n522), .A3(new_n529), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n528), .A2(new_n530), .B1(new_n515), .B2(new_n517), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n525), .B1(new_n531), .B2(new_n524), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n511), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n523), .B1(new_n515), .B2(new_n517), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n529), .B1(new_n519), .B2(G50gat), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n521), .A2(G43gat), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n527), .B(new_n526), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n518), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n534), .B1(new_n538), .B2(new_n523), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n507), .A2(new_n510), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n533), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G229gat), .A2(G233gat), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n542), .B(KEYINPUT13), .Z(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT17), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n545), .B(new_n525), .C1(new_n531), .C2(new_n524), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT91), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT91), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n539), .A2(new_n548), .A3(new_n545), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n532), .A2(KEYINPUT17), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n550), .A2(new_n506), .A3(new_n551), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n552), .A2(new_n540), .A3(KEYINPUT18), .A4(new_n542), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n552), .A2(new_n540), .A3(new_n542), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT18), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n544), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G113gat), .B(G141gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(G197gat), .ZN(new_n559));
  XOR2_X1   g358(.A(KEYINPUT11), .B(G169gat), .Z(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT12), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n557), .A2(KEYINPUT89), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n562), .B1(new_n557), .B2(KEYINPUT89), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AND2_X1   g364(.A1(new_n499), .A2(new_n565), .ZN(new_n566));
  AND2_X1   g365(.A1(KEYINPUT93), .A2(G64gat), .ZN(new_n567));
  NOR2_X1   g366(.A1(KEYINPUT93), .A2(G64gat), .ZN(new_n568));
  OAI21_X1  g367(.A(G57gat), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT94), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT94), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n571), .B(G57gat), .C1(new_n567), .C2(new_n568), .ZN(new_n572));
  INV_X1    g371(.A(G64gat), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n570), .B(new_n572), .C1(G57gat), .C2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(G71gat), .A2(G78gat), .ZN(new_n575));
  OR2_X1    g374(.A1(G71gat), .A2(G78gat), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT9), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G57gat), .B(G64gat), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n575), .B(new_n576), .C1(new_n580), .C2(new_n577), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(KEYINPUT21), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n511), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT97), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT97), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n511), .A2(new_n587), .A3(new_n584), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  XOR2_X1   g388(.A(G127gat), .B(G155gat), .Z(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT96), .ZN(new_n591));
  NAND2_X1  g390(.A1(G231gat), .A2(G233gat), .ZN(new_n592));
  XOR2_X1   g391(.A(new_n592), .B(KEYINPUT95), .Z(new_n593));
  XNOR2_X1  g392(.A(new_n591), .B(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n589), .B(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT21), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(G183gat), .B(G211gat), .Z(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n596), .B(new_n602), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n547), .A2(new_n549), .ZN(new_n604));
  INV_X1    g403(.A(G92gat), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n605), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(G92gat), .ZN(new_n608));
  NOR2_X1   g407(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n606), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(G99gat), .A2(G106gat), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT99), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT99), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n613), .A2(G99gat), .A3(G106gat), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n612), .A2(new_n614), .A3(KEYINPUT8), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G99gat), .B(G106gat), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT101), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n616), .A2(KEYINPUT101), .A3(new_n618), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n610), .A2(new_n615), .A3(new_n617), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT100), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n551), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(KEYINPUT102), .B1(new_n604), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT100), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n623), .B(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT101), .ZN(new_n629));
  AOI211_X1 g428(.A(new_n629), .B(new_n617), .C1(new_n610), .C2(new_n615), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n619), .A2(new_n630), .ZN(new_n631));
  AOI22_X1  g430(.A1(new_n628), .A2(new_n631), .B1(KEYINPUT17), .B2(new_n532), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT102), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n632), .A2(new_n550), .A3(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n628), .A2(new_n631), .A3(new_n539), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT103), .ZN(new_n636));
  NAND3_X1  g435(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n636), .B1(new_n635), .B2(new_n637), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n626), .B(new_n634), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G190gat), .B(G218gat), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n642), .ZN(new_n644));
  AND3_X1   g443(.A1(new_n632), .A2(new_n550), .A3(new_n633), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n633), .B1(new_n632), .B2(new_n550), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n640), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n638), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n644), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT98), .ZN(new_n652));
  XNOR2_X1  g451(.A(G134gat), .B(G162gat), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n652), .B(new_n653), .Z(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  OR3_X1    g454(.A1(new_n643), .A2(new_n650), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT105), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n647), .A2(new_n649), .A3(new_n644), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n658), .B1(new_n650), .B2(KEYINPUT104), .ZN(new_n659));
  OR3_X1    g458(.A1(new_n641), .A2(KEYINPUT104), .A3(new_n642), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n657), .B1(new_n661), .B2(new_n655), .ZN(new_n662));
  AOI211_X1 g461(.A(KEYINPUT105), .B(new_n654), .C1(new_n659), .C2(new_n660), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n603), .B(new_n656), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT106), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(KEYINPUT104), .B1(new_n641), .B2(new_n642), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n667), .A2(new_n643), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n641), .A2(KEYINPUT104), .A3(new_n642), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n655), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(KEYINPUT105), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n661), .A2(new_n657), .A3(new_n655), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n673), .A2(KEYINPUT106), .A3(new_n603), .A4(new_n656), .ZN(new_n674));
  XNOR2_X1  g473(.A(G120gat), .B(G148gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(G176gat), .B(G204gat), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n675), .B(new_n676), .Z(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n616), .A2(new_n618), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n583), .A2(new_n623), .A3(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n582), .B1(new_n622), .B2(new_n624), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(G230gat), .A2(G233gat), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT107), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT10), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n680), .A2(new_n689), .A3(new_n681), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n583), .A2(KEYINPUT10), .A3(new_n628), .A4(new_n631), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n684), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n678), .B1(new_n688), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n692), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n687), .A2(new_n677), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n666), .A2(new_n674), .A3(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT108), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n666), .A2(new_n674), .A3(KEYINPUT108), .A4(new_n697), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n566), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n703), .A2(new_n453), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(new_n501), .ZN(G1324gat));
  NOR2_X1   g504(.A1(new_n703), .A2(new_n326), .ZN(new_n706));
  XNOR2_X1  g505(.A(KEYINPUT109), .B(KEYINPUT16), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(new_n505), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT42), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n706), .A2(KEYINPUT42), .A3(new_n708), .ZN(new_n712));
  OAI21_X1  g511(.A(G8gat), .B1(new_n703), .B2(new_n326), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(G1325gat));
  INV_X1    g513(.A(new_n703), .ZN(new_n715));
  AOI21_X1  g514(.A(G15gat), .B1(new_n715), .B2(new_n378), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n463), .A2(G15gat), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n717), .B(KEYINPUT110), .Z(new_n718));
  AOI21_X1  g517(.A(new_n716), .B1(new_n715), .B2(new_n718), .ZN(G1326gat));
  INV_X1    g518(.A(KEYINPUT111), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n720), .B1(new_n703), .B2(new_n260), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n566), .A2(KEYINPUT111), .A3(new_n481), .A4(new_n702), .ZN(new_n722));
  XNOR2_X1  g521(.A(KEYINPUT43), .B(G22gat), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n723), .B1(new_n721), .B2(new_n722), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n724), .A2(new_n725), .ZN(G1327gat));
  NAND2_X1  g525(.A1(new_n673), .A2(new_n656), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n440), .B1(new_n450), .B2(new_n423), .ZN(new_n728));
  OAI21_X1  g527(.A(KEYINPUT112), .B1(new_n728), .B2(new_n260), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT112), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n730), .B(new_n481), .C1(new_n496), .C2(new_n440), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n494), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n727), .B1(new_n457), .B2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI211_X1 g534(.A(KEYINPUT44), .B(new_n727), .C1(new_n457), .C2(new_n498), .ZN(new_n736));
  INV_X1    g535(.A(new_n603), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n697), .ZN(new_n738));
  INV_X1    g537(.A(new_n565), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n735), .A2(new_n736), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(G29gat), .B1(new_n741), .B2(new_n453), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n743));
  INV_X1    g542(.A(new_n727), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n744), .A2(new_n738), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n499), .A2(new_n565), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n453), .A2(G29gat), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n743), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n566), .A2(KEYINPUT45), .A3(new_n745), .A4(new_n747), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n742), .A2(new_n749), .A3(new_n750), .ZN(G1328gat));
  NOR3_X1   g550(.A1(new_n746), .A2(G36gat), .A3(new_n326), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT46), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(KEYINPUT113), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(G36gat), .B1(new_n741), .B2(new_n326), .ZN(new_n755));
  XNOR2_X1  g554(.A(KEYINPUT113), .B(KEYINPUT46), .ZN(new_n756));
  OAI211_X1 g555(.A(new_n754), .B(new_n755), .C1(new_n752), .C2(new_n756), .ZN(G1329gat));
  OAI21_X1  g556(.A(new_n519), .B1(new_n746), .B2(new_n377), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n463), .A2(G43gat), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n758), .B1(new_n741), .B2(new_n759), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g560(.A(new_n521), .B1(new_n746), .B2(new_n260), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n481), .A2(G50gat), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n762), .B1(new_n741), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT48), .ZN(G1331gat));
  OR2_X1    g564(.A1(new_n457), .A2(new_n732), .ZN(new_n766));
  AND4_X1   g565(.A1(new_n739), .A2(new_n666), .A3(new_n674), .A4(new_n696), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n496), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g570(.A(new_n326), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(KEYINPUT114), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n773), .A2(KEYINPUT114), .ZN(new_n776));
  OAI22_X1  g575(.A1(new_n775), .A2(new_n776), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n777));
  INV_X1    g576(.A(new_n776), .ZN(new_n778));
  NOR2_X1   g577(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n778), .A2(new_n774), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n777), .A2(new_n780), .ZN(G1333gat));
  OR3_X1    g580(.A1(new_n458), .A2(new_n460), .A3(new_n462), .ZN(new_n782));
  OAI21_X1  g581(.A(G71gat), .B1(new_n768), .B2(new_n782), .ZN(new_n783));
  OR2_X1    g582(.A1(new_n377), .A2(G71gat), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n783), .B1(new_n768), .B2(new_n784), .ZN(new_n785));
  XOR2_X1   g584(.A(new_n785), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g585(.A1(new_n768), .A2(new_n260), .ZN(new_n787));
  XOR2_X1   g586(.A(KEYINPUT115), .B(G78gat), .Z(new_n788));
  XNOR2_X1  g587(.A(new_n787), .B(new_n788), .ZN(G1335gat));
  NOR2_X1   g588(.A1(new_n603), .A2(new_n565), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n766), .A2(KEYINPUT51), .A3(new_n727), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT116), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n727), .B(new_n790), .C1(new_n457), .C2(new_n732), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT51), .ZN(new_n794));
  OR3_X1    g593(.A1(new_n793), .A2(KEYINPUT116), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n792), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n453), .A2(G85gat), .A3(new_n697), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n790), .A2(new_n696), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n735), .A2(new_n736), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(G85gat), .B1(new_n802), .B2(new_n453), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n799), .A2(new_n803), .ZN(G1336gat));
  NOR3_X1   g603(.A1(new_n697), .A2(G92gat), .A3(new_n326), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n797), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n735), .A2(new_n440), .A3(new_n736), .A4(new_n801), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT52), .B1(new_n807), .B2(G92gat), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT117), .ZN(new_n810));
  AND3_X1   g609(.A1(new_n807), .A2(new_n810), .A3(G92gat), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n810), .B1(new_n807), .B2(G92gat), .ZN(new_n812));
  INV_X1    g611(.A(new_n805), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n813), .B1(new_n791), .B2(new_n796), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n811), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n809), .B1(new_n815), .B2(new_n816), .ZN(G1337gat));
  NOR3_X1   g616(.A1(new_n697), .A2(G99gat), .A3(new_n377), .ZN(new_n818));
  XOR2_X1   g617(.A(new_n818), .B(KEYINPUT118), .Z(new_n819));
  NAND2_X1  g618(.A1(new_n797), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(G99gat), .B1(new_n802), .B2(new_n782), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(G1338gat));
  NOR3_X1   g621(.A1(new_n697), .A2(G106gat), .A3(new_n260), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n797), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n735), .A2(new_n481), .A3(new_n736), .A4(new_n801), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(G106gat), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n791), .A2(new_n796), .ZN(new_n829));
  AOI22_X1  g628(.A1(new_n829), .A2(new_n823), .B1(new_n825), .B2(G106gat), .ZN(new_n830));
  OAI22_X1  g629(.A1(new_n824), .A2(new_n828), .B1(new_n827), .B2(new_n830), .ZN(G1339gat));
  NAND3_X1  g630(.A1(new_n690), .A2(new_n684), .A3(new_n691), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n694), .A2(KEYINPUT54), .A3(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n677), .B1(new_n692), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n833), .A2(KEYINPUT55), .A3(new_n835), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n836), .A2(new_n695), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n833), .A2(new_n835), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT55), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n541), .A2(new_n543), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n542), .B1(new_n552), .B2(new_n540), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n561), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n544), .A2(new_n556), .A3(new_n553), .A4(new_n562), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XOR2_X1   g645(.A(new_n846), .B(KEYINPUT119), .Z(new_n847));
  AND3_X1   g646(.A1(new_n727), .A2(new_n841), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n837), .A2(new_n565), .A3(new_n840), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n696), .A2(new_n846), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n727), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n737), .B1(new_n848), .B2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n666), .A2(new_n674), .A3(new_n739), .A4(new_n697), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n853), .B1(new_n852), .B2(new_n854), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n856), .A2(new_n481), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n453), .A2(new_n440), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n378), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n861), .A2(new_n331), .A3(new_n739), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n860), .A2(new_n444), .A3(new_n565), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n862), .B1(new_n331), .B2(new_n863), .ZN(G1340gat));
  NOR3_X1   g663(.A1(new_n861), .A2(new_n332), .A3(new_n697), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n860), .A2(new_n444), .A3(new_n696), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n865), .B1(new_n332), .B2(new_n866), .ZN(G1341gat));
  OAI21_X1  g666(.A(G127gat), .B1(new_n861), .B2(new_n737), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n858), .A2(new_n444), .A3(new_n859), .ZN(new_n869));
  OR2_X1    g668(.A1(new_n737), .A2(G127gat), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(G1342gat));
  OAI21_X1  g670(.A(G134gat), .B1(new_n861), .B2(new_n744), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n744), .A2(G134gat), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  OR3_X1    g673(.A1(new_n869), .A2(KEYINPUT56), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(KEYINPUT56), .B1(new_n869), .B2(new_n874), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n872), .A2(new_n875), .A3(new_n876), .ZN(G1343gat));
  NAND2_X1  g676(.A1(new_n782), .A2(new_n481), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n878), .B(KEYINPUT123), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n859), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n856), .A2(new_n880), .A3(new_n857), .ZN(new_n881));
  AOI21_X1  g680(.A(G141gat), .B1(new_n881), .B2(new_n565), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n859), .A2(new_n782), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n852), .A2(new_n854), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(KEYINPUT120), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n481), .A3(new_n855), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT57), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n840), .B(KEYINPUT121), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n837), .A2(new_n565), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n850), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n744), .A2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n727), .A2(new_n841), .A3(new_n847), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n744), .A2(new_n891), .A3(KEYINPUT122), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n854), .B1(new_n897), .B2(new_n603), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n260), .A2(new_n887), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n883), .B1(new_n888), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n739), .A2(new_n219), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n882), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT124), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT58), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT58), .ZN(new_n906));
  INV_X1    g705(.A(new_n902), .ZN(new_n907));
  AOI211_X1 g706(.A(new_n883), .B(new_n907), .C1(new_n888), .C2(new_n900), .ZN(new_n908));
  OAI211_X1 g707(.A(KEYINPUT124), .B(new_n906), .C1(new_n908), .C2(new_n882), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n905), .A2(new_n909), .ZN(G1344gat));
  NAND3_X1  g709(.A1(new_n881), .A2(new_n216), .A3(new_n696), .ZN(new_n911));
  XOR2_X1   g710(.A(KEYINPUT125), .B(KEYINPUT59), .Z(new_n912));
  INV_X1    g711(.A(new_n883), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n885), .A2(new_n855), .A3(new_n899), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n700), .A2(new_n739), .A3(new_n701), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n892), .A2(new_n895), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n737), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(KEYINPUT57), .B1(new_n918), .B2(new_n481), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT126), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n914), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AOI211_X1 g720(.A(KEYINPUT126), .B(KEYINPUT57), .C1(new_n918), .C2(new_n481), .ZN(new_n922));
  OAI211_X1 g721(.A(new_n696), .B(new_n913), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n912), .B1(new_n923), .B2(G148gat), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n216), .A2(KEYINPUT59), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n925), .B1(new_n901), .B2(new_n696), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n911), .B1(new_n924), .B2(new_n926), .ZN(G1345gat));
  INV_X1    g726(.A(new_n901), .ZN(new_n928));
  OAI21_X1  g727(.A(G155gat), .B1(new_n928), .B2(new_n737), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n881), .A2(new_n225), .A3(new_n603), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1346gat));
  OAI21_X1  g730(.A(G162gat), .B1(new_n928), .B2(new_n744), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n881), .A2(new_n226), .A3(new_n727), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1347gat));
  NOR2_X1   g733(.A1(new_n496), .A2(new_n326), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n936), .A2(new_n377), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n858), .A2(new_n937), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n938), .A2(new_n265), .A3(new_n739), .ZN(new_n939));
  NOR4_X1   g738(.A1(new_n856), .A2(new_n857), .A3(new_n445), .A4(new_n936), .ZN(new_n940));
  AOI21_X1  g739(.A(G169gat), .B1(new_n940), .B2(new_n565), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n939), .A2(new_n941), .ZN(G1348gat));
  OAI21_X1  g741(.A(G176gat), .B1(new_n938), .B2(new_n697), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n940), .A2(new_n266), .A3(new_n696), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1349gat));
  OAI21_X1  g744(.A(G183gat), .B1(new_n938), .B2(new_n737), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT127), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n737), .A2(new_n280), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n947), .B1(new_n940), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g750(.A(G190gat), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n940), .A2(new_n952), .A3(new_n727), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n858), .A2(new_n727), .A3(new_n937), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT61), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n954), .A2(new_n955), .A3(G190gat), .ZN(new_n956));
  INV_X1    g755(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n955), .B1(new_n954), .B2(G190gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n953), .B1(new_n957), .B2(new_n958), .ZN(G1351gat));
  NOR2_X1   g758(.A1(new_n936), .A2(new_n463), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n885), .A2(new_n481), .A3(new_n855), .A4(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  AOI21_X1  g761(.A(G197gat), .B1(new_n962), .B2(new_n565), .ZN(new_n963));
  OR2_X1    g762(.A1(new_n921), .A2(new_n922), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n964), .A2(new_n960), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n739), .A2(new_n206), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n963), .B1(new_n965), .B2(new_n966), .ZN(G1352gat));
  NAND2_X1  g766(.A1(new_n696), .A2(new_n207), .ZN(new_n968));
  OR2_X1    g767(.A1(new_n961), .A2(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT62), .ZN(new_n970));
  XNOR2_X1  g769(.A(new_n969), .B(new_n970), .ZN(new_n971));
  AND3_X1   g770(.A1(new_n964), .A2(new_n696), .A3(new_n960), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n971), .B1(new_n972), .B2(new_n207), .ZN(G1353gat));
  OR3_X1    g772(.A1(new_n961), .A2(G211gat), .A3(new_n737), .ZN(new_n974));
  OAI211_X1 g773(.A(new_n603), .B(new_n960), .C1(new_n921), .C2(new_n922), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n975), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n976));
  AOI21_X1  g775(.A(KEYINPUT63), .B1(new_n975), .B2(G211gat), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n974), .B1(new_n976), .B2(new_n977), .ZN(G1354gat));
  NAND3_X1  g777(.A1(new_n964), .A2(new_n727), .A3(new_n960), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(G218gat), .ZN(new_n980));
  OR3_X1    g779(.A1(new_n961), .A2(G218gat), .A3(new_n744), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(G1355gat));
endmodule


