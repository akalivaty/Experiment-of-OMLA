

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748;

  XNOR2_X1 U373 ( .A(G902), .B(KEYINPUT15), .ZN(n614) );
  XNOR2_X2 U374 ( .A(n582), .B(n581), .ZN(n596) );
  XNOR2_X2 U375 ( .A(n540), .B(n357), .ZN(n389) );
  NOR2_X2 U376 ( .A1(n710), .A2(n543), .ZN(n540) );
  XNOR2_X1 U377 ( .A(n360), .B(n359), .ZN(n709) );
  NOR2_X1 U378 ( .A1(n562), .A2(n561), .ZN(n466) );
  INV_X1 U379 ( .A(n594), .ZN(n695) );
  NOR2_X1 U380 ( .A1(n716), .A2(n715), .ZN(n396) );
  AND2_X1 U381 ( .A1(n401), .A2(n405), .ZN(n403) );
  AND2_X1 U382 ( .A1(n384), .A2(n382), .ZN(n388) );
  XNOR2_X1 U383 ( .A(n362), .B(KEYINPUT32), .ZN(n747) );
  NOR2_X1 U384 ( .A1(n709), .A2(n397), .ZN(n583) );
  OR2_X1 U385 ( .A1(n542), .A2(n435), .ZN(n436) );
  XNOR2_X1 U386 ( .A(n427), .B(n426), .ZN(n531) );
  OR2_X1 U387 ( .A1(n617), .A2(G902), .ZN(n512) );
  XNOR2_X1 U388 ( .A(n486), .B(G472), .ZN(n594) );
  OR2_X1 U389 ( .A1(n497), .A2(n469), .ZN(n471) );
  XNOR2_X1 U390 ( .A(n478), .B(n477), .ZN(n508) );
  XNOR2_X1 U391 ( .A(n443), .B(G140), .ZN(n444) );
  XNOR2_X1 U392 ( .A(n456), .B(G134), .ZN(n478) );
  XNOR2_X1 U393 ( .A(KEYINPUT68), .B(G131), .ZN(n476) );
  NAND2_X2 U394 ( .A1(n404), .A2(n402), .ZN(n717) );
  NAND2_X1 U395 ( .A1(n403), .A2(n626), .ZN(n402) );
  XNOR2_X2 U396 ( .A(n517), .B(KEYINPUT66), .ZN(n579) );
  BUF_X1 U397 ( .A(n580), .Z(n352) );
  NAND2_X1 U398 ( .A1(n353), .A2(n379), .ZN(n378) );
  INV_X1 U399 ( .A(KEYINPUT104), .ZN(n379) );
  NAND2_X1 U400 ( .A1(n388), .A2(n386), .ZN(n568) );
  NAND2_X1 U401 ( .A1(n387), .A2(KEYINPUT46), .ZN(n386) );
  NAND2_X1 U402 ( .A1(n409), .A2(n406), .ZN(n592) );
  AND2_X1 U403 ( .A1(n747), .A2(n361), .ZN(n406) );
  XOR2_X1 U404 ( .A(KEYINPUT12), .B(G104), .Z(n438) );
  XNOR2_X1 U405 ( .A(G143), .B(G122), .ZN(n437) );
  XOR2_X1 U406 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n440) );
  NOR2_X1 U407 ( .A1(n399), .A2(G953), .ZN(n398) );
  INV_X1 U408 ( .A(G224), .ZN(n399) );
  NOR2_X1 U409 ( .A1(n730), .A2(n614), .ZN(n369) );
  XNOR2_X1 U410 ( .A(n368), .B(n367), .ZN(n685) );
  INV_X1 U411 ( .A(KEYINPUT107), .ZN(n367) );
  NAND2_X1 U412 ( .A1(n681), .A2(n682), .ZN(n368) );
  INV_X1 U413 ( .A(KEYINPUT33), .ZN(n359) );
  INV_X1 U414 ( .A(n682), .ZN(n364) );
  INV_X1 U415 ( .A(KEYINPUT3), .ZN(n419) );
  XNOR2_X1 U416 ( .A(G119), .B(G101), .ZN(n417) );
  INV_X2 U417 ( .A(G953), .ZN(n739) );
  AND2_X1 U418 ( .A1(n566), .A2(n383), .ZN(n382) );
  NAND2_X1 U419 ( .A1(G234), .A2(G237), .ZN(n430) );
  OR2_X1 U420 ( .A1(G237), .A2(G902), .ZN(n428) );
  XOR2_X1 U421 ( .A(KEYINPUT5), .B(KEYINPUT75), .Z(n480) );
  INV_X1 U422 ( .A(KEYINPUT48), .ZN(n567) );
  NOR2_X1 U423 ( .A1(G237), .A2(G953), .ZN(n447) );
  INV_X1 U424 ( .A(KEYINPUT74), .ZN(n581) );
  NAND2_X1 U425 ( .A1(n380), .A2(n376), .ZN(n375) );
  NAND2_X1 U426 ( .A1(n378), .A2(n377), .ZN(n376) );
  NAND2_X1 U427 ( .A1(n526), .A2(KEYINPUT104), .ZN(n377) );
  NAND2_X1 U428 ( .A1(n374), .A2(n373), .ZN(n372) );
  NAND2_X1 U429 ( .A1(n526), .A2(n379), .ZN(n373) );
  NAND2_X1 U430 ( .A1(n353), .A2(KEYINPUT104), .ZN(n374) );
  OR2_X1 U431 ( .A1(n534), .A2(n526), .ZN(n392) );
  XNOR2_X1 U432 ( .A(G110), .B(KEYINPUT92), .ZN(n492) );
  XNOR2_X1 U433 ( .A(KEYINPUT24), .B(G119), .ZN(n493) );
  XNOR2_X1 U434 ( .A(KEYINPUT93), .B(KEYINPUT23), .ZN(n488) );
  XNOR2_X1 U435 ( .A(G116), .B(G122), .ZN(n455) );
  XNOR2_X1 U436 ( .A(G113), .B(KEYINPUT97), .ZN(n439) );
  XOR2_X1 U437 ( .A(G146), .B(G140), .Z(n503) );
  XOR2_X1 U438 ( .A(KEYINPUT17), .B(KEYINPUT85), .Z(n411) );
  XNOR2_X1 U439 ( .A(n400), .B(n398), .ZN(n412) );
  XNOR2_X1 U440 ( .A(KEYINPUT4), .B(KEYINPUT18), .ZN(n400) );
  XNOR2_X1 U441 ( .A(n366), .B(n356), .ZN(n710) );
  NOR2_X1 U442 ( .A1(n685), .A2(n684), .ZN(n366) );
  XNOR2_X1 U443 ( .A(n530), .B(KEYINPUT77), .ZN(n564) );
  NAND2_X1 U444 ( .A1(n390), .A2(n391), .ZN(n530) );
  AND2_X1 U445 ( .A1(n529), .A2(n392), .ZN(n391) );
  NAND2_X1 U446 ( .A1(n375), .A2(n371), .ZN(n390) );
  XNOR2_X1 U447 ( .A(n363), .B(n354), .ZN(n542) );
  NOR2_X1 U448 ( .A1(n531), .A2(n364), .ZN(n363) );
  NOR2_X1 U449 ( .A1(G902), .A2(n645), .ZN(n486) );
  XNOR2_X1 U450 ( .A(n421), .B(G122), .ZN(n422) );
  XOR2_X1 U451 ( .A(KEYINPUT16), .B(KEYINPUT73), .Z(n421) );
  AND2_X1 U452 ( .A1(n620), .A2(G953), .ZN(n722) );
  NAND2_X1 U453 ( .A1(n569), .A2(n664), .ZN(n533) );
  NOR2_X1 U454 ( .A1(n573), .A2(n571), .ZN(n553) );
  NAND2_X1 U455 ( .A1(n589), .A2(n407), .ZN(n362) );
  NOR2_X1 U456 ( .A1(n542), .A2(n543), .ZN(n665) );
  INV_X1 U457 ( .A(KEYINPUT53), .ZN(n393) );
  INV_X1 U458 ( .A(G137), .ZN(n365) );
  INV_X1 U459 ( .A(n361), .ZN(n658) );
  NAND2_X1 U460 ( .A1(n534), .A2(n526), .ZN(n353) );
  XOR2_X1 U461 ( .A(n429), .B(KEYINPUT19), .Z(n354) );
  XNOR2_X1 U462 ( .A(KEYINPUT6), .B(n594), .ZN(n590) );
  XNOR2_X1 U463 ( .A(n532), .B(KEYINPUT39), .ZN(n569) );
  AND2_X1 U464 ( .A1(n586), .A2(n585), .ZN(n355) );
  XNOR2_X1 U465 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n356) );
  XOR2_X1 U466 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n357) );
  NAND2_X1 U467 ( .A1(n358), .A2(n584), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n583), .B(KEYINPUT34), .ZN(n358) );
  NAND2_X1 U469 ( .A1(n596), .A2(n590), .ZN(n360) );
  XNOR2_X1 U470 ( .A(n502), .B(KEYINPUT91), .ZN(n504) );
  NAND2_X1 U471 ( .A1(n370), .A2(n369), .ZN(n401) );
  NOR2_X2 U472 ( .A1(n648), .A2(n722), .ZN(n651) );
  NOR2_X2 U473 ( .A1(n641), .A2(n722), .ZN(n642) );
  XNOR2_X1 U474 ( .A(n420), .B(n419), .ZN(n479) );
  NAND2_X1 U475 ( .A1(n589), .A2(n355), .ZN(n361) );
  NOR2_X1 U476 ( .A1(n389), .A2(KEYINPUT46), .ZN(n385) );
  XNOR2_X1 U477 ( .A(n389), .B(n365), .ZN(G39) );
  NOR2_X2 U478 ( .A1(n738), .A2(n730), .ZN(n678) );
  INV_X1 U479 ( .A(n738), .ZN(n370) );
  NAND2_X1 U480 ( .A1(n678), .A2(KEYINPUT2), .ZN(n626) );
  NAND2_X1 U481 ( .A1(n678), .A2(n610), .ZN(n613) );
  NAND2_X1 U482 ( .A1(n593), .A2(n372), .ZN(n371) );
  INV_X1 U483 ( .A(n593), .ZN(n380) );
  NAND2_X1 U484 ( .A1(n615), .A2(n626), .ZN(n404) );
  XNOR2_X2 U485 ( .A(n573), .B(KEYINPUT38), .ZN(n681) );
  XNOR2_X1 U486 ( .A(n381), .B(G137), .ZN(n489) );
  XNOR2_X2 U487 ( .A(G128), .B(KEYINPUT80), .ZN(n381) );
  NAND2_X1 U488 ( .A1(n389), .A2(KEYINPUT46), .ZN(n383) );
  NAND2_X1 U489 ( .A1(n541), .A2(n385), .ZN(n384) );
  XNOR2_X2 U490 ( .A(n533), .B(KEYINPUT40), .ZN(n541) );
  INV_X1 U491 ( .A(n541), .ZN(n387) );
  XNOR2_X1 U492 ( .A(n394), .B(n393), .ZN(G75) );
  NAND2_X1 U493 ( .A1(n395), .A2(n739), .ZN(n394) );
  XNOR2_X1 U494 ( .A(n396), .B(KEYINPUT122), .ZN(n395) );
  NOR2_X1 U495 ( .A1(n397), .A2(n684), .ZN(n472) );
  NOR2_X1 U496 ( .A1(n397), .A2(n700), .ZN(n597) );
  OR2_X1 U497 ( .A1(n397), .A2(n595), .ZN(n654) );
  XNOR2_X2 U498 ( .A(n436), .B(KEYINPUT0), .ZN(n397) );
  OR2_X1 U499 ( .A1(n403), .A2(n615), .ZN(n629) );
  INV_X1 U500 ( .A(KEYINPUT82), .ZN(n405) );
  AND2_X1 U501 ( .A1(n588), .A2(n408), .ZN(n407) );
  INV_X1 U502 ( .A(n590), .ZN(n408) );
  INV_X1 U503 ( .A(n746), .ZN(n409) );
  XNOR2_X2 U504 ( .A(n410), .B(KEYINPUT35), .ZN(n746) );
  NOR2_X2 U505 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X2 U506 ( .A(n445), .B(n444), .ZN(n736) );
  XNOR2_X1 U507 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U508 ( .A(n508), .B(n479), .ZN(n485) );
  INV_X1 U509 ( .A(KEYINPUT78), .ZN(n526) );
  XNOR2_X1 U510 ( .A(n412), .B(n411), .ZN(n414) );
  XNOR2_X2 U511 ( .A(G146), .B(G125), .ZN(n445) );
  XNOR2_X2 U512 ( .A(G128), .B(G143), .ZN(n456) );
  XOR2_X1 U513 ( .A(n445), .B(n456), .Z(n413) );
  XNOR2_X1 U514 ( .A(n414), .B(n413), .ZN(n416) );
  XOR2_X1 U515 ( .A(G107), .B(G104), .Z(n415) );
  XNOR2_X1 U516 ( .A(n415), .B(G110), .ZN(n723) );
  XNOR2_X1 U517 ( .A(n723), .B(KEYINPUT70), .ZN(n507) );
  XNOR2_X1 U518 ( .A(n416), .B(n507), .ZN(n423) );
  XOR2_X1 U519 ( .A(G113), .B(G116), .Z(n418) );
  XNOR2_X1 U520 ( .A(n418), .B(n417), .ZN(n420) );
  XNOR2_X1 U521 ( .A(n479), .B(n422), .ZN(n724) );
  XNOR2_X1 U522 ( .A(n423), .B(n724), .ZN(n631) );
  NAND2_X1 U523 ( .A1(n631), .A2(n614), .ZN(n427) );
  XOR2_X1 U524 ( .A(KEYINPUT87), .B(KEYINPUT86), .Z(n425) );
  NAND2_X1 U525 ( .A1(G210), .A2(n428), .ZN(n424) );
  XNOR2_X1 U526 ( .A(n425), .B(n424), .ZN(n426) );
  NAND2_X1 U527 ( .A1(G214), .A2(n428), .ZN(n682) );
  XOR2_X1 U528 ( .A(KEYINPUT65), .B(KEYINPUT79), .Z(n429) );
  XNOR2_X1 U529 ( .A(n430), .B(KEYINPUT14), .ZN(n432) );
  NAND2_X1 U530 ( .A1(G952), .A2(n432), .ZN(n708) );
  NOR2_X1 U531 ( .A1(n708), .A2(G953), .ZN(n523) );
  NOR2_X1 U532 ( .A1(G898), .A2(n739), .ZN(n431) );
  XOR2_X1 U533 ( .A(KEYINPUT88), .B(n431), .Z(n725) );
  NAND2_X1 U534 ( .A1(G902), .A2(n432), .ZN(n520) );
  NOR2_X1 U535 ( .A1(n725), .A2(n520), .ZN(n433) );
  NOR2_X1 U536 ( .A1(n523), .A2(n433), .ZN(n434) );
  XOR2_X1 U537 ( .A(KEYINPUT89), .B(n434), .Z(n435) );
  XNOR2_X1 U538 ( .A(n438), .B(n437), .ZN(n442) );
  XNOR2_X1 U539 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U540 ( .A(n442), .B(n441), .ZN(n446) );
  INV_X1 U541 ( .A(KEYINPUT10), .ZN(n443) );
  XNOR2_X1 U542 ( .A(n446), .B(n736), .ZN(n451) );
  XNOR2_X1 U543 ( .A(n447), .B(KEYINPUT76), .ZN(n481) );
  NAND2_X1 U544 ( .A1(n481), .A2(G214), .ZN(n449) );
  XNOR2_X1 U545 ( .A(n476), .B(KEYINPUT11), .ZN(n448) );
  XNOR2_X1 U546 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U547 ( .A(n451), .B(n450), .ZN(n638) );
  NOR2_X1 U548 ( .A1(G902), .A2(n638), .ZN(n453) );
  XNOR2_X1 U549 ( .A(KEYINPUT98), .B(KEYINPUT13), .ZN(n452) );
  XNOR2_X1 U550 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U551 ( .A(n454), .B(G475), .ZN(n562) );
  XNOR2_X1 U552 ( .A(n455), .B(G107), .ZN(n457) );
  XOR2_X1 U553 ( .A(n457), .B(n478), .Z(n461) );
  NAND2_X1 U554 ( .A1(n739), .A2(G234), .ZN(n459) );
  XNOR2_X1 U555 ( .A(KEYINPUT8), .B(KEYINPUT67), .ZN(n458) );
  XNOR2_X1 U556 ( .A(n459), .B(n458), .ZN(n487) );
  NAND2_X1 U557 ( .A1(n487), .A2(G217), .ZN(n460) );
  XNOR2_X1 U558 ( .A(n461), .B(n460), .ZN(n463) );
  XOR2_X1 U559 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n462) );
  XNOR2_X1 U560 ( .A(n463), .B(n462), .ZN(n718) );
  NOR2_X1 U561 ( .A1(G902), .A2(n718), .ZN(n465) );
  XNOR2_X1 U562 ( .A(KEYINPUT99), .B(G478), .ZN(n464) );
  XNOR2_X1 U563 ( .A(n465), .B(n464), .ZN(n561) );
  XOR2_X1 U564 ( .A(n466), .B(KEYINPUT100), .Z(n684) );
  NAND2_X1 U565 ( .A1(n614), .A2(G234), .ZN(n468) );
  INV_X1 U566 ( .A(KEYINPUT20), .ZN(n467) );
  XNOR2_X1 U567 ( .A(n468), .B(n467), .ZN(n497) );
  INV_X1 U568 ( .A(G221), .ZN(n469) );
  INV_X1 U569 ( .A(KEYINPUT21), .ZN(n470) );
  XNOR2_X1 U570 ( .A(n471), .B(n470), .ZN(n691) );
  NAND2_X1 U571 ( .A1(n472), .A2(n691), .ZN(n474) );
  XOR2_X1 U572 ( .A(KEYINPUT72), .B(KEYINPUT22), .Z(n473) );
  XNOR2_X2 U573 ( .A(n474), .B(n473), .ZN(n589) );
  XNOR2_X1 U574 ( .A(G137), .B(KEYINPUT4), .ZN(n475) );
  XNOR2_X1 U575 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U576 ( .A(n480), .B(G146), .ZN(n483) );
  NAND2_X1 U577 ( .A1(G210), .A2(n481), .ZN(n482) );
  XNOR2_X1 U578 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U579 ( .A(n485), .B(n484), .ZN(n645) );
  NAND2_X1 U580 ( .A1(n487), .A2(G221), .ZN(n491) );
  XNOR2_X1 U581 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U582 ( .A(n491), .B(n490), .ZN(n496) );
  XNOR2_X1 U583 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U584 ( .A(n736), .B(n494), .ZN(n495) );
  XNOR2_X1 U585 ( .A(n496), .B(n495), .ZN(n622) );
  OR2_X2 U586 ( .A1(n622), .A2(G902), .ZN(n501) );
  INV_X1 U587 ( .A(n497), .ZN(n498) );
  NAND2_X1 U588 ( .A1(n498), .A2(G217), .ZN(n499) );
  XNOR2_X1 U589 ( .A(n499), .B(KEYINPUT25), .ZN(n500) );
  XNOR2_X2 U590 ( .A(n501), .B(n500), .ZN(n516) );
  INV_X1 U591 ( .A(n516), .ZN(n692) );
  NAND2_X1 U592 ( .A1(n408), .A2(n692), .ZN(n513) );
  NAND2_X1 U593 ( .A1(G227), .A2(n739), .ZN(n502) );
  XNOR2_X1 U594 ( .A(n505), .B(G101), .ZN(n506) );
  XNOR2_X1 U595 ( .A(n506), .B(n507), .ZN(n509) );
  XNOR2_X1 U596 ( .A(n508), .B(KEYINPUT90), .ZN(n737) );
  XNOR2_X1 U597 ( .A(n509), .B(n737), .ZN(n617) );
  INV_X1 U598 ( .A(KEYINPUT69), .ZN(n510) );
  XNOR2_X1 U599 ( .A(n510), .B(G469), .ZN(n511) );
  XNOR2_X2 U600 ( .A(n512), .B(n511), .ZN(n538) );
  XNOR2_X1 U601 ( .A(n538), .B(KEYINPUT1), .ZN(n580) );
  NOR2_X1 U602 ( .A1(n513), .A2(n352), .ZN(n514) );
  NAND2_X1 U603 ( .A1(n589), .A2(n514), .ZN(n601) );
  XNOR2_X1 U604 ( .A(n601), .B(G101), .ZN(G3) );
  INV_X1 U605 ( .A(n691), .ZN(n515) );
  NAND2_X1 U606 ( .A1(n579), .A2(n538), .ZN(n519) );
  INV_X1 U607 ( .A(KEYINPUT94), .ZN(n518) );
  XNOR2_X2 U608 ( .A(n519), .B(n518), .ZN(n593) );
  OR2_X1 U609 ( .A1(n739), .A2(n520), .ZN(n521) );
  XOR2_X1 U610 ( .A(KEYINPUT103), .B(n521), .Z(n522) );
  OR2_X1 U611 ( .A1(n522), .A2(G900), .ZN(n525) );
  INV_X1 U612 ( .A(n523), .ZN(n524) );
  NAND2_X1 U613 ( .A1(n525), .A2(n524), .ZN(n534) );
  NAND2_X1 U614 ( .A1(n695), .A2(n682), .ZN(n528) );
  XNOR2_X1 U615 ( .A(KEYINPUT105), .B(KEYINPUT30), .ZN(n527) );
  XNOR2_X1 U616 ( .A(n528), .B(n527), .ZN(n529) );
  BUF_X2 U617 ( .A(n531), .Z(n573) );
  NAND2_X1 U618 ( .A1(n564), .A2(n681), .ZN(n532) );
  INV_X1 U619 ( .A(n561), .ZN(n544) );
  AND2_X1 U620 ( .A1(n562), .A2(n544), .ZN(n664) );
  XNOR2_X1 U621 ( .A(n541), .B(G131), .ZN(G33) );
  AND2_X1 U622 ( .A1(n534), .A2(n691), .ZN(n535) );
  NAND2_X1 U623 ( .A1(n516), .A2(n535), .ZN(n550) );
  NOR2_X1 U624 ( .A1(n594), .A2(n550), .ZN(n537) );
  XNOR2_X1 U625 ( .A(KEYINPUT106), .B(KEYINPUT28), .ZN(n536) );
  XNOR2_X1 U626 ( .A(n537), .B(n536), .ZN(n539) );
  NAND2_X1 U627 ( .A1(n539), .A2(n538), .ZN(n543) );
  NAND2_X1 U628 ( .A1(n665), .A2(KEYINPUT47), .ZN(n548) );
  INV_X1 U629 ( .A(KEYINPUT47), .ZN(n556) );
  OR2_X1 U630 ( .A1(n562), .A2(n544), .ZN(n671) );
  INV_X1 U631 ( .A(n671), .ZN(n659) );
  NOR2_X1 U632 ( .A1(n659), .A2(n664), .ZN(n686) );
  NOR2_X1 U633 ( .A1(n686), .A2(KEYINPUT81), .ZN(n545) );
  NAND2_X1 U634 ( .A1(n665), .A2(n545), .ZN(n546) );
  NAND2_X1 U635 ( .A1(n556), .A2(n546), .ZN(n547) );
  NAND2_X1 U636 ( .A1(n548), .A2(n547), .ZN(n555) );
  AND2_X1 U637 ( .A1(n590), .A2(n682), .ZN(n549) );
  AND2_X1 U638 ( .A1(n664), .A2(n549), .ZN(n552) );
  INV_X1 U639 ( .A(n550), .ZN(n551) );
  NAND2_X1 U640 ( .A1(n552), .A2(n551), .ZN(n571) );
  XNOR2_X1 U641 ( .A(n553), .B(KEYINPUT36), .ZN(n554) );
  NAND2_X1 U642 ( .A1(n554), .A2(n352), .ZN(n674) );
  AND2_X1 U643 ( .A1(n555), .A2(n674), .ZN(n560) );
  NAND2_X1 U644 ( .A1(n665), .A2(KEYINPUT81), .ZN(n557) );
  NAND2_X1 U645 ( .A1(n557), .A2(n556), .ZN(n558) );
  NAND2_X1 U646 ( .A1(n558), .A2(n686), .ZN(n559) );
  NAND2_X1 U647 ( .A1(n560), .A2(n559), .ZN(n565) );
  NAND2_X1 U648 ( .A1(n562), .A2(n561), .ZN(n578) );
  NOR2_X1 U649 ( .A1(n573), .A2(n578), .ZN(n563) );
  AND2_X1 U650 ( .A1(n564), .A2(n563), .ZN(n663) );
  NOR2_X1 U651 ( .A1(n565), .A2(n663), .ZN(n566) );
  XNOR2_X1 U652 ( .A(n568), .B(n567), .ZN(n577) );
  NAND2_X1 U653 ( .A1(n569), .A2(n659), .ZN(n570) );
  XNOR2_X1 U654 ( .A(n570), .B(KEYINPUT110), .ZN(n748) );
  INV_X1 U655 ( .A(n748), .ZN(n575) );
  OR2_X1 U656 ( .A1(n571), .A2(n352), .ZN(n572) );
  XNOR2_X1 U657 ( .A(n572), .B(KEYINPUT43), .ZN(n574) );
  AND2_X1 U658 ( .A1(n574), .A2(n573), .ZN(n676) );
  NOR2_X1 U659 ( .A1(n575), .A2(n676), .ZN(n576) );
  NAND2_X1 U660 ( .A1(n577), .A2(n576), .ZN(n738) );
  INV_X1 U661 ( .A(n578), .ZN(n584) );
  NAND2_X1 U662 ( .A1(n580), .A2(n579), .ZN(n582) );
  NOR2_X1 U663 ( .A1(n695), .A2(n692), .ZN(n586) );
  INV_X1 U664 ( .A(n352), .ZN(n585) );
  NAND2_X1 U665 ( .A1(n352), .A2(n516), .ZN(n587) );
  XOR2_X1 U666 ( .A(KEYINPUT102), .B(n587), .Z(n588) );
  NOR2_X1 U667 ( .A1(KEYINPUT71), .A2(KEYINPUT44), .ZN(n591) );
  XNOR2_X1 U668 ( .A(n592), .B(n591), .ZN(n606) );
  NAND2_X1 U669 ( .A1(KEYINPUT71), .A2(KEYINPUT44), .ZN(n604) );
  XNOR2_X1 U670 ( .A(n686), .B(KEYINPUT81), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n593), .A2(n594), .ZN(n595) );
  NAND2_X1 U672 ( .A1(n695), .A2(n596), .ZN(n700) );
  XNOR2_X1 U673 ( .A(n597), .B(KEYINPUT31), .ZN(n670) );
  NAND2_X1 U674 ( .A1(n654), .A2(n670), .ZN(n598) );
  NAND2_X1 U675 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U676 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U677 ( .A(KEYINPUT101), .B(n602), .ZN(n603) );
  AND2_X1 U678 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U679 ( .A1(n606), .A2(n605), .ZN(n608) );
  INV_X1 U680 ( .A(KEYINPUT45), .ZN(n607) );
  XNOR2_X2 U681 ( .A(n608), .B(n607), .ZN(n730) );
  INV_X1 U682 ( .A(n614), .ZN(n609) );
  AND2_X1 U683 ( .A1(KEYINPUT82), .A2(n609), .ZN(n610) );
  INV_X1 U684 ( .A(KEYINPUT2), .ZN(n611) );
  OR2_X1 U685 ( .A1(n614), .A2(n611), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n613), .A2(n612), .ZN(n615) );
  NAND2_X1 U687 ( .A1(n717), .A2(G469), .ZN(n619) );
  XOR2_X1 U688 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n616) );
  XNOR2_X1 U689 ( .A(n617), .B(n616), .ZN(n618) );
  XNOR2_X1 U690 ( .A(n619), .B(n618), .ZN(n621) );
  INV_X1 U691 ( .A(G952), .ZN(n620) );
  NOR2_X1 U692 ( .A1(n621), .A2(n722), .ZN(G54) );
  NAND2_X1 U693 ( .A1(n717), .A2(G217), .ZN(n624) );
  XOR2_X1 U694 ( .A(KEYINPUT125), .B(n622), .Z(n623) );
  XNOR2_X1 U695 ( .A(n624), .B(n623), .ZN(n625) );
  NOR2_X1 U696 ( .A1(n625), .A2(n722), .ZN(G66) );
  INV_X1 U697 ( .A(n626), .ZN(n680) );
  INV_X1 U698 ( .A(G210), .ZN(n627) );
  NOR2_X1 U699 ( .A1(n680), .A2(n627), .ZN(n628) );
  NAND2_X1 U700 ( .A1(n629), .A2(n628), .ZN(n633) );
  XNOR2_X1 U701 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n630) );
  XNOR2_X1 U702 ( .A(n631), .B(n630), .ZN(n632) );
  XNOR2_X1 U703 ( .A(n633), .B(n632), .ZN(n634) );
  NOR2_X1 U704 ( .A1(n634), .A2(n722), .ZN(n635) );
  XNOR2_X1 U705 ( .A(n635), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U706 ( .A1(n717), .A2(G475), .ZN(n640) );
  XNOR2_X1 U707 ( .A(KEYINPUT64), .B(KEYINPUT123), .ZN(n636) );
  XNOR2_X1 U708 ( .A(n636), .B(KEYINPUT59), .ZN(n637) );
  XNOR2_X1 U709 ( .A(n638), .B(n637), .ZN(n639) );
  XNOR2_X1 U710 ( .A(n640), .B(n639), .ZN(n641) );
  XNOR2_X1 U711 ( .A(n642), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U712 ( .A1(n717), .A2(G472), .ZN(n647) );
  XNOR2_X1 U713 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n643) );
  XOR2_X1 U714 ( .A(n643), .B(KEYINPUT62), .Z(n644) );
  XNOR2_X1 U715 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U716 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U717 ( .A(KEYINPUT84), .B(KEYINPUT63), .ZN(n649) );
  XNOR2_X1 U718 ( .A(n649), .B(KEYINPUT83), .ZN(n650) );
  XNOR2_X1 U719 ( .A(n651), .B(n650), .ZN(G57) );
  INV_X1 U720 ( .A(n664), .ZN(n668) );
  NOR2_X1 U721 ( .A1(n668), .A2(n654), .ZN(n653) );
  XNOR2_X1 U722 ( .A(G104), .B(KEYINPUT113), .ZN(n652) );
  XNOR2_X1 U723 ( .A(n653), .B(n652), .ZN(G6) );
  NOR2_X1 U724 ( .A1(n671), .A2(n654), .ZN(n656) );
  XNOR2_X1 U725 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n655) );
  XNOR2_X1 U726 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U727 ( .A(G107), .B(n657), .ZN(G9) );
  XOR2_X1 U728 ( .A(G110), .B(n658), .Z(G12) );
  XOR2_X1 U729 ( .A(KEYINPUT114), .B(KEYINPUT29), .Z(n661) );
  NAND2_X1 U730 ( .A1(n665), .A2(n659), .ZN(n660) );
  XNOR2_X1 U731 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U732 ( .A(G128), .B(n662), .ZN(G30) );
  XOR2_X1 U733 ( .A(G143), .B(n663), .Z(G45) );
  XOR2_X1 U734 ( .A(G146), .B(KEYINPUT115), .Z(n667) );
  NAND2_X1 U735 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U736 ( .A(n667), .B(n666), .ZN(G48) );
  NOR2_X1 U737 ( .A1(n668), .A2(n670), .ZN(n669) );
  XOR2_X1 U738 ( .A(G113), .B(n669), .Z(G15) );
  NOR2_X1 U739 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U740 ( .A(G116), .B(n672), .Z(G18) );
  XOR2_X1 U741 ( .A(KEYINPUT37), .B(KEYINPUT116), .Z(n673) );
  XNOR2_X1 U742 ( .A(n674), .B(n673), .ZN(n675) );
  XNOR2_X1 U743 ( .A(G125), .B(n675), .ZN(G27) );
  XNOR2_X1 U744 ( .A(G140), .B(n676), .ZN(n677) );
  XNOR2_X1 U745 ( .A(n677), .B(KEYINPUT117), .ZN(G42) );
  NOR2_X1 U746 ( .A1(n678), .A2(KEYINPUT2), .ZN(n679) );
  NOR2_X1 U747 ( .A1(n680), .A2(n679), .ZN(n716) );
  NOR2_X1 U748 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U749 ( .A1(n684), .A2(n683), .ZN(n688) );
  NOR2_X1 U750 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U751 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U752 ( .A1(n709), .A2(n689), .ZN(n705) );
  NOR2_X1 U753 ( .A1(n352), .A2(n579), .ZN(n690) );
  XOR2_X1 U754 ( .A(KEYINPUT50), .B(n690), .Z(n698) );
  NOR2_X1 U755 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U756 ( .A(KEYINPUT49), .B(n693), .Z(n694) );
  NOR2_X1 U757 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U758 ( .A(KEYINPUT118), .B(n696), .ZN(n697) );
  NAND2_X1 U759 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U760 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U761 ( .A(KEYINPUT51), .B(n701), .ZN(n702) );
  NOR2_X1 U762 ( .A1(n710), .A2(n702), .ZN(n703) );
  XOR2_X1 U763 ( .A(KEYINPUT119), .B(n703), .Z(n704) );
  NOR2_X1 U764 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U765 ( .A(n706), .B(KEYINPUT52), .ZN(n707) );
  NOR2_X1 U766 ( .A1(n708), .A2(n707), .ZN(n713) );
  NOR2_X1 U767 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U768 ( .A(n711), .B(KEYINPUT120), .ZN(n712) );
  NOR2_X1 U769 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U770 ( .A(KEYINPUT121), .B(n714), .ZN(n715) );
  NAND2_X1 U771 ( .A1(n717), .A2(G478), .ZN(n720) );
  XNOR2_X1 U772 ( .A(n718), .B(KEYINPUT124), .ZN(n719) );
  XNOR2_X1 U773 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U774 ( .A1(n722), .A2(n721), .ZN(G63) );
  XNOR2_X1 U775 ( .A(n724), .B(n723), .ZN(n726) );
  NAND2_X1 U776 ( .A1(n726), .A2(n725), .ZN(n735) );
  NAND2_X1 U777 ( .A1(G224), .A2(G953), .ZN(n727) );
  XNOR2_X1 U778 ( .A(n727), .B(KEYINPUT126), .ZN(n728) );
  XNOR2_X1 U779 ( .A(KEYINPUT61), .B(n728), .ZN(n729) );
  NAND2_X1 U780 ( .A1(n729), .A2(G898), .ZN(n733) );
  NOR2_X1 U781 ( .A1(G953), .A2(n730), .ZN(n731) );
  XNOR2_X1 U782 ( .A(KEYINPUT127), .B(n731), .ZN(n732) );
  NAND2_X1 U783 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U784 ( .A(n735), .B(n734), .Z(G69) );
  XNOR2_X1 U785 ( .A(n737), .B(n736), .ZN(n741) );
  XNOR2_X1 U786 ( .A(n738), .B(n741), .ZN(n740) );
  NAND2_X1 U787 ( .A1(n740), .A2(n739), .ZN(n745) );
  XNOR2_X1 U788 ( .A(n741), .B(G227), .ZN(n742) );
  NAND2_X1 U789 ( .A1(n742), .A2(G900), .ZN(n743) );
  NAND2_X1 U790 ( .A1(n743), .A2(G953), .ZN(n744) );
  NAND2_X1 U791 ( .A1(n745), .A2(n744), .ZN(G72) );
  XOR2_X1 U792 ( .A(n746), .B(G122), .Z(G24) );
  XNOR2_X1 U793 ( .A(G119), .B(n747), .ZN(G21) );
  XNOR2_X1 U794 ( .A(G134), .B(n748), .ZN(G36) );
endmodule

