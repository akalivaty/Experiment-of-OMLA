

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U553 ( .A1(n539), .A2(n538), .ZN(G164) );
  AND2_X1 U554 ( .A1(n532), .A2(n531), .ZN(G160) );
  NAND2_X1 U555 ( .A1(n985), .A2(n802), .ZN(n521) );
  NOR2_X1 U556 ( .A1(n729), .A2(n947), .ZN(n687) );
  NOR2_X1 U557 ( .A1(n692), .A2(n967), .ZN(n693) );
  XNOR2_X1 U558 ( .A(n693), .B(KEYINPUT64), .ZN(n695) );
  INV_X1 U559 ( .A(KEYINPUT102), .ZN(n709) );
  XNOR2_X1 U560 ( .A(n710), .B(n709), .ZN(n714) );
  NAND2_X1 U561 ( .A1(n767), .A2(n685), .ZN(n729) );
  NOR2_X1 U562 ( .A1(n789), .A2(n521), .ZN(n790) );
  NOR2_X1 U563 ( .A1(G651), .A2(n635), .ZN(n651) );
  AND2_X1 U564 ( .A1(n822), .A2(n821), .ZN(n824) );
  NOR2_X1 U565 ( .A1(n550), .A2(n549), .ZN(G171) );
  INV_X1 U566 ( .A(G2105), .ZN(n526) );
  INV_X1 U567 ( .A(G2104), .ZN(n522) );
  NOR2_X1 U568 ( .A1(n526), .A2(n522), .ZN(n874) );
  NAND2_X1 U569 ( .A1(n874), .A2(G113), .ZN(n525) );
  NOR2_X2 U570 ( .A1(G2105), .A2(n522), .ZN(n869) );
  NAND2_X1 U571 ( .A1(G101), .A2(n869), .ZN(n523) );
  XOR2_X1 U572 ( .A(KEYINPUT23), .B(n523), .Z(n524) );
  AND2_X1 U573 ( .A1(n525), .A2(n524), .ZN(n532) );
  NOR2_X1 U574 ( .A1(G2104), .A2(n526), .ZN(n877) );
  NAND2_X1 U575 ( .A1(G125), .A2(n877), .ZN(n530) );
  XNOR2_X1 U576 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n528) );
  NOR2_X1 U577 ( .A1(G2105), .A2(G2104), .ZN(n527) );
  XNOR2_X2 U578 ( .A(n528), .B(n527), .ZN(n870) );
  NAND2_X1 U579 ( .A1(G137), .A2(n870), .ZN(n529) );
  AND2_X1 U580 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U581 ( .A1(G138), .A2(n870), .ZN(n533) );
  XOR2_X1 U582 ( .A(n533), .B(KEYINPUT90), .Z(n539) );
  NAND2_X1 U583 ( .A1(n877), .A2(G126), .ZN(n537) );
  NAND2_X1 U584 ( .A1(G114), .A2(n874), .ZN(n535) );
  NAND2_X1 U585 ( .A1(G102), .A2(n869), .ZN(n534) );
  AND2_X1 U586 ( .A1(n535), .A2(n534), .ZN(n536) );
  NAND2_X1 U587 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U588 ( .A(KEYINPUT9), .B(KEYINPUT69), .ZN(n543) );
  XOR2_X1 U589 ( .A(KEYINPUT0), .B(G543), .Z(n635) );
  INV_X1 U590 ( .A(G651), .ZN(n544) );
  NOR2_X1 U591 ( .A1(n635), .A2(n544), .ZN(n646) );
  NAND2_X1 U592 ( .A1(G77), .A2(n646), .ZN(n541) );
  NOR2_X1 U593 ( .A1(G651), .A2(G543), .ZN(n647) );
  NAND2_X1 U594 ( .A1(G90), .A2(n647), .ZN(n540) );
  NAND2_X1 U595 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U596 ( .A(n543), .B(n542), .ZN(n550) );
  NOR2_X1 U597 ( .A1(G543), .A2(n544), .ZN(n545) );
  XOR2_X1 U598 ( .A(KEYINPUT1), .B(n545), .Z(n650) );
  NAND2_X1 U599 ( .A1(n650), .A2(G64), .ZN(n546) );
  XNOR2_X1 U600 ( .A(n546), .B(KEYINPUT68), .ZN(n548) );
  NAND2_X1 U601 ( .A1(G52), .A2(n651), .ZN(n547) );
  NAND2_X1 U602 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U603 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U604 ( .A(G57), .ZN(G237) );
  INV_X1 U605 ( .A(G120), .ZN(G236) );
  INV_X1 U606 ( .A(G69), .ZN(G235) );
  NAND2_X1 U607 ( .A1(n647), .A2(G89), .ZN(n551) );
  XNOR2_X1 U608 ( .A(n551), .B(KEYINPUT4), .ZN(n553) );
  NAND2_X1 U609 ( .A1(G76), .A2(n646), .ZN(n552) );
  NAND2_X1 U610 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U611 ( .A(n554), .B(KEYINPUT5), .ZN(n559) );
  NAND2_X1 U612 ( .A1(G63), .A2(n650), .ZN(n556) );
  NAND2_X1 U613 ( .A1(G51), .A2(n651), .ZN(n555) );
  NAND2_X1 U614 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U615 ( .A(KEYINPUT6), .B(n557), .Z(n558) );
  NAND2_X1 U616 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U617 ( .A(n560), .B(KEYINPUT7), .ZN(G168) );
  XNOR2_X1 U618 ( .A(G168), .B(KEYINPUT8), .ZN(n561) );
  XNOR2_X1 U619 ( .A(n561), .B(KEYINPUT77), .ZN(G286) );
  NAND2_X1 U620 ( .A1(G7), .A2(G661), .ZN(n562) );
  XNOR2_X1 U621 ( .A(n562), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U622 ( .A(G223), .B(KEYINPUT71), .ZN(n825) );
  NAND2_X1 U623 ( .A1(n825), .A2(G567), .ZN(n563) );
  XOR2_X1 U624 ( .A(KEYINPUT11), .B(n563), .Z(G234) );
  NAND2_X1 U625 ( .A1(n647), .A2(G81), .ZN(n564) );
  XNOR2_X1 U626 ( .A(n564), .B(KEYINPUT12), .ZN(n566) );
  NAND2_X1 U627 ( .A1(G68), .A2(n646), .ZN(n565) );
  NAND2_X1 U628 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U629 ( .A(KEYINPUT13), .B(n567), .ZN(n573) );
  NAND2_X1 U630 ( .A1(G56), .A2(n650), .ZN(n568) );
  XOR2_X1 U631 ( .A(KEYINPUT14), .B(n568), .Z(n571) );
  NAND2_X1 U632 ( .A1(n651), .A2(G43), .ZN(n569) );
  XOR2_X1 U633 ( .A(KEYINPUT72), .B(n569), .Z(n570) );
  NOR2_X1 U634 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U635 ( .A1(n573), .A2(n572), .ZN(n967) );
  INV_X1 U636 ( .A(G860), .ZN(n597) );
  OR2_X1 U637 ( .A1(n967), .A2(n597), .ZN(G153) );
  INV_X1 U638 ( .A(G868), .ZN(n667) );
  NOR2_X1 U639 ( .A1(n667), .A2(G171), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n574), .B(KEYINPUT73), .ZN(n586) );
  NAND2_X1 U641 ( .A1(G79), .A2(n646), .ZN(n576) );
  NAND2_X1 U642 ( .A1(G54), .A2(n651), .ZN(n575) );
  NAND2_X1 U643 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U644 ( .A(KEYINPUT74), .B(n577), .ZN(n581) );
  NAND2_X1 U645 ( .A1(G92), .A2(n647), .ZN(n579) );
  NAND2_X1 U646 ( .A1(G66), .A2(n650), .ZN(n578) );
  NAND2_X1 U647 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U648 ( .A1(n581), .A2(n580), .ZN(n583) );
  XNOR2_X1 U649 ( .A(KEYINPUT75), .B(KEYINPUT76), .ZN(n582) );
  XNOR2_X1 U650 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U651 ( .A(KEYINPUT15), .B(n584), .ZN(n970) );
  OR2_X1 U652 ( .A1(G868), .A2(n970), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n586), .A2(n585), .ZN(G284) );
  NAND2_X1 U654 ( .A1(G78), .A2(n646), .ZN(n588) );
  NAND2_X1 U655 ( .A1(G91), .A2(n647), .ZN(n587) );
  NAND2_X1 U656 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U657 ( .A1(n651), .A2(G53), .ZN(n589) );
  XOR2_X1 U658 ( .A(KEYINPUT70), .B(n589), .Z(n590) );
  NOR2_X1 U659 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U660 ( .A1(n650), .A2(G65), .ZN(n592) );
  NAND2_X1 U661 ( .A1(n593), .A2(n592), .ZN(G299) );
  NOR2_X1 U662 ( .A1(G286), .A2(n667), .ZN(n594) );
  XNOR2_X1 U663 ( .A(n594), .B(KEYINPUT78), .ZN(n596) );
  NOR2_X1 U664 ( .A1(G299), .A2(G868), .ZN(n595) );
  NOR2_X1 U665 ( .A1(n596), .A2(n595), .ZN(G297) );
  NAND2_X1 U666 ( .A1(n597), .A2(G559), .ZN(n598) );
  NAND2_X1 U667 ( .A1(n598), .A2(n970), .ZN(n599) );
  XNOR2_X1 U668 ( .A(n599), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U669 ( .A1(G868), .A2(n967), .ZN(n600) );
  XOR2_X1 U670 ( .A(KEYINPUT79), .B(n600), .Z(n603) );
  NAND2_X1 U671 ( .A1(G868), .A2(n970), .ZN(n601) );
  NOR2_X1 U672 ( .A1(G559), .A2(n601), .ZN(n602) );
  NOR2_X1 U673 ( .A1(n603), .A2(n602), .ZN(G282) );
  NAND2_X1 U674 ( .A1(G111), .A2(n874), .ZN(n605) );
  NAND2_X1 U675 ( .A1(G99), .A2(n869), .ZN(n604) );
  NAND2_X1 U676 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U677 ( .A(KEYINPUT80), .B(n606), .ZN(n609) );
  NAND2_X1 U678 ( .A1(n877), .A2(G123), .ZN(n607) );
  XOR2_X1 U679 ( .A(KEYINPUT18), .B(n607), .Z(n608) );
  NOR2_X1 U680 ( .A1(n609), .A2(n608), .ZN(n611) );
  NAND2_X1 U681 ( .A1(n870), .A2(G135), .ZN(n610) );
  NAND2_X1 U682 ( .A1(n611), .A2(n610), .ZN(n921) );
  XOR2_X1 U683 ( .A(n921), .B(G2096), .Z(n613) );
  XNOR2_X1 U684 ( .A(G2100), .B(KEYINPUT81), .ZN(n612) );
  NAND2_X1 U685 ( .A1(n613), .A2(n612), .ZN(G156) );
  NAND2_X1 U686 ( .A1(G559), .A2(n970), .ZN(n665) );
  XNOR2_X1 U687 ( .A(n967), .B(n665), .ZN(n614) );
  NOR2_X1 U688 ( .A1(n614), .A2(G860), .ZN(n622) );
  NAND2_X1 U689 ( .A1(G93), .A2(n647), .ZN(n615) );
  XNOR2_X1 U690 ( .A(n615), .B(KEYINPUT82), .ZN(n617) );
  NAND2_X1 U691 ( .A1(n646), .A2(G80), .ZN(n616) );
  NAND2_X1 U692 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U693 ( .A1(G67), .A2(n650), .ZN(n619) );
  NAND2_X1 U694 ( .A1(G55), .A2(n651), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n619), .A2(n618), .ZN(n620) );
  OR2_X1 U696 ( .A1(n621), .A2(n620), .ZN(n668) );
  XOR2_X1 U697 ( .A(n622), .B(n668), .Z(G145) );
  XOR2_X1 U698 ( .A(KEYINPUT84), .B(KEYINPUT2), .Z(n624) );
  NAND2_X1 U699 ( .A1(G73), .A2(n646), .ZN(n623) );
  XNOR2_X1 U700 ( .A(n624), .B(n623), .ZN(n629) );
  NAND2_X1 U701 ( .A1(G86), .A2(n647), .ZN(n626) );
  NAND2_X1 U702 ( .A1(G61), .A2(n650), .ZN(n625) );
  NAND2_X1 U703 ( .A1(n626), .A2(n625), .ZN(n627) );
  XOR2_X1 U704 ( .A(KEYINPUT83), .B(n627), .Z(n628) );
  NOR2_X1 U705 ( .A1(n629), .A2(n628), .ZN(n631) );
  NAND2_X1 U706 ( .A1(n651), .A2(G48), .ZN(n630) );
  NAND2_X1 U707 ( .A1(n631), .A2(n630), .ZN(G305) );
  NAND2_X1 U708 ( .A1(G49), .A2(n651), .ZN(n633) );
  NAND2_X1 U709 ( .A1(G74), .A2(G651), .ZN(n632) );
  NAND2_X1 U710 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U711 ( .A1(n650), .A2(n634), .ZN(n637) );
  NAND2_X1 U712 ( .A1(n635), .A2(G87), .ZN(n636) );
  NAND2_X1 U713 ( .A1(n637), .A2(n636), .ZN(G288) );
  NAND2_X1 U714 ( .A1(n647), .A2(G85), .ZN(n644) );
  NAND2_X1 U715 ( .A1(G60), .A2(n650), .ZN(n639) );
  NAND2_X1 U716 ( .A1(G47), .A2(n651), .ZN(n638) );
  NAND2_X1 U717 ( .A1(n639), .A2(n638), .ZN(n642) );
  NAND2_X1 U718 ( .A1(G72), .A2(n646), .ZN(n640) );
  XOR2_X1 U719 ( .A(KEYINPUT66), .B(n640), .Z(n641) );
  NOR2_X1 U720 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U721 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U722 ( .A(KEYINPUT67), .B(n645), .Z(G290) );
  NAND2_X1 U723 ( .A1(G75), .A2(n646), .ZN(n649) );
  NAND2_X1 U724 ( .A1(G88), .A2(n647), .ZN(n648) );
  NAND2_X1 U725 ( .A1(n649), .A2(n648), .ZN(n655) );
  NAND2_X1 U726 ( .A1(G62), .A2(n650), .ZN(n653) );
  NAND2_X1 U727 ( .A1(G50), .A2(n651), .ZN(n652) );
  NAND2_X1 U728 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U729 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U730 ( .A(KEYINPUT85), .B(n656), .Z(G166) );
  XOR2_X1 U731 ( .A(n967), .B(G305), .Z(n660) );
  XNOR2_X1 U732 ( .A(KEYINPUT86), .B(KEYINPUT87), .ZN(n658) );
  XNOR2_X1 U733 ( .A(G288), .B(KEYINPUT19), .ZN(n657) );
  XNOR2_X1 U734 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U735 ( .A(n660), .B(n659), .ZN(n662) );
  XNOR2_X1 U736 ( .A(G290), .B(G166), .ZN(n661) );
  XNOR2_X1 U737 ( .A(n662), .B(n661), .ZN(n663) );
  XOR2_X1 U738 ( .A(n668), .B(n663), .Z(n664) );
  XNOR2_X1 U739 ( .A(n664), .B(G299), .ZN(n894) );
  XOR2_X1 U740 ( .A(n894), .B(n665), .Z(n666) );
  NOR2_X1 U741 ( .A1(n667), .A2(n666), .ZN(n670) );
  NOR2_X1 U742 ( .A1(G868), .A2(n668), .ZN(n669) );
  NOR2_X1 U743 ( .A1(n670), .A2(n669), .ZN(G295) );
  NAND2_X1 U744 ( .A1(G2078), .A2(G2084), .ZN(n671) );
  XOR2_X1 U745 ( .A(KEYINPUT20), .B(n671), .Z(n672) );
  NAND2_X1 U746 ( .A1(G2090), .A2(n672), .ZN(n673) );
  XNOR2_X1 U747 ( .A(KEYINPUT21), .B(n673), .ZN(n674) );
  NAND2_X1 U748 ( .A1(n674), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U749 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U750 ( .A1(G235), .A2(G236), .ZN(n675) );
  NAND2_X1 U751 ( .A1(G108), .A2(n675), .ZN(n676) );
  NOR2_X1 U752 ( .A1(n676), .A2(G237), .ZN(n677) );
  XNOR2_X1 U753 ( .A(n677), .B(KEYINPUT89), .ZN(n913) );
  NAND2_X1 U754 ( .A1(n913), .A2(G567), .ZN(n683) );
  NAND2_X1 U755 ( .A1(G132), .A2(G82), .ZN(n678) );
  XNOR2_X1 U756 ( .A(n678), .B(KEYINPUT22), .ZN(n679) );
  XNOR2_X1 U757 ( .A(n679), .B(KEYINPUT88), .ZN(n680) );
  NOR2_X1 U758 ( .A1(G218), .A2(n680), .ZN(n681) );
  NAND2_X1 U759 ( .A1(G96), .A2(n681), .ZN(n914) );
  NAND2_X1 U760 ( .A1(n914), .A2(G2106), .ZN(n682) );
  NAND2_X1 U761 ( .A1(n683), .A2(n682), .ZN(n829) );
  NAND2_X1 U762 ( .A1(G483), .A2(G661), .ZN(n684) );
  NOR2_X1 U763 ( .A1(n829), .A2(n684), .ZN(n828) );
  NAND2_X1 U764 ( .A1(n828), .A2(G36), .ZN(G176) );
  XNOR2_X1 U765 ( .A(KEYINPUT91), .B(G166), .ZN(G303) );
  NOR2_X1 U766 ( .A1(G164), .A2(G1384), .ZN(n767) );
  NAND2_X1 U767 ( .A1(G160), .A2(G40), .ZN(n768) );
  INV_X1 U768 ( .A(n768), .ZN(n685) );
  NAND2_X1 U769 ( .A1(G8), .A2(n729), .ZN(n798) );
  INV_X1 U770 ( .A(G1996), .ZN(n947) );
  XOR2_X1 U771 ( .A(KEYINPUT26), .B(KEYINPUT98), .Z(n686) );
  XNOR2_X1 U772 ( .A(n687), .B(n686), .ZN(n689) );
  NAND2_X1 U773 ( .A1(n729), .A2(G1341), .ZN(n688) );
  NAND2_X1 U774 ( .A1(n689), .A2(n688), .ZN(n691) );
  INV_X1 U775 ( .A(KEYINPUT99), .ZN(n690) );
  XNOR2_X1 U776 ( .A(n691), .B(n690), .ZN(n692) );
  NOR2_X1 U777 ( .A1(n970), .A2(n695), .ZN(n694) );
  XNOR2_X1 U778 ( .A(n694), .B(KEYINPUT101), .ZN(n702) );
  NAND2_X1 U779 ( .A1(n970), .A2(n695), .ZN(n700) );
  NAND2_X1 U780 ( .A1(n729), .A2(G1348), .ZN(n696) );
  XNOR2_X1 U781 ( .A(n696), .B(KEYINPUT100), .ZN(n698) );
  INV_X1 U782 ( .A(n729), .ZN(n717) );
  NAND2_X1 U783 ( .A1(n717), .A2(G2067), .ZN(n697) );
  NAND2_X1 U784 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U785 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U786 ( .A1(n702), .A2(n701), .ZN(n708) );
  INV_X1 U787 ( .A(G2072), .ZN(n930) );
  NOR2_X1 U788 ( .A1(n729), .A2(n930), .ZN(n704) );
  XOR2_X1 U789 ( .A(KEYINPUT97), .B(KEYINPUT27), .Z(n703) );
  XNOR2_X1 U790 ( .A(n704), .B(n703), .ZN(n706) );
  NAND2_X1 U791 ( .A1(n729), .A2(G1956), .ZN(n705) );
  NAND2_X1 U792 ( .A1(n706), .A2(n705), .ZN(n711) );
  OR2_X1 U793 ( .A1(G299), .A2(n711), .ZN(n707) );
  NAND2_X1 U794 ( .A1(n708), .A2(n707), .ZN(n710) );
  NAND2_X1 U795 ( .A1(G299), .A2(n711), .ZN(n712) );
  XOR2_X1 U796 ( .A(KEYINPUT28), .B(n712), .Z(n713) );
  NOR2_X1 U797 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U798 ( .A(n715), .B(KEYINPUT29), .ZN(n721) );
  INV_X1 U799 ( .A(G1961), .ZN(n1010) );
  NAND2_X1 U800 ( .A1(n729), .A2(n1010), .ZN(n719) );
  XNOR2_X1 U801 ( .A(G2078), .B(KEYINPUT25), .ZN(n716) );
  XNOR2_X1 U802 ( .A(n716), .B(KEYINPUT96), .ZN(n946) );
  NAND2_X1 U803 ( .A1(n717), .A2(n946), .ZN(n718) );
  NAND2_X1 U804 ( .A1(n719), .A2(n718), .ZN(n725) );
  NAND2_X1 U805 ( .A1(G171), .A2(n725), .ZN(n720) );
  NAND2_X1 U806 ( .A1(n721), .A2(n720), .ZN(n742) );
  NOR2_X1 U807 ( .A1(G1966), .A2(n798), .ZN(n744) );
  NOR2_X1 U808 ( .A1(G2084), .A2(n729), .ZN(n743) );
  NOR2_X1 U809 ( .A1(n744), .A2(n743), .ZN(n722) );
  NAND2_X1 U810 ( .A1(G8), .A2(n722), .ZN(n723) );
  XNOR2_X1 U811 ( .A(KEYINPUT30), .B(n723), .ZN(n724) );
  NOR2_X1 U812 ( .A1(G168), .A2(n724), .ZN(n727) );
  NOR2_X1 U813 ( .A1(G171), .A2(n725), .ZN(n726) );
  NOR2_X1 U814 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U815 ( .A(KEYINPUT31), .B(n728), .Z(n741) );
  INV_X1 U816 ( .A(G8), .ZN(n734) );
  NOR2_X1 U817 ( .A1(G1971), .A2(n798), .ZN(n731) );
  NOR2_X1 U818 ( .A1(G2090), .A2(n729), .ZN(n730) );
  NOR2_X1 U819 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U820 ( .A1(n732), .A2(G303), .ZN(n733) );
  OR2_X1 U821 ( .A1(n734), .A2(n733), .ZN(n736) );
  AND2_X1 U822 ( .A1(n741), .A2(n736), .ZN(n735) );
  NAND2_X1 U823 ( .A1(n742), .A2(n735), .ZN(n739) );
  INV_X1 U824 ( .A(n736), .ZN(n737) );
  OR2_X1 U825 ( .A1(n737), .A2(G286), .ZN(n738) );
  NAND2_X1 U826 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U827 ( .A(n740), .B(KEYINPUT32), .ZN(n749) );
  AND2_X1 U828 ( .A1(n742), .A2(n741), .ZN(n747) );
  AND2_X1 U829 ( .A1(G8), .A2(n743), .ZN(n745) );
  OR2_X1 U830 ( .A1(n745), .A2(n744), .ZN(n746) );
  OR2_X1 U831 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U832 ( .A1(n749), .A2(n748), .ZN(n794) );
  NOR2_X1 U833 ( .A1(G1976), .A2(G288), .ZN(n973) );
  NOR2_X1 U834 ( .A1(G1971), .A2(G303), .ZN(n750) );
  NOR2_X1 U835 ( .A1(n973), .A2(n750), .ZN(n751) );
  NAND2_X1 U836 ( .A1(n794), .A2(n751), .ZN(n752) );
  NAND2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n974) );
  NAND2_X1 U838 ( .A1(n752), .A2(n974), .ZN(n753) );
  NOR2_X1 U839 ( .A1(n798), .A2(n753), .ZN(n754) );
  NOR2_X1 U840 ( .A1(KEYINPUT33), .A2(n754), .ZN(n755) );
  INV_X1 U841 ( .A(n755), .ZN(n791) );
  NAND2_X1 U842 ( .A1(n973), .A2(KEYINPUT33), .ZN(n756) );
  NOR2_X1 U843 ( .A1(n756), .A2(n798), .ZN(n789) );
  XOR2_X1 U844 ( .A(G1981), .B(G305), .Z(n985) );
  NAND2_X1 U845 ( .A1(n870), .A2(G140), .ZN(n757) );
  XOR2_X1 U846 ( .A(KEYINPUT93), .B(n757), .Z(n759) );
  NAND2_X1 U847 ( .A1(n869), .A2(G104), .ZN(n758) );
  NAND2_X1 U848 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U849 ( .A(KEYINPUT34), .B(n760), .ZN(n765) );
  NAND2_X1 U850 ( .A1(G116), .A2(n874), .ZN(n762) );
  NAND2_X1 U851 ( .A1(G128), .A2(n877), .ZN(n761) );
  NAND2_X1 U852 ( .A1(n762), .A2(n761), .ZN(n763) );
  XOR2_X1 U853 ( .A(KEYINPUT35), .B(n763), .Z(n764) );
  NOR2_X1 U854 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U855 ( .A(KEYINPUT36), .B(n766), .ZN(n891) );
  XNOR2_X1 U856 ( .A(G2067), .B(KEYINPUT37), .ZN(n803) );
  NOR2_X1 U857 ( .A1(n891), .A2(n803), .ZN(n927) );
  NOR2_X1 U858 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U859 ( .A(n769), .B(KEYINPUT92), .ZN(n818) );
  NAND2_X1 U860 ( .A1(n927), .A2(n818), .ZN(n811) );
  INV_X1 U861 ( .A(n818), .ZN(n787) );
  NAND2_X1 U862 ( .A1(G117), .A2(n874), .ZN(n771) );
  NAND2_X1 U863 ( .A1(G129), .A2(n877), .ZN(n770) );
  NAND2_X1 U864 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U865 ( .A(KEYINPUT94), .B(n772), .ZN(n775) );
  NAND2_X1 U866 ( .A1(n869), .A2(G105), .ZN(n773) );
  XOR2_X1 U867 ( .A(KEYINPUT38), .B(n773), .Z(n774) );
  NOR2_X1 U868 ( .A1(n775), .A2(n774), .ZN(n777) );
  NAND2_X1 U869 ( .A1(n870), .A2(G141), .ZN(n776) );
  NAND2_X1 U870 ( .A1(n777), .A2(n776), .ZN(n868) );
  NAND2_X1 U871 ( .A1(n868), .A2(G1996), .ZN(n785) );
  NAND2_X1 U872 ( .A1(G107), .A2(n874), .ZN(n779) );
  NAND2_X1 U873 ( .A1(G95), .A2(n869), .ZN(n778) );
  NAND2_X1 U874 ( .A1(n779), .A2(n778), .ZN(n783) );
  NAND2_X1 U875 ( .A1(G119), .A2(n877), .ZN(n781) );
  NAND2_X1 U876 ( .A1(G131), .A2(n870), .ZN(n780) );
  NAND2_X1 U877 ( .A1(n781), .A2(n780), .ZN(n782) );
  OR2_X1 U878 ( .A1(n783), .A2(n782), .ZN(n888) );
  NAND2_X1 U879 ( .A1(G1991), .A2(n888), .ZN(n784) );
  NAND2_X1 U880 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U881 ( .A(n786), .B(KEYINPUT95), .ZN(n920) );
  NOR2_X1 U882 ( .A1(n787), .A2(n920), .ZN(n807) );
  INV_X1 U883 ( .A(n807), .ZN(n788) );
  AND2_X1 U884 ( .A1(n811), .A2(n788), .ZN(n802) );
  NAND2_X1 U885 ( .A1(n791), .A2(n790), .ZN(n817) );
  NOR2_X1 U886 ( .A1(G2090), .A2(G303), .ZN(n792) );
  NAND2_X1 U887 ( .A1(G8), .A2(n792), .ZN(n793) );
  NAND2_X1 U888 ( .A1(n794), .A2(n793), .ZN(n795) );
  NAND2_X1 U889 ( .A1(n795), .A2(n798), .ZN(n800) );
  NOR2_X1 U890 ( .A1(G1981), .A2(G305), .ZN(n796) );
  XOR2_X1 U891 ( .A(n796), .B(KEYINPUT24), .Z(n797) );
  OR2_X1 U892 ( .A1(n798), .A2(n797), .ZN(n799) );
  NAND2_X1 U893 ( .A1(n800), .A2(n799), .ZN(n801) );
  AND2_X1 U894 ( .A1(n802), .A2(n801), .ZN(n815) );
  NAND2_X1 U895 ( .A1(n891), .A2(n803), .ZN(n936) );
  NOR2_X1 U896 ( .A1(G1996), .A2(n868), .ZN(n917) );
  NOR2_X1 U897 ( .A1(G1991), .A2(n888), .ZN(n924) );
  NOR2_X1 U898 ( .A1(G1986), .A2(G290), .ZN(n804) );
  NOR2_X1 U899 ( .A1(n924), .A2(n804), .ZN(n805) );
  XOR2_X1 U900 ( .A(KEYINPUT103), .B(n805), .Z(n806) );
  NOR2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n808) );
  NOR2_X1 U902 ( .A1(n917), .A2(n808), .ZN(n809) );
  XNOR2_X1 U903 ( .A(KEYINPUT104), .B(n809), .ZN(n810) );
  XNOR2_X1 U904 ( .A(n810), .B(KEYINPUT39), .ZN(n812) );
  NAND2_X1 U905 ( .A1(n812), .A2(n811), .ZN(n813) );
  NAND2_X1 U906 ( .A1(n936), .A2(n813), .ZN(n814) );
  AND2_X1 U907 ( .A1(n814), .A2(n818), .ZN(n820) );
  NOR2_X1 U908 ( .A1(n815), .A2(n820), .ZN(n816) );
  NAND2_X1 U909 ( .A1(n817), .A2(n816), .ZN(n822) );
  XNOR2_X1 U910 ( .A(G1986), .B(G290), .ZN(n969) );
  NAND2_X1 U911 ( .A1(n969), .A2(n818), .ZN(n819) );
  OR2_X1 U912 ( .A1(n820), .A2(n819), .ZN(n821) );
  XOR2_X1 U913 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n823) );
  XNOR2_X1 U914 ( .A(n824), .B(n823), .ZN(G329) );
  NAND2_X1 U915 ( .A1(G2106), .A2(n825), .ZN(G217) );
  AND2_X1 U916 ( .A1(G15), .A2(G2), .ZN(n826) );
  NAND2_X1 U917 ( .A1(G661), .A2(n826), .ZN(G259) );
  NAND2_X1 U918 ( .A1(G3), .A2(G1), .ZN(n827) );
  NAND2_X1 U919 ( .A1(n828), .A2(n827), .ZN(G188) );
  INV_X1 U920 ( .A(n829), .ZN(G319) );
  XOR2_X1 U921 ( .A(KEYINPUT107), .B(G1976), .Z(n831) );
  XNOR2_X1 U922 ( .A(G1986), .B(G1956), .ZN(n830) );
  XNOR2_X1 U923 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U924 ( .A(n832), .B(KEYINPUT41), .Z(n834) );
  XNOR2_X1 U925 ( .A(G1996), .B(G1991), .ZN(n833) );
  XNOR2_X1 U926 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U927 ( .A(G1981), .B(G1971), .Z(n836) );
  XNOR2_X1 U928 ( .A(G1966), .B(G1961), .ZN(n835) );
  XNOR2_X1 U929 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U930 ( .A(n838), .B(n837), .Z(n840) );
  XNOR2_X1 U931 ( .A(G2474), .B(KEYINPUT108), .ZN(n839) );
  XNOR2_X1 U932 ( .A(n840), .B(n839), .ZN(G229) );
  XOR2_X1 U933 ( .A(G2100), .B(G2096), .Z(n842) );
  XNOR2_X1 U934 ( .A(KEYINPUT42), .B(G2678), .ZN(n841) );
  XNOR2_X1 U935 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U936 ( .A(KEYINPUT43), .B(G2090), .Z(n844) );
  XNOR2_X1 U937 ( .A(G2067), .B(G2072), .ZN(n843) );
  XNOR2_X1 U938 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U939 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U940 ( .A(G2078), .B(G2084), .ZN(n847) );
  XNOR2_X1 U941 ( .A(n848), .B(n847), .ZN(G227) );
  NAND2_X1 U942 ( .A1(G136), .A2(n870), .ZN(n855) );
  NAND2_X1 U943 ( .A1(G112), .A2(n874), .ZN(n850) );
  NAND2_X1 U944 ( .A1(G100), .A2(n869), .ZN(n849) );
  NAND2_X1 U945 ( .A1(n850), .A2(n849), .ZN(n853) );
  NAND2_X1 U946 ( .A1(n877), .A2(G124), .ZN(n851) );
  XOR2_X1 U947 ( .A(KEYINPUT44), .B(n851), .Z(n852) );
  NOR2_X1 U948 ( .A1(n853), .A2(n852), .ZN(n854) );
  NAND2_X1 U949 ( .A1(n855), .A2(n854), .ZN(n856) );
  XNOR2_X1 U950 ( .A(n856), .B(KEYINPUT109), .ZN(G162) );
  XNOR2_X1 U951 ( .A(KEYINPUT113), .B(KEYINPUT47), .ZN(n861) );
  NAND2_X1 U952 ( .A1(n874), .A2(G115), .ZN(n857) );
  XNOR2_X1 U953 ( .A(n857), .B(KEYINPUT112), .ZN(n859) );
  NAND2_X1 U954 ( .A1(G127), .A2(n877), .ZN(n858) );
  NAND2_X1 U955 ( .A1(n859), .A2(n858), .ZN(n860) );
  XNOR2_X1 U956 ( .A(n861), .B(n860), .ZN(n866) );
  NAND2_X1 U957 ( .A1(G103), .A2(n869), .ZN(n863) );
  NAND2_X1 U958 ( .A1(G139), .A2(n870), .ZN(n862) );
  NAND2_X1 U959 ( .A1(n863), .A2(n862), .ZN(n864) );
  XOR2_X1 U960 ( .A(KEYINPUT111), .B(n864), .Z(n865) );
  NOR2_X1 U961 ( .A1(n866), .A2(n865), .ZN(n929) );
  XOR2_X1 U962 ( .A(G160), .B(n929), .Z(n867) );
  XNOR2_X1 U963 ( .A(n868), .B(n867), .ZN(n884) );
  NAND2_X1 U964 ( .A1(G106), .A2(n869), .ZN(n872) );
  NAND2_X1 U965 ( .A1(G142), .A2(n870), .ZN(n871) );
  NAND2_X1 U966 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U967 ( .A(n873), .B(KEYINPUT45), .ZN(n876) );
  NAND2_X1 U968 ( .A1(G118), .A2(n874), .ZN(n875) );
  NAND2_X1 U969 ( .A1(n876), .A2(n875), .ZN(n880) );
  NAND2_X1 U970 ( .A1(n877), .A2(G130), .ZN(n878) );
  XOR2_X1 U971 ( .A(KEYINPUT110), .B(n878), .Z(n879) );
  NOR2_X1 U972 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U973 ( .A(G164), .B(n881), .Z(n882) );
  XNOR2_X1 U974 ( .A(n921), .B(n882), .ZN(n883) );
  XNOR2_X1 U975 ( .A(n884), .B(n883), .ZN(n890) );
  XOR2_X1 U976 ( .A(KEYINPUT114), .B(KEYINPUT48), .Z(n886) );
  XNOR2_X1 U977 ( .A(G162), .B(KEYINPUT46), .ZN(n885) );
  XNOR2_X1 U978 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U979 ( .A(n888), .B(n887), .ZN(n889) );
  XNOR2_X1 U980 ( .A(n890), .B(n889), .ZN(n892) );
  XNOR2_X1 U981 ( .A(n892), .B(n891), .ZN(n893) );
  NOR2_X1 U982 ( .A1(G37), .A2(n893), .ZN(G395) );
  XNOR2_X1 U983 ( .A(G286), .B(n970), .ZN(n895) );
  XNOR2_X1 U984 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U985 ( .A(n896), .B(G171), .ZN(n897) );
  NOR2_X1 U986 ( .A1(G37), .A2(n897), .ZN(G397) );
  XOR2_X1 U987 ( .A(G2438), .B(G2435), .Z(n899) );
  XNOR2_X1 U988 ( .A(G2443), .B(G2430), .ZN(n898) );
  XNOR2_X1 U989 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U990 ( .A(n900), .B(G2454), .Z(n902) );
  XNOR2_X1 U991 ( .A(G1348), .B(G1341), .ZN(n901) );
  XNOR2_X1 U992 ( .A(n902), .B(n901), .ZN(n906) );
  XOR2_X1 U993 ( .A(G2451), .B(G2427), .Z(n904) );
  XNOR2_X1 U994 ( .A(KEYINPUT106), .B(G2446), .ZN(n903) );
  XNOR2_X1 U995 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U996 ( .A(n906), .B(n905), .Z(n907) );
  NAND2_X1 U997 ( .A1(G14), .A2(n907), .ZN(n915) );
  NAND2_X1 U998 ( .A1(G319), .A2(n915), .ZN(n910) );
  NOR2_X1 U999 ( .A1(G229), .A2(G227), .ZN(n908) );
  XNOR2_X1 U1000 ( .A(KEYINPUT49), .B(n908), .ZN(n909) );
  NOR2_X1 U1001 ( .A1(n910), .A2(n909), .ZN(n912) );
  NOR2_X1 U1002 ( .A1(G395), .A2(G397), .ZN(n911) );
  NAND2_X1 U1003 ( .A1(n912), .A2(n911), .ZN(G225) );
  XNOR2_X1 U1004 ( .A(KEYINPUT115), .B(G225), .ZN(G308) );
  XOR2_X1 U1005 ( .A(G108), .B(KEYINPUT116), .Z(G238) );
  INV_X1 U1007 ( .A(G132), .ZN(G219) );
  INV_X1 U1008 ( .A(G82), .ZN(G220) );
  NOR2_X1 U1009 ( .A1(n914), .A2(n913), .ZN(G325) );
  INV_X1 U1010 ( .A(G325), .ZN(G261) );
  INV_X1 U1011 ( .A(G171), .ZN(G301) );
  INV_X1 U1012 ( .A(G96), .ZN(G221) );
  INV_X1 U1013 ( .A(n915), .ZN(G401) );
  XOR2_X1 U1014 ( .A(G2090), .B(G162), .Z(n916) );
  NOR2_X1 U1015 ( .A1(n917), .A2(n916), .ZN(n918) );
  XOR2_X1 U1016 ( .A(KEYINPUT51), .B(n918), .Z(n919) );
  NAND2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(n939) );
  XNOR2_X1 U1018 ( .A(G160), .B(G2084), .ZN(n922) );
  NAND2_X1 U1019 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1021 ( .A(n925), .B(KEYINPUT117), .ZN(n926) );
  NOR2_X1 U1022 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1023 ( .A(KEYINPUT118), .B(n928), .Z(n935) );
  XOR2_X1 U1024 ( .A(G164), .B(G2078), .Z(n932) );
  XNOR2_X1 U1025 ( .A(n930), .B(n929), .ZN(n931) );
  NOR2_X1 U1026 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1027 ( .A(KEYINPUT50), .B(n933), .Z(n934) );
  NOR2_X1 U1028 ( .A1(n935), .A2(n934), .ZN(n937) );
  NAND2_X1 U1029 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1030 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1031 ( .A(KEYINPUT52), .B(n940), .ZN(n941) );
  INV_X1 U1032 ( .A(KEYINPUT55), .ZN(n963) );
  NAND2_X1 U1033 ( .A1(n941), .A2(n963), .ZN(n942) );
  NAND2_X1 U1034 ( .A1(n942), .A2(G29), .ZN(n1026) );
  XOR2_X1 U1035 ( .A(G34), .B(KEYINPUT120), .Z(n944) );
  XNOR2_X1 U1036 ( .A(G2084), .B(KEYINPUT54), .ZN(n943) );
  XNOR2_X1 U1037 ( .A(n944), .B(n943), .ZN(n961) );
  XNOR2_X1 U1038 ( .A(G2090), .B(G35), .ZN(n959) );
  XOR2_X1 U1039 ( .A(G1991), .B(G25), .Z(n945) );
  NAND2_X1 U1040 ( .A1(n945), .A2(G28), .ZN(n956) );
  XNOR2_X1 U1041 ( .A(n946), .B(G27), .ZN(n949) );
  XNOR2_X1 U1042 ( .A(n947), .B(G32), .ZN(n948) );
  NAND2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1044 ( .A(KEYINPUT119), .B(n950), .ZN(n954) );
  XNOR2_X1 U1045 ( .A(G2067), .B(G26), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(G2072), .B(G33), .ZN(n951) );
  NOR2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1050 ( .A(KEYINPUT53), .B(n957), .ZN(n958) );
  NOR2_X1 U1051 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1052 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1053 ( .A(n963), .B(n962), .ZN(n965) );
  INV_X1 U1054 ( .A(G29), .ZN(n964) );
  NAND2_X1 U1055 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1056 ( .A1(G11), .A2(n966), .ZN(n1024) );
  XNOR2_X1 U1057 ( .A(G16), .B(KEYINPUT56), .ZN(n994) );
  XNOR2_X1 U1058 ( .A(G1341), .B(n967), .ZN(n968) );
  NOR2_X1 U1059 ( .A1(n969), .A2(n968), .ZN(n992) );
  XNOR2_X1 U1060 ( .A(G1348), .B(n970), .ZN(n984) );
  XNOR2_X1 U1061 ( .A(G1961), .B(G171), .ZN(n971) );
  XNOR2_X1 U1062 ( .A(n971), .B(KEYINPUT122), .ZN(n979) );
  XOR2_X1 U1063 ( .A(G1956), .B(KEYINPUT123), .Z(n972) );
  XNOR2_X1 U1064 ( .A(G299), .B(n972), .ZN(n977) );
  INV_X1 U1065 ( .A(n973), .ZN(n975) );
  NAND2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1068 ( .A1(n979), .A2(n978), .ZN(n982) );
  XNOR2_X1 U1069 ( .A(G1971), .B(G303), .ZN(n980) );
  XNOR2_X1 U1070 ( .A(KEYINPUT124), .B(n980), .ZN(n981) );
  NOR2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1072 ( .A1(n984), .A2(n983), .ZN(n990) );
  XNOR2_X1 U1073 ( .A(G1966), .B(G168), .ZN(n986) );
  NAND2_X1 U1074 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1075 ( .A(KEYINPUT121), .B(n987), .ZN(n988) );
  XNOR2_X1 U1076 ( .A(KEYINPUT57), .B(n988), .ZN(n989) );
  NOR2_X1 U1077 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1078 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1079 ( .A1(n994), .A2(n993), .ZN(n1022) );
  INV_X1 U1080 ( .A(G16), .ZN(n1020) );
  XOR2_X1 U1081 ( .A(G1986), .B(G24), .Z(n996) );
  XOR2_X1 U1082 ( .A(G1971), .B(G22), .Z(n995) );
  NAND2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n998) );
  XNOR2_X1 U1084 ( .A(G23), .B(G1976), .ZN(n997) );
  NOR2_X1 U1085 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1086 ( .A(KEYINPUT58), .B(n999), .Z(n1017) );
  XNOR2_X1 U1087 ( .A(KEYINPUT125), .B(G1981), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(n1000), .B(G6), .ZN(n1006) );
  XOR2_X1 U1089 ( .A(KEYINPUT126), .B(G4), .Z(n1002) );
  XNOR2_X1 U1090 ( .A(G1348), .B(KEYINPUT59), .ZN(n1001) );
  XNOR2_X1 U1091 ( .A(n1002), .B(n1001), .ZN(n1004) );
  XNOR2_X1 U1092 ( .A(G1341), .B(G19), .ZN(n1003) );
  NOR2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1008) );
  XNOR2_X1 U1095 ( .A(G20), .B(G1956), .ZN(n1007) );
  NOR2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1097 ( .A(KEYINPUT60), .B(n1009), .ZN(n1012) );
  XNOR2_X1 U1098 ( .A(n1010), .B(G5), .ZN(n1011) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  XNOR2_X1 U1100 ( .A(G21), .B(G1966), .ZN(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1102 ( .A(KEYINPUT127), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(KEYINPUT61), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1107 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1108 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1027), .Z(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

