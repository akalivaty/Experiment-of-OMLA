//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 0 1 1 1 0 0 1 1 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 0 1 1 1 0 1 0 0 1 1 1 1 0 0 0 0 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1256, new_n1257, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(KEYINPUT64), .ZN(new_n202));
  XNOR2_X1  g0002(.A(new_n201), .B(new_n202), .ZN(new_n203));
  INV_X1    g0003(.A(G77), .ZN(new_n204));
  AND2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G250), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  INV_X1    g0011(.A(G264), .ZN(new_n212));
  AOI211_X1 g0012(.A(new_n207), .B(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  OR2_X1    g0013(.A1(new_n213), .A2(KEYINPUT0), .ZN(new_n214));
  NOR2_X1   g0014(.A1(G58), .A2(G68), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  INV_X1    g0019(.A(G20), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n213), .A2(KEYINPUT0), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n214), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT65), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n226));
  INV_X1    g0026(.A(G68), .ZN(new_n227));
  INV_X1    g0027(.A(G238), .ZN(new_n228));
  INV_X1    g0028(.A(G87), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n226), .B1(new_n227), .B2(new_n228), .C1(new_n229), .C2(new_n207), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n231));
  INV_X1    g0031(.A(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G107), .ZN(new_n233));
  OAI221_X1 g0033(.A(new_n231), .B1(new_n204), .B2(new_n232), .C1(new_n233), .C2(new_n212), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n208), .B1(new_n230), .B2(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(KEYINPUT1), .Z(new_n236));
  NAND2_X1  g0036(.A1(new_n225), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G264), .B(G270), .Z(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G68), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  AOI21_X1  g0053(.A(new_n219), .B1(G33), .B2(G41), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n228), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n232), .A2(G1698), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT3), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n260), .A2(new_n262), .A3(KEYINPUT76), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT76), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(new_n259), .A3(G33), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n258), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G116), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n261), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n254), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G41), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(G1), .A3(G13), .ZN(new_n271));
  AND2_X1   g0071(.A1(new_n271), .A2(G274), .ZN(new_n272));
  INV_X1    g0072(.A(G45), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(G1), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(new_n207), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n272), .A2(new_n274), .B1(new_n275), .B2(new_n271), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n269), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT82), .ZN(new_n278));
  INV_X1    g0078(.A(G179), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT82), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n269), .A2(new_n280), .A3(new_n276), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n278), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT83), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n278), .A2(new_n281), .ZN(new_n285));
  INV_X1    g0085(.A(G169), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n278), .A2(KEYINPUT83), .A3(new_n279), .A4(new_n281), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT68), .B1(new_n208), .B2(new_n261), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT68), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n290), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n289), .A2(new_n219), .A3(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n263), .A2(new_n265), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n294), .A2(new_n220), .A3(G68), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n261), .A2(G20), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT19), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n296), .A2(new_n297), .A3(G97), .ZN(new_n298));
  NOR2_X1   g0098(.A1(G97), .A2(G107), .ZN(new_n299));
  NAND2_X1  g0099(.A1(G33), .A2(G97), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n299), .A2(new_n229), .B1(new_n300), .B2(new_n220), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n298), .B1(new_n301), .B2(new_n297), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n293), .B1(new_n295), .B2(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(KEYINPUT15), .B(G87), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G1), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n306), .A2(G13), .A3(G20), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n289), .A2(new_n219), .A3(new_n291), .A4(new_n307), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n306), .A2(G33), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n309), .B1(new_n304), .B2(new_n313), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n284), .A2(new_n287), .A3(new_n288), .A4(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n285), .A2(G200), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n313), .A2(new_n229), .ZN(new_n317));
  NOR3_X1   g0117(.A1(new_n317), .A2(new_n303), .A3(new_n308), .ZN(new_n318));
  INV_X1    g0118(.A(G190), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n316), .B(new_n318), .C1(new_n319), .C2(new_n285), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT84), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n315), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n306), .B1(G41), .B2(G45), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  AND3_X1   g0124(.A1(new_n324), .A2(new_n271), .A3(G274), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n271), .A2(new_n323), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n325), .B1(G226), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT3), .B(G33), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n330), .A2(G222), .A3(new_n255), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT67), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n331), .B(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n330), .A2(G1698), .ZN(new_n334));
  INV_X1    g0134(.A(G223), .ZN(new_n335));
  OAI22_X1  g0135(.A1(new_n334), .A2(new_n335), .B1(new_n204), .B2(new_n330), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n329), .B1(new_n338), .B2(new_n254), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G200), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n307), .A2(G50), .ZN(new_n342));
  NOR2_X1   g0142(.A1(G20), .A2(G33), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(G150), .ZN(new_n344));
  NOR2_X1   g0144(.A1(KEYINPUT8), .A2(G58), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  XNOR2_X1  g0146(.A(KEYINPUT69), .B(G58), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT8), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n296), .ZN(new_n350));
  OAI221_X1 g0150(.A(new_n344), .B1(new_n349), .B2(new_n350), .C1(new_n203), .C2(new_n220), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n342), .B1(new_n351), .B2(new_n292), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT70), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n310), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n310), .A2(new_n353), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n306), .A2(G20), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n355), .A2(new_n356), .A3(G50), .A4(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n352), .A2(KEYINPUT9), .A3(new_n358), .ZN(new_n359));
  OR2_X1    g0159(.A1(new_n331), .A2(new_n332), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n331), .A2(new_n332), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n336), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OAI211_X1 g0162(.A(G190), .B(new_n328), .C1(new_n362), .C2(new_n271), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT73), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n363), .A2(KEYINPUT73), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n341), .B(new_n359), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  AOI211_X1 g0167(.A(KEYINPUT72), .B(KEYINPUT9), .C1(new_n352), .C2(new_n358), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT72), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n351), .A2(new_n292), .ZN(new_n370));
  INV_X1    g0170(.A(new_n342), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(new_n358), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT9), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n369), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n368), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(KEYINPUT10), .B1(new_n367), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n372), .A2(new_n373), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT72), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n372), .A2(new_n369), .A3(new_n373), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT10), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT73), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n339), .A2(new_n382), .A3(G190), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n383), .A2(new_n364), .B1(new_n340), .B2(G200), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n380), .A2(new_n381), .A3(new_n359), .A4(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n376), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n340), .A2(new_n286), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n339), .A2(new_n279), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n387), .A2(new_n372), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(G226), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n255), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n330), .B(new_n392), .C1(G232), .C2(new_n255), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n300), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n254), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n324), .A2(new_n271), .A3(G274), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n326), .B2(new_n228), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT13), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n395), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT74), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n271), .B1(new_n393), .B2(new_n300), .ZN(new_n402));
  OAI21_X1  g0202(.A(KEYINPUT13), .B1(new_n402), .B2(new_n397), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n400), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  OAI211_X1 g0204(.A(KEYINPUT74), .B(KEYINPUT13), .C1(new_n402), .C2(new_n397), .ZN(new_n405));
  AND2_X1   g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT75), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT14), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n406), .A2(new_n407), .A3(new_n408), .A4(G169), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n404), .A2(new_n405), .A3(G169), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT75), .B1(new_n410), .B2(KEYINPUT14), .ZN(new_n411));
  AND3_X1   g0211(.A1(new_n400), .A2(G179), .A3(new_n403), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n412), .B1(new_n410), .B2(KEYINPUT14), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n409), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n350), .A2(new_n204), .ZN(new_n415));
  INV_X1    g0215(.A(new_n343), .ZN(new_n416));
  INV_X1    g0216(.A(G50), .ZN(new_n417));
  OAI22_X1  g0217(.A1(new_n416), .A2(new_n417), .B1(new_n220), .B2(G68), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n292), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT11), .ZN(new_n420));
  OR2_X1    g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n420), .ZN(new_n422));
  INV_X1    g0222(.A(new_n307), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n227), .ZN(new_n424));
  XNOR2_X1  g0224(.A(new_n424), .B(KEYINPUT12), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n311), .A2(G68), .A3(new_n357), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n421), .A2(new_n422), .A3(new_n425), .A4(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n414), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n406), .A2(G200), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n403), .A2(G190), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n427), .B1(new_n430), .B2(new_n400), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n216), .B1(new_n347), .B2(new_n227), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n434), .A2(G20), .B1(G159), .B2(new_n343), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT7), .ZN(new_n436));
  NOR3_X1   g0236(.A1(new_n261), .A2(KEYINPUT76), .A3(KEYINPUT3), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n437), .B1(new_n330), .B2(KEYINPUT76), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n436), .B1(new_n438), .B2(new_n220), .ZN(new_n439));
  AND2_X1   g0239(.A1(KEYINPUT77), .A2(KEYINPUT7), .ZN(new_n440));
  NOR2_X1   g0240(.A1(KEYINPUT77), .A2(KEYINPUT7), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n263), .A2(new_n220), .A3(new_n442), .A4(new_n265), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G68), .ZN(new_n444));
  OAI211_X1 g0244(.A(KEYINPUT16), .B(new_n435), .C1(new_n439), .C2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT16), .ZN(new_n446));
  INV_X1    g0246(.A(G58), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(KEYINPUT69), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT69), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(G58), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n215), .B1(new_n451), .B2(G68), .ZN(new_n452));
  INV_X1    g0252(.A(G159), .ZN(new_n453));
  OAI22_X1  g0253(.A1(new_n452), .A2(new_n220), .B1(new_n453), .B2(new_n416), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n442), .B1(new_n330), .B2(G20), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n259), .A2(G33), .ZN(new_n457));
  OAI211_X1 g0257(.A(KEYINPUT7), .B(new_n220), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n227), .B1(new_n455), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n446), .B1(new_n454), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n445), .A2(new_n460), .A3(new_n292), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n271), .A2(G232), .A3(new_n323), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n396), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n261), .A2(new_n229), .ZN(new_n464));
  NOR2_X1   g0264(.A1(G223), .A2(G1698), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n465), .B1(new_n391), .B2(G1698), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n464), .B1(new_n294), .B2(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n319), .B(new_n463), .C1(new_n467), .C2(new_n271), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n396), .A2(new_n462), .ZN(new_n469));
  INV_X1    g0269(.A(new_n464), .ZN(new_n470));
  INV_X1    g0270(.A(new_n466), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n470), .B1(new_n438), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n469), .B1(new_n472), .B2(new_n254), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n468), .B1(new_n473), .B2(G200), .ZN(new_n474));
  INV_X1    g0274(.A(new_n349), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n356), .A2(new_n357), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n475), .B1(new_n476), .B2(new_n354), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n349), .A2(new_n307), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n461), .A2(new_n474), .A3(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT78), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n461), .A2(new_n474), .A3(KEYINPUT78), .A4(new_n479), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(KEYINPUT17), .A3(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT17), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n461), .A2(new_n474), .A3(new_n485), .A4(new_n479), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n486), .A2(KEYINPUT79), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n461), .A2(new_n479), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT18), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n473), .A2(G179), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n491), .B1(new_n286), .B2(new_n473), .ZN(new_n492));
  AND3_X1   g0292(.A1(new_n489), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n490), .B1(new_n489), .B2(new_n492), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT79), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n482), .A2(new_n496), .A3(KEYINPUT17), .A4(new_n483), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n488), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n330), .A2(G232), .A3(new_n255), .ZN(new_n499));
  OAI221_X1 g0299(.A(new_n499), .B1(new_n233), .B2(new_n330), .C1(new_n334), .C2(new_n228), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n254), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n325), .B1(G244), .B2(new_n327), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n501), .A2(new_n279), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n311), .A2(G77), .A3(new_n357), .ZN(new_n504));
  XNOR2_X1  g0304(.A(KEYINPUT8), .B(G58), .ZN(new_n505));
  OAI22_X1  g0305(.A1(new_n505), .A2(new_n416), .B1(new_n220), .B2(new_n204), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n304), .A2(new_n350), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n292), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n423), .A2(new_n204), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n504), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  AND2_X1   g0310(.A1(new_n501), .A2(new_n502), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n503), .B(new_n510), .C1(new_n511), .C2(G169), .ZN(new_n512));
  INV_X1    g0312(.A(new_n510), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n501), .A2(G190), .A3(new_n502), .ZN(new_n514));
  INV_X1    g0314(.A(G200), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n513), .B(new_n514), .C1(new_n511), .C2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g0317(.A(new_n517), .B(KEYINPUT71), .ZN(new_n518));
  NOR4_X1   g0318(.A1(new_n390), .A2(new_n433), .A3(new_n498), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n315), .A2(new_n320), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT84), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n268), .A2(new_n220), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n233), .A2(KEYINPUT23), .A3(G20), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT23), .B1(new_n233), .B2(G20), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n229), .A2(G20), .ZN(new_n526));
  AOI21_X1  g0326(.A(KEYINPUT22), .B1(new_n330), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n294), .A2(KEYINPUT22), .A3(new_n220), .A4(G87), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT24), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n530), .B1(new_n528), .B2(new_n529), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n292), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(G13), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n535), .A2(G1), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n220), .A2(G107), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n538), .A2(KEYINPUT86), .A3(KEYINPUT25), .ZN(new_n539));
  OR2_X1    g0339(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n540));
  NAND2_X1  g0340(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n536), .A2(new_n537), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n539), .B(new_n542), .C1(new_n313), .C2(new_n233), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  AND2_X1   g0344(.A1(KEYINPUT5), .A2(G41), .ZN(new_n545));
  NOR2_X1   g0345(.A1(KEYINPUT5), .A2(G41), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n274), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n271), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n548), .A2(new_n212), .ZN(new_n549));
  NAND2_X1  g0349(.A1(G33), .A2(G294), .ZN(new_n550));
  NOR2_X1   g0350(.A1(G250), .A2(G1698), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n551), .B1(new_n211), .B2(G1698), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n550), .B1(new_n438), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n549), .B1(new_n554), .B2(new_n254), .ZN(new_n555));
  XNOR2_X1  g0355(.A(KEYINPUT5), .B(G41), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n556), .A2(new_n271), .A3(G274), .A4(new_n274), .ZN(new_n557));
  AOI21_X1  g0357(.A(G200), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n254), .B1(new_n274), .B2(new_n556), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(G264), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n294), .A2(new_n552), .B1(G33), .B2(G294), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n557), .B(new_n560), .C1(new_n561), .C2(new_n271), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n562), .A2(G190), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n534), .B(new_n544), .C1(new_n558), .C2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n311), .A2(G116), .A3(new_n312), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n423), .A2(new_n267), .ZN(new_n566));
  AOI21_X1  g0366(.A(G20), .B1(G33), .B2(G283), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n261), .A2(G97), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n567), .A2(new_n568), .B1(G20), .B2(new_n267), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n292), .A2(KEYINPUT20), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(KEYINPUT20), .B1(new_n292), .B2(new_n569), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n565), .B(new_n566), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n212), .A2(G1698), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(G257), .B2(G1698), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n574), .B1(new_n265), .B2(new_n263), .ZN(new_n575));
  INV_X1    g0375(.A(G303), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n330), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n254), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT85), .B1(new_n559), .B2(G270), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT85), .ZN(new_n580));
  INV_X1    g0380(.A(G270), .ZN(new_n581));
  NOR3_X1   g0381(.A1(new_n548), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n578), .B(new_n557), .C1(new_n579), .C2(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n572), .B1(new_n583), .B2(G200), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n319), .B2(new_n583), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n343), .A2(G77), .ZN(new_n586));
  XOR2_X1   g0386(.A(new_n586), .B(KEYINPUT80), .Z(new_n587));
  INV_X1    g0387(.A(KEYINPUT6), .ZN(new_n588));
  INV_X1    g0388(.A(G97), .ZN(new_n589));
  NOR3_X1   g0389(.A1(new_n588), .A2(new_n589), .A3(G107), .ZN(new_n590));
  XNOR2_X1  g0390(.A(G97), .B(G107), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n590), .B1(new_n588), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n587), .B1(new_n220), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n233), .B1(new_n455), .B2(new_n458), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n292), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n307), .A2(G97), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(new_n313), .B2(new_n589), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n232), .A2(G1698), .ZN(new_n601));
  AOI21_X1  g0401(.A(KEYINPUT4), .B1(new_n294), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n330), .A2(G250), .A3(G1698), .ZN(new_n603));
  NAND2_X1  g0403(.A1(G33), .A2(G283), .ZN(new_n604));
  AND2_X1   g0404(.A1(KEYINPUT4), .A2(G244), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n260), .A2(new_n262), .A3(new_n605), .A4(new_n255), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n603), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n254), .B1(new_n602), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n547), .A2(G257), .A3(new_n271), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n557), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(KEYINPUT81), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT81), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n609), .A2(new_n612), .A3(new_n557), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n608), .A2(new_n279), .A3(new_n611), .A4(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n607), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT4), .ZN(new_n616));
  INV_X1    g0416(.A(new_n601), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n616), .B1(new_n438), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n271), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n286), .B1(new_n619), .B2(new_n610), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n600), .A2(new_n614), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n455), .A2(new_n458), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(G107), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n623), .B(new_n587), .C1(new_n220), .C2(new_n592), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n598), .B1(new_n624), .B2(new_n292), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n611), .A2(new_n613), .ZN(new_n626));
  OAI21_X1  g0426(.A(G200), .B1(new_n626), .B2(new_n619), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n606), .A2(new_n604), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n617), .B1(new_n263), .B2(new_n265), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n628), .B(new_n603), .C1(new_n629), .C2(KEYINPUT4), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n610), .B1(new_n630), .B2(new_n254), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(G190), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n625), .A2(new_n627), .A3(new_n632), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n564), .A2(new_n585), .A3(new_n621), .A4(new_n633), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n578), .A2(new_n557), .ZN(new_n635));
  INV_X1    g0435(.A(new_n582), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n580), .B1(new_n548), .B2(new_n581), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n635), .A2(new_n572), .A3(new_n638), .A4(G179), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n583), .A2(new_n572), .A3(KEYINPUT21), .A4(G169), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n562), .A2(new_n286), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n555), .A2(new_n279), .A3(new_n557), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n528), .A2(new_n529), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(KEYINPUT24), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n293), .B1(new_n645), .B2(new_n531), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n642), .B(new_n643), .C1(new_n646), .C2(new_n543), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n583), .A2(G169), .A3(new_n572), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT21), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n641), .A2(new_n647), .A3(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n634), .A2(new_n651), .ZN(new_n652));
  AND4_X1   g0452(.A1(new_n322), .A2(new_n519), .A3(new_n521), .A4(new_n652), .ZN(G372));
  INV_X1    g0453(.A(new_n389), .ZN(new_n654));
  INV_X1    g0454(.A(new_n432), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(new_n512), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n656), .B1(new_n427), .B2(new_n414), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n488), .A2(new_n497), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n495), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n654), .B1(new_n659), .B2(new_n386), .ZN(new_n660));
  INV_X1    g0460(.A(new_n519), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT87), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n651), .A2(new_n662), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n564), .A2(new_n633), .A3(new_n621), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n277), .A2(G200), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n318), .B(new_n665), .C1(new_n285), .C2(new_n319), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n277), .A2(new_n286), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n314), .A2(new_n282), .A3(new_n667), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n641), .A2(new_n647), .A3(KEYINPUT87), .A4(new_n650), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n663), .A2(new_n664), .A3(new_n669), .A4(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n668), .ZN(new_n672));
  INV_X1    g0472(.A(new_n621), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n673), .A2(new_n668), .A3(new_n666), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT26), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n521), .A2(KEYINPUT26), .A3(new_n322), .A4(new_n673), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n672), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n660), .B1(new_n661), .B2(new_n678), .ZN(G369));
  NAND2_X1  g0479(.A1(new_n536), .A2(new_n220), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G213), .A3(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(G343), .ZN(new_n684));
  OR3_X1    g0484(.A1(new_n683), .A2(KEYINPUT88), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(KEYINPUT88), .B1(new_n683), .B2(new_n684), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n572), .ZN(new_n688));
  XOR2_X1   g0488(.A(new_n688), .B(KEYINPUT89), .Z(new_n689));
  AND2_X1   g0489(.A1(new_n641), .A2(new_n650), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(new_n690), .A3(new_n585), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n690), .B2(new_n689), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n692), .A2(G330), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n646), .A2(new_n543), .ZN(new_n694));
  INV_X1    g0494(.A(new_n687), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n647), .B(new_n564), .C1(new_n694), .C2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n647), .B2(new_n695), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n690), .A2(new_n687), .ZN(new_n699));
  INV_X1    g0499(.A(new_n696), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n647), .A2(new_n687), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n698), .A2(new_n704), .ZN(G399));
  NOR2_X1   g0505(.A1(new_n210), .A2(G41), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n299), .A2(new_n229), .A3(new_n267), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n706), .A2(new_n707), .A3(new_n306), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n708), .B1(new_n218), .B2(new_n706), .ZN(new_n709));
  XOR2_X1   g0509(.A(new_n709), .B(KEYINPUT28), .Z(new_n710));
  NAND3_X1  g0510(.A1(new_n664), .A2(new_n669), .A3(new_n651), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n674), .A2(KEYINPUT26), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n711), .A2(new_n668), .A3(new_n712), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n521), .A2(new_n675), .A3(new_n322), .A4(new_n673), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n715), .A2(KEYINPUT29), .A3(new_n695), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n678), .A2(new_n687), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n716), .B1(new_n717), .B2(KEYINPUT29), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT31), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n278), .A2(new_n631), .A3(new_n281), .A4(new_n555), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n635), .A2(G179), .A3(new_n638), .ZN(new_n721));
  OAI21_X1  g0521(.A(KEYINPUT30), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n610), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n555), .A2(new_n608), .A3(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n583), .A2(new_n279), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n269), .A2(new_n280), .A3(new_n276), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n280), .B1(new_n269), .B2(new_n276), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT30), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n725), .A2(new_n726), .A3(new_n729), .A4(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(G179), .B1(new_n269), .B2(new_n276), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n583), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n562), .B1(new_n626), .B2(new_n619), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT90), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI211_X1 g0536(.A(KEYINPUT90), .B(new_n562), .C1(new_n626), .C2(new_n619), .ZN(new_n737));
  AOI22_X1  g0537(.A1(new_n722), .A2(new_n731), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT91), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n687), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n722), .A2(new_n731), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n736), .A2(new_n737), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n741), .A2(new_n739), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n719), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n521), .A2(new_n652), .A3(new_n322), .A4(new_n695), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n724), .A2(new_n728), .A3(new_n727), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n730), .B1(new_n746), .B2(new_n726), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n720), .A2(KEYINPUT30), .A3(new_n721), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n742), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n749), .A2(KEYINPUT31), .A3(new_n687), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n744), .A2(new_n745), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G330), .ZN(new_n752));
  AND2_X1   g0552(.A1(new_n718), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n710), .B1(new_n753), .B2(G1), .ZN(G364));
  NOR2_X1   g0554(.A1(new_n535), .A2(G20), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n306), .B1(new_n755), .B2(G45), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n706), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT92), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n219), .B1(G20), .B2(new_n286), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n220), .A2(G179), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(G190), .A3(G200), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n229), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n319), .A2(G179), .A3(G200), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n220), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n765), .B1(G97), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G190), .A2(G200), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n763), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G159), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n763), .A2(new_n319), .A3(G200), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n769), .B1(KEYINPUT32), .B2(new_n773), .C1(new_n233), .C2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n220), .A2(new_n279), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(new_n770), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n776), .A2(G190), .A3(new_n515), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n330), .B1(new_n777), .B2(new_n204), .C1(new_n347), .C2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n776), .A2(G200), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n319), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n773), .A2(KEYINPUT32), .B1(new_n782), .B2(G50), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n781), .A2(G190), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  OAI211_X1 g0585(.A(new_n780), .B(new_n783), .C1(new_n227), .C2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(G283), .ZN(new_n787));
  INV_X1    g0587(.A(G329), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n774), .A2(new_n787), .B1(new_n771), .B2(new_n788), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n789), .B(KEYINPUT96), .Z(new_n790));
  INV_X1    g0590(.A(G322), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n778), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n777), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n330), .B(new_n792), .C1(G311), .C2(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(G294), .A2(new_n768), .B1(new_n782), .B2(G326), .ZN(new_n795));
  XNOR2_X1  g0595(.A(KEYINPUT33), .B(G317), .ZN(new_n796));
  INV_X1    g0596(.A(new_n764), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n784), .A2(new_n796), .B1(new_n797), .B2(G303), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n790), .A2(new_n794), .A3(new_n795), .A4(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n762), .B1(new_n786), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(G13), .A2(G33), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(G20), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n761), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT95), .ZN(new_n805));
  INV_X1    g0605(.A(new_n330), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(new_n210), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n807), .A2(G355), .B1(new_n267), .B2(new_n210), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n808), .B(KEYINPUT93), .Z(new_n809));
  NAND2_X1  g0609(.A1(new_n252), .A2(G45), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT94), .Z(new_n811));
  NOR2_X1   g0611(.A1(new_n294), .A2(new_n210), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(G45), .B2(new_n217), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n809), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n760), .B(new_n800), .C1(new_n805), .C2(new_n814), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(KEYINPUT97), .Z(new_n816));
  INV_X1    g0616(.A(new_n803), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n816), .B1(new_n692), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n693), .A2(new_n758), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(G330), .B2(new_n692), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT98), .ZN(G396));
  NAND2_X1  g0622(.A1(new_n687), .A2(new_n510), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n512), .A2(new_n516), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(KEYINPUT99), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT99), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n512), .A2(new_n516), .A3(new_n823), .A4(new_n826), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n512), .A2(new_n695), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n825), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n825), .A2(new_n827), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n695), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n717), .A2(new_n829), .B1(new_n678), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n758), .B1(new_n832), .B2(new_n752), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n752), .B2(new_n832), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n762), .A2(new_n802), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n759), .B1(G77), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n782), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n837), .A2(new_n576), .B1(new_n764), .B2(new_n233), .ZN(new_n838));
  INV_X1    g0638(.A(new_n774), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n838), .B1(G87), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n778), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n330), .B1(new_n841), .B2(G294), .ZN(new_n842));
  AOI22_X1  g0642(.A1(G116), .A2(new_n793), .B1(new_n772), .B2(G311), .ZN(new_n843));
  AOI22_X1  g0643(.A1(G97), .A2(new_n768), .B1(new_n784), .B2(G283), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n840), .A2(new_n842), .A3(new_n843), .A4(new_n844), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n841), .A2(G143), .B1(new_n793), .B2(G159), .ZN(new_n846));
  INV_X1    g0646(.A(G137), .ZN(new_n847));
  INV_X1    g0647(.A(G150), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n846), .B1(new_n837), .B2(new_n847), .C1(new_n848), .C2(new_n785), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT34), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n438), .B1(G132), .B2(new_n772), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n774), .A2(new_n227), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n347), .B2(new_n767), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(G50), .B2(new_n797), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n851), .A2(new_n852), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n849), .A2(new_n850), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n845), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n836), .B1(new_n859), .B2(new_n761), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n829), .B2(new_n802), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n834), .A2(new_n861), .ZN(G384));
  NOR2_X1   g0662(.A1(new_n755), .A2(new_n306), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n519), .B(new_n716), .C1(new_n717), .C2(KEYINPUT29), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n660), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n865), .B(KEYINPUT102), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n683), .B(KEYINPUT100), .ZN(new_n867));
  OR2_X1    g0667(.A1(new_n495), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n445), .A2(new_n292), .ZN(new_n869));
  OAI21_X1  g0669(.A(KEYINPUT7), .B1(new_n294), .B2(G20), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n870), .A2(G68), .A3(new_n443), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT16), .B1(new_n871), .B2(new_n435), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n479), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n683), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n498), .A2(new_n875), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n491), .B(new_n683), .C1(new_n286), .C2(new_n473), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n482), .A2(new_n878), .A3(new_n483), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT37), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT101), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT37), .B1(new_n489), .B2(new_n492), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n489), .A2(new_n867), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n882), .A2(new_n482), .A3(new_n483), .A4(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n880), .A2(new_n881), .A3(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n881), .B1(new_n880), .B2(new_n884), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n876), .B(KEYINPUT38), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n880), .A2(new_n884), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT101), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n885), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT38), .B1(new_n892), .B2(new_n876), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n687), .A2(new_n427), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n428), .A2(new_n432), .A3(new_n895), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n427), .B(new_n687), .C1(new_n655), .C2(new_n414), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n677), .A2(new_n676), .ZN(new_n899));
  INV_X1    g0699(.A(new_n668), .ZN(new_n900));
  AND3_X1   g0700(.A1(new_n664), .A2(new_n670), .A3(new_n669), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n900), .B1(new_n901), .B2(new_n663), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n831), .B1(new_n899), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n512), .A2(new_n687), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n898), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n883), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n498), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n489), .A2(new_n492), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n908), .A2(new_n883), .A3(new_n480), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT37), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n884), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n907), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT38), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n888), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT39), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n876), .B1(new_n886), .B2(new_n887), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n913), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(KEYINPUT39), .A3(new_n888), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n428), .A2(new_n687), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  OAI221_X1 g0723(.A(new_n868), .B1(new_n894), .B2(new_n905), .C1(new_n921), .C2(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n866), .B(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(G330), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT38), .B1(new_n907), .B2(new_n911), .ZN(new_n927));
  AOI22_X1  g0727(.A1(new_n891), .A2(new_n885), .B1(new_n498), .B2(new_n875), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n927), .B1(KEYINPUT38), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n749), .A2(KEYINPUT91), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n741), .A2(new_n739), .A3(new_n742), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n930), .A2(KEYINPUT31), .A3(new_n687), .A4(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n744), .A2(new_n745), .A3(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n829), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n934), .B1(new_n896), .B2(new_n897), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(KEYINPUT40), .B1(new_n929), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n919), .A2(new_n888), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT40), .ZN(new_n939));
  AND3_X1   g0739(.A1(new_n933), .A2(new_n935), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n519), .A2(new_n933), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n926), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n943), .B2(new_n942), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n863), .B1(new_n925), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n925), .B2(new_n945), .ZN(new_n947));
  INV_X1    g0747(.A(new_n592), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n948), .A2(KEYINPUT35), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(KEYINPUT35), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n949), .A2(G116), .A3(new_n221), .A4(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT36), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n218), .B(G77), .C1(new_n227), .C2(new_n347), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(G50), .B2(new_n227), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n954), .A2(G1), .A3(new_n535), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n947), .A2(new_n952), .A3(new_n955), .ZN(G367));
  OAI21_X1  g0756(.A(new_n805), .B1(new_n209), .B2(new_n304), .ZN(new_n957));
  INV_X1    g0757(.A(new_n812), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n958), .A2(new_n245), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n759), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n841), .A2(G150), .B1(new_n772), .B2(G137), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n961), .B(new_n330), .C1(new_n417), .C2(new_n777), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n784), .A2(G159), .B1(new_n839), .B2(G77), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n347), .B2(new_n764), .ZN(new_n964));
  INV_X1    g0764(.A(G143), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n837), .A2(new_n965), .B1(new_n227), .B2(new_n767), .ZN(new_n966));
  NOR3_X1   g0766(.A1(new_n962), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT108), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n764), .A2(new_n267), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT46), .ZN(new_n970));
  XNOR2_X1  g0770(.A(KEYINPUT107), .B(G311), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n837), .A2(new_n971), .B1(new_n774), .B2(new_n589), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(G294), .B2(new_n784), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n778), .A2(new_n576), .B1(new_n777), .B2(new_n787), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(G317), .B2(new_n772), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n294), .B1(new_n768), .B2(G107), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n973), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n968), .B1(new_n970), .B2(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT47), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n960), .B1(new_n979), .B2(new_n761), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n695), .A2(new_n318), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n669), .A2(new_n981), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n981), .A2(new_n668), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n980), .B1(new_n817), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n673), .A2(new_n687), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n633), .B(new_n621), .C1(new_n625), .C2(new_n695), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n704), .A2(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n989), .B(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT44), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n988), .B1(KEYINPUT105), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n703), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n992), .A2(KEYINPUT105), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n994), .A2(new_n995), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n991), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n1000), .A2(new_n698), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n698), .ZN(new_n1002));
  NOR3_X1   g0802(.A1(new_n991), .A2(new_n999), .A3(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n693), .A2(KEYINPUT106), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n701), .B1(new_n697), .B2(new_n699), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n693), .B(KEYINPUT106), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1007), .B1(new_n1008), .B2(new_n1006), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1004), .A2(new_n753), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(new_n753), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n706), .B(KEYINPUT41), .Z(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n757), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n699), .A2(new_n700), .A3(new_n988), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT42), .Z(new_n1016));
  INV_X1    g0816(.A(KEYINPUT43), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n984), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n621), .B1(new_n987), .B2(new_n647), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n695), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .A4(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT103), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1024));
  AND2_X1   g0824(.A1(new_n1016), .A2(new_n1020), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n984), .B(KEYINPUT43), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1023), .B(new_n1024), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1002), .A2(new_n988), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1027), .B(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n985), .B1(new_n1014), .B2(new_n1029), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT109), .Z(G387));
  NAND2_X1  g0831(.A1(new_n1009), .A2(new_n757), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n791), .A2(new_n837), .B1(new_n785), .B2(new_n971), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1033), .A2(KEYINPUT111), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(KEYINPUT111), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n841), .A2(G317), .B1(new_n793), .B2(G303), .ZN(new_n1036));
  AND3_X1   g0836(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1037), .A2(KEYINPUT48), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(KEYINPUT48), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n768), .A2(G283), .B1(new_n797), .B2(G294), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT49), .Z(new_n1042));
  AOI21_X1  g0842(.A(new_n294), .B1(G326), .B2(new_n772), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n267), .B2(new_n774), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n475), .A2(new_n784), .B1(G68), .B2(new_n793), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT110), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n305), .A2(new_n768), .B1(new_n782), .B2(G159), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n764), .A2(new_n204), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(G97), .B2(new_n839), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n841), .A2(G50), .B1(new_n772), .B2(G150), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1048), .A2(new_n1050), .A3(new_n294), .A4(new_n1051), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1047), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n761), .B1(new_n1045), .B2(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n807), .A2(new_n707), .B1(new_n233), .B2(new_n210), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n242), .A2(new_n273), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n505), .A2(G50), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT50), .Z(new_n1058));
  INV_X1    g0858(.A(new_n707), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1059), .B(new_n273), .C1(new_n227), .C2(new_n204), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n812), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1055), .B1(new_n1056), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n760), .B1(new_n1062), .B2(new_n805), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1054), .B(new_n1063), .C1(new_n697), .C2(new_n817), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n753), .A2(new_n1009), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n706), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n753), .A2(new_n1009), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1032), .B(new_n1064), .C1(new_n1066), .C2(new_n1067), .ZN(G393));
  OAI21_X1  g0868(.A(new_n1065), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1069), .A2(new_n706), .A3(new_n1010), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1004), .A2(new_n757), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n805), .B1(new_n589), .B2(new_n209), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n958), .A2(new_n249), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n759), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n837), .A2(new_n848), .B1(new_n453), .B2(new_n778), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT51), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n777), .A2(new_n505), .B1(new_n771), .B2(new_n965), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1077), .A2(new_n438), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n784), .A2(G50), .B1(new_n839), .B2(G87), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n768), .A2(G77), .B1(new_n797), .B2(G68), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1076), .A2(new_n1078), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(G317), .A2(new_n782), .B1(new_n841), .B2(G311), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT52), .Z(new_n1083));
  AOI22_X1  g0883(.A1(new_n768), .A2(G116), .B1(new_n793), .B2(G294), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1083), .B(new_n1084), .C1(new_n576), .C2(new_n785), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n806), .B1(new_n771), .B2(new_n791), .C1(new_n233), .C2(new_n774), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(G283), .B2(new_n797), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT112), .Z(new_n1088));
  OAI21_X1  g0888(.A(new_n1081), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1074), .B1(new_n1089), .B2(new_n761), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n988), .B2(new_n817), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1070), .A2(new_n1071), .A3(new_n1091), .ZN(G390));
  NAND3_X1  g0892(.A1(new_n933), .A2(new_n935), .A3(G330), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(KEYINPUT113), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT113), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n933), .A2(new_n935), .A3(new_n1095), .A4(G330), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n917), .A2(new_n920), .B1(new_n905), .B2(new_n923), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n831), .B1(new_n713), .B2(new_n714), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n898), .B1(new_n1099), .B2(new_n904), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1100), .A2(new_n915), .A3(new_n923), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1097), .B1(new_n1098), .B2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n751), .A2(new_n829), .A3(G330), .A4(new_n898), .ZN(new_n1104));
  AOI21_X1  g0904(.A(KEYINPUT39), .B1(new_n914), .B2(new_n888), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n894), .B2(KEYINPUT39), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n678), .A2(new_n831), .B1(new_n512), .B2(new_n687), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n922), .B1(new_n1107), .B2(new_n898), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1101), .B(new_n1104), .C1(new_n1106), .C2(new_n1108), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n1103), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n757), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n759), .B1(new_n475), .B2(new_n835), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(G128), .A2(new_n782), .B1(new_n841), .B2(G132), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT117), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n806), .B1(new_n772), .B2(G125), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n785), .B2(new_n847), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n767), .A2(new_n453), .B1(new_n774), .B2(new_n417), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  XOR2_X1   g0918(.A(KEYINPUT54), .B(G143), .Z(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT116), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n793), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n764), .A2(new_n848), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT53), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1114), .A2(new_n1118), .A3(new_n1121), .A4(new_n1123), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n785), .A2(new_n233), .B1(new_n777), .B2(new_n589), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT118), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n1125), .A2(new_n1126), .B1(new_n787), .B2(new_n837), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(new_n1126), .B2(new_n1125), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT119), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n767), .A2(new_n204), .B1(new_n778), .B2(new_n267), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT120), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n330), .B(new_n765), .C1(G294), .C2(new_n772), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1131), .A2(new_n854), .A3(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1124), .B1(new_n1129), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1112), .B1(new_n1134), .B2(new_n761), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n1106), .B2(new_n802), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT115), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n751), .A2(G330), .A3(new_n829), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n898), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1094), .A2(new_n1140), .A3(new_n1096), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1099), .A2(new_n904), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n1104), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n933), .A2(G330), .A3(new_n829), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n1139), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n1141), .A2(new_n1107), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n519), .A2(G330), .A3(new_n933), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n864), .A2(new_n660), .A3(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1137), .B1(new_n1110), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1141), .A2(new_n1107), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1148), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1103), .A2(new_n1153), .A3(new_n1109), .A4(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT114), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1155), .A2(new_n1156), .A3(new_n706), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1103), .A2(new_n1109), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1158), .A2(new_n1159), .A3(KEYINPUT115), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1150), .A2(new_n1157), .A3(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1156), .B1(new_n1155), .B2(new_n706), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1111), .B(new_n1136), .C1(new_n1161), .C2(new_n1162), .ZN(G378));
  INV_X1    g0963(.A(KEYINPUT123), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n372), .A2(new_n874), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n390), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n386), .A2(new_n389), .A3(new_n1165), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1169), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1165), .B1(new_n386), .B2(new_n389), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n654), .B(new_n1166), .C1(new_n376), .C2(new_n385), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1171), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1170), .A2(new_n1174), .ZN(new_n1175));
  AND2_X1   g0975(.A1(new_n933), .A2(new_n935), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n915), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1177), .A2(KEYINPUT40), .B1(new_n938), .B2(new_n940), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1175), .B1(new_n1178), .B2(new_n926), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n917), .A2(new_n922), .A3(new_n920), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n868), .B1(new_n894), .B2(new_n905), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1175), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n942), .A2(G330), .A3(new_n1183), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1179), .A2(new_n1182), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1182), .B1(new_n1179), .B2(new_n1184), .ZN(new_n1186));
  OAI21_X1  g0986(.A(KEYINPUT57), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1148), .B1(new_n1110), .B2(new_n1149), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1164), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1183), .B1(new_n942), .B2(G330), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n926), .B(new_n1175), .C1(new_n937), .C2(new_n941), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n924), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1179), .A2(new_n1182), .A3(new_n1184), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1154), .B1(new_n1158), .B2(new_n1146), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT57), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1194), .A2(new_n1195), .A3(KEYINPUT123), .A4(KEYINPUT57), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1189), .A2(new_n1198), .A3(new_n706), .A4(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1175), .A2(new_n801), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n758), .B1(G50), .B2(new_n835), .ZN(new_n1202));
  OR2_X1    g1002(.A1(new_n294), .A2(G41), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1203), .B(new_n417), .C1(G33), .C2(G41), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(G68), .A2(new_n768), .B1(new_n782), .B2(G116), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT121), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1049), .B1(G97), .B2(new_n784), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n347), .B2(new_n774), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n305), .A2(new_n793), .B1(new_n772), .B2(G283), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n233), .B2(new_n778), .ZN(new_n1210));
  NOR4_X1   g1010(.A1(new_n1206), .A2(new_n1208), .A3(new_n1203), .A4(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1204), .B1(new_n1211), .B2(KEYINPUT58), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT122), .ZN(new_n1213));
  OR2_X1    g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1120), .A2(new_n797), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n784), .A2(G132), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n841), .A2(G128), .B1(new_n793), .B2(G137), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G150), .A2(new_n768), .B1(new_n782), .B2(G125), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  OR2_X1    g1020(.A1(new_n1220), .A2(KEYINPUT59), .ZN(new_n1221));
  AOI211_X1 g1021(.A(G33), .B(G41), .C1(new_n772), .C2(G124), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n453), .B2(new_n774), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(new_n1220), .B2(KEYINPUT59), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1211), .A2(KEYINPUT58), .B1(new_n1221), .B2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1214), .A2(new_n1215), .A3(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1202), .B1(new_n1226), .B2(new_n761), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n1194), .A2(new_n757), .B1(new_n1201), .B2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1200), .A2(new_n1228), .ZN(G375));
  NAND2_X1  g1029(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1159), .A2(new_n1013), .A3(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n759), .B1(G68), .B2(new_n835), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n778), .A2(new_n787), .B1(new_n777), .B2(new_n233), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n330), .B(new_n1233), .C1(G303), .C2(new_n772), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n797), .A2(G97), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n784), .A2(G116), .B1(new_n782), .B2(G294), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n768), .A2(new_n305), .B1(new_n839), .B2(G77), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT124), .ZN(new_n1239));
  OR2_X1    g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n841), .A2(G137), .B1(new_n772), .B2(G128), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n848), .B2(new_n777), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(new_n784), .B2(new_n1120), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n767), .A2(new_n417), .B1(new_n764), .B2(new_n453), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n438), .B(new_n1244), .C1(new_n451), .C2(new_n839), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n782), .A2(G132), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1246), .B(KEYINPUT125), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1243), .A2(new_n1245), .A3(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1240), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1232), .B1(new_n1250), .B2(new_n761), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n898), .B2(new_n802), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n1146), .B2(new_n756), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1231), .A2(new_n1254), .ZN(G381));
  OR2_X1    g1055(.A1(G393), .A2(G396), .ZN(new_n1256));
  OR4_X1    g1056(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1256), .ZN(new_n1257));
  OR4_X1    g1057(.A1(G387), .A2(new_n1257), .A3(G378), .A4(G375), .ZN(G407));
  NAND2_X1  g1058(.A1(new_n1111), .A2(new_n1136), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1150), .A2(new_n1157), .A3(new_n1160), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1162), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1259), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n684), .A2(G213), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1265));
  OAI211_X1 g1065(.A(G407), .B(G213), .C1(G375), .C2(new_n1265), .ZN(G409));
  INV_X1    g1066(.A(KEYINPUT61), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1200), .A2(G378), .A3(new_n1228), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1194), .A2(new_n1195), .A3(new_n1013), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(KEYINPUT126), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT126), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1194), .A2(new_n1195), .A3(new_n1271), .A4(new_n1013), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1270), .A2(new_n1228), .A3(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1262), .A2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1264), .B1(new_n1268), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT60), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1230), .B1(new_n1149), .B2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1146), .A2(KEYINPUT60), .A3(new_n1148), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1277), .A2(new_n706), .A3(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1279), .A2(G384), .A3(new_n1254), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(G384), .B1(new_n1279), .B2(new_n1254), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1264), .A2(G2897), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  OAI211_X1 g1085(.A(G2897), .B(new_n1264), .C1(new_n1281), .C2(new_n1282), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1267), .B1(new_n1275), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1275), .A2(new_n1283), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT63), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(G393), .A2(G396), .ZN(new_n1293));
  AOI21_X1  g1093(.A(KEYINPUT109), .B1(new_n1256), .B2(new_n1293), .ZN(new_n1294));
  OR2_X1    g1094(.A1(new_n1294), .A2(G390), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1256), .A2(new_n1293), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(G390), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1295), .A2(new_n1030), .A3(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1030), .B1(new_n1295), .B2(new_n1297), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1275), .A2(KEYINPUT63), .A3(new_n1283), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1289), .A2(new_n1292), .A3(new_n1301), .A4(new_n1302), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1304));
  AND3_X1   g1104(.A1(new_n1275), .A2(new_n1283), .A3(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT127), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(KEYINPUT62), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1307), .B1(new_n1275), .B2(new_n1283), .ZN(new_n1308));
  NOR3_X1   g1108(.A1(new_n1305), .A2(new_n1288), .A3(new_n1308), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1303), .B1(new_n1309), .B2(new_n1301), .ZN(G405));
  NAND2_X1  g1110(.A1(G375), .A2(new_n1262), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n1268), .ZN(new_n1312));
  OR2_X1    g1112(.A1(new_n1312), .A2(new_n1283), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1283), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1301), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1313), .A2(new_n1301), .A3(new_n1314), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(G402));
endmodule


