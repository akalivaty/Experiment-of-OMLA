//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 0 1 1 0 0 0 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 1 0 0 1 1 1 0 0 1 1 0 0 1 1 1 0 1 0 0 1 0 1 1 0 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n796, new_n797, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975;
  INV_X1    g000(.A(KEYINPUT90), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT6), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT5), .ZN(new_n204));
  INV_X1    g003(.A(G134gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G127gat), .ZN(new_n206));
  INV_X1    g005(.A(G127gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G134gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G113gat), .B(G120gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n209), .B1(new_n210), .B2(KEYINPUT1), .ZN(new_n211));
  INV_X1    g010(.A(G120gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G113gat), .ZN(new_n213));
  INV_X1    g012(.A(G113gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G120gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G127gat), .B(G134gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT1), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n211), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221));
  INV_X1    g020(.A(G155gat), .ZN(new_n222));
  INV_X1    g021(.A(G162gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n221), .B1(new_n224), .B2(KEYINPUT2), .ZN(new_n225));
  AND2_X1   g024(.A1(G141gat), .A2(G148gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(G141gat), .A2(G148gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n221), .A2(KEYINPUT2), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT74), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT74), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n221), .A2(new_n232), .A3(KEYINPUT2), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n231), .A2(new_n228), .A3(new_n233), .ZN(new_n234));
  AND2_X1   g033(.A1(new_n224), .A2(new_n221), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n229), .A3(new_n236), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n234), .A2(new_n235), .B1(new_n228), .B2(new_n225), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n237), .B1(new_n238), .B2(new_n220), .ZN(new_n239));
  NAND2_X1  g038(.A1(G225gat), .A2(G233gat), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n204), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT4), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n220), .A2(new_n244), .A3(new_n229), .A4(new_n236), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT75), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n237), .A2(KEYINPUT4), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n229), .A2(new_n211), .A3(new_n219), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n249), .A2(KEYINPUT75), .A3(new_n244), .A4(new_n236), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n247), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n236), .A2(new_n229), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n220), .B1(new_n252), .B2(KEYINPUT3), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT3), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n236), .A2(new_n254), .A3(new_n229), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n241), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n251), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT76), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT76), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n251), .A2(new_n259), .A3(new_n256), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n243), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n248), .A2(new_n245), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n256), .A2(new_n204), .A3(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G1gat), .B(G29gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(KEYINPUT0), .ZN(new_n265));
  XNOR2_X1  g064(.A(G57gat), .B(G85gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n263), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n203), .B1(new_n261), .B2(new_n269), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n251), .A2(new_n259), .A3(new_n256), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n259), .B1(new_n251), .B2(new_n256), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n242), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n268), .B1(new_n273), .B2(new_n263), .ZN(new_n274));
  OAI21_X1  g073(.A(KEYINPUT80), .B1(new_n270), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n263), .ZN(new_n276));
  OAI211_X1 g075(.A(KEYINPUT6), .B(new_n267), .C1(new_n261), .C2(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n267), .B1(new_n261), .B2(new_n276), .ZN(new_n278));
  INV_X1    g077(.A(new_n269), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT6), .B1(new_n273), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT80), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n278), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n275), .A2(new_n277), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G211gat), .ZN(new_n284));
  INV_X1    g083(.A(G218gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(G211gat), .A2(G218gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT22), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G197gat), .B(G204gat), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n288), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n288), .A2(new_n291), .A3(new_n290), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G226gat), .A2(G233gat), .ZN(new_n297));
  XOR2_X1   g096(.A(new_n297), .B(KEYINPUT72), .Z(new_n298));
  INV_X1    g097(.A(KEYINPUT24), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n299), .A2(G183gat), .A3(G190gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(G169gat), .A2(G176gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT23), .ZN(new_n302));
  XNOR2_X1  g101(.A(G183gat), .B(G190gat), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n300), .B(new_n302), .C1(new_n303), .C2(new_n299), .ZN(new_n304));
  NAND2_X1  g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT66), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT66), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n307), .A2(G169gat), .A3(G176gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n309), .B1(KEYINPUT23), .B2(new_n301), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT25), .B1(new_n304), .B2(new_n310), .ZN(new_n311));
  XOR2_X1   g110(.A(KEYINPUT65), .B(G169gat), .Z(new_n312));
  INV_X1    g111(.A(G176gat), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n313), .A2(KEYINPUT23), .ZN(new_n314));
  AOI21_X1  g113(.A(KEYINPUT25), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  OR2_X1    g114(.A1(new_n303), .A2(new_n299), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n301), .A2(KEYINPUT23), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n317), .B1(new_n306), .B2(new_n308), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n315), .A2(new_n316), .A3(new_n318), .A4(new_n300), .ZN(new_n319));
  XNOR2_X1  g118(.A(KEYINPUT27), .B(G183gat), .ZN(new_n320));
  INV_X1    g119(.A(G190gat), .ZN(new_n321));
  AND3_X1   g120(.A1(new_n320), .A2(KEYINPUT28), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT28), .ZN(new_n323));
  INV_X1    g122(.A(G183gat), .ZN(new_n324));
  OAI21_X1  g123(.A(KEYINPUT67), .B1(new_n324), .B2(KEYINPUT27), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n321), .B(new_n325), .C1(new_n320), .C2(KEYINPUT67), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n322), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(KEYINPUT68), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT26), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n301), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n309), .A2(new_n331), .ZN(new_n332));
  OAI22_X1  g131(.A1(new_n329), .A2(new_n332), .B1(new_n324), .B2(new_n321), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n311), .B(new_n319), .C1(new_n327), .C2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(KEYINPUT73), .B(KEYINPUT29), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n298), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  AND2_X1   g135(.A1(new_n319), .A2(new_n311), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT68), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n328), .B(new_n338), .ZN(new_n339));
  AOI22_X1  g138(.A1(new_n306), .A2(new_n308), .B1(new_n330), .B2(new_n301), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n339), .A2(new_n340), .B1(G183gat), .B2(G190gat), .ZN(new_n341));
  XOR2_X1   g140(.A(KEYINPUT27), .B(G183gat), .Z(new_n342));
  INV_X1    g141(.A(KEYINPUT67), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AND2_X1   g143(.A1(new_n325), .A2(new_n321), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT28), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n341), .B1(new_n346), .B2(new_n322), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n297), .B1(new_n337), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n296), .B1(new_n336), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n298), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT29), .B1(new_n337), .B2(new_n347), .ZN(new_n351));
  INV_X1    g150(.A(new_n297), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n295), .B(new_n350), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G8gat), .B(G36gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(G64gat), .B(G92gat), .ZN(new_n357));
  XOR2_X1   g156(.A(new_n356), .B(new_n357), .Z(new_n358));
  NAND2_X1  g157(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT30), .ZN(new_n360));
  INV_X1    g159(.A(new_n358), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n360), .B1(new_n354), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n355), .A2(new_n360), .A3(new_n358), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n283), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT82), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT82), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n283), .A2(new_n368), .A3(new_n365), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  XOR2_X1   g169(.A(G15gat), .B(G43gat), .Z(new_n371));
  XNOR2_X1  g170(.A(G71gat), .B(G99gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G227gat), .A2(G233gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n374), .B(KEYINPUT64), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n220), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n334), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n347), .A2(new_n220), .A3(new_n311), .A4(new_n319), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n376), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n373), .B1(new_n380), .B2(KEYINPUT33), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT32), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  OR2_X1    g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n378), .A2(new_n379), .ZN(new_n385));
  INV_X1    g184(.A(new_n374), .ZN(new_n386));
  OAI21_X1  g185(.A(KEYINPUT34), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT69), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n375), .A2(KEYINPUT34), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n378), .A2(new_n388), .A3(new_n379), .A4(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n378), .A2(new_n379), .A3(new_n389), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT69), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n387), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  AOI221_X4 g192(.A(new_n382), .B1(KEYINPUT33), .B2(new_n373), .C1(new_n385), .C2(new_n375), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n384), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT71), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n381), .A2(new_n383), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n399), .A2(new_n394), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n400), .A2(KEYINPUT71), .A3(new_n393), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n387), .A2(new_n390), .A3(new_n392), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n403), .B1(new_n399), .B2(new_n394), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(G228gat), .A2(G233gat), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n295), .B1(new_n255), .B2(new_n335), .ZN(new_n407));
  INV_X1    g206(.A(new_n294), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n335), .B1(new_n408), .B2(new_n292), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n238), .B1(new_n409), .B2(new_n254), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n406), .B1(new_n407), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n406), .B1(new_n252), .B2(KEYINPUT3), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT29), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n295), .A2(new_n252), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n335), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n415), .B1(new_n238), .B2(new_n254), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n412), .B(new_n414), .C1(new_n295), .C2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(G22gat), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n411), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n418), .B1(new_n411), .B2(new_n417), .ZN(new_n420));
  OAI21_X1  g219(.A(G78gat), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n411), .A2(new_n417), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(G22gat), .ZN(new_n423));
  INV_X1    g222(.A(G78gat), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n411), .A2(new_n417), .A3(new_n418), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT31), .B(G50gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n427), .B(KEYINPUT77), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n428), .B(G106gat), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n421), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n429), .B1(new_n421), .B2(new_n426), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NOR3_X1   g232(.A1(new_n405), .A2(KEYINPUT35), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n393), .A2(KEYINPUT70), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT70), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n403), .A2(new_n436), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n435), .B(new_n437), .C1(new_n399), .C2(new_n394), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT71), .B1(new_n400), .B2(new_n393), .ZN(new_n439));
  NOR4_X1   g238(.A1(new_n399), .A2(new_n403), .A3(new_n394), .A4(new_n397), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n432), .B(new_n438), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT83), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT83), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n402), .A2(new_n443), .A3(new_n432), .A4(new_n438), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n277), .B1(new_n270), .B2(new_n274), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n365), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n442), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  AOI22_X1  g247(.A1(new_n370), .A2(new_n434), .B1(new_n448), .B2(KEYINPUT35), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n354), .A2(new_n361), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n354), .A2(new_n361), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n361), .A2(KEYINPUT37), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n295), .B1(new_n336), .B2(new_n348), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n296), .B(new_n350), .C1(new_n351), .C2(new_n352), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n454), .A2(new_n455), .A3(KEYINPUT37), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT38), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n450), .B1(new_n453), .B2(new_n458), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n275), .A2(new_n277), .A3(new_n282), .A4(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT81), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n453), .A2(new_n458), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n462), .A2(new_n277), .A3(new_n359), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT81), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n463), .A2(new_n464), .A3(new_n275), .A4(new_n282), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n354), .A2(KEYINPUT37), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n361), .B1(new_n354), .B2(KEYINPUT37), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT38), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n461), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n365), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT39), .B1(new_n239), .B2(new_n241), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT79), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n253), .A2(new_n255), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n240), .B1(new_n262), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n471), .A2(new_n472), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n473), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT39), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n267), .B1(new_n475), .B2(new_n479), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n478), .A2(KEYINPUT40), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT40), .B1(new_n478), .B2(new_n480), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n481), .A2(new_n482), .A3(new_n274), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n470), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(new_n432), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n469), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT36), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT78), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n490), .B1(new_n430), .B2(new_n431), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n421), .A2(new_n426), .ZN(new_n492));
  INV_X1    g291(.A(new_n429), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n421), .A2(new_n426), .A3(new_n429), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n494), .A2(KEYINPUT78), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(new_n446), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT36), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n402), .A2(new_n499), .A3(new_n404), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n489), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n449), .B1(new_n487), .B2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G15gat), .B(G22gat), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT87), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(G1gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n504), .A2(new_n505), .A3(G1gat), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT16), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n508), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(G8gat), .ZN(new_n513));
  NOR2_X1   g312(.A1(G29gat), .A2(G36gat), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT14), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n514), .B(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(G29gat), .A2(G36gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n517), .B(KEYINPUT85), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT15), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n516), .A2(KEYINPUT15), .A3(new_n518), .ZN(new_n522));
  XNOR2_X1  g321(.A(G43gat), .B(G50gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  OR2_X1    g323(.A1(new_n522), .A2(new_n523), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n513), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(KEYINPUT86), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT17), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n526), .A2(KEYINPUT86), .A3(KEYINPUT17), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(G8gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n512), .B(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n527), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(G229gat), .A2(G233gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT18), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n513), .A2(new_n526), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n527), .A2(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n536), .B(KEYINPUT13), .Z(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(KEYINPUT89), .A3(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n541), .B1(new_n527), .B2(new_n539), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT89), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI22_X1  g344(.A1(new_n537), .A2(new_n538), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT88), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n535), .A2(new_n547), .A3(KEYINPUT18), .A4(new_n536), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n526), .A2(KEYINPUT86), .A3(KEYINPUT17), .ZN(new_n549));
  AOI21_X1  g348(.A(KEYINPUT17), .B1(new_n526), .B2(KEYINPUT86), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n534), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n527), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n551), .A2(KEYINPUT18), .A3(new_n536), .A4(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT88), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n548), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n546), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G113gat), .B(G141gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G169gat), .B(G197gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n561), .B(KEYINPUT12), .Z(new_n562));
  NAND2_X1  g361(.A1(new_n556), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n562), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n546), .A2(new_n555), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n202), .B1(new_n503), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n370), .A2(new_n434), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n448), .A2(KEYINPUT35), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n468), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n572), .B1(new_n460), .B2(KEYINPUT81), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n485), .B1(new_n573), .B2(new_n465), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n571), .B1(new_n574), .B2(new_n501), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n575), .A2(KEYINPUT90), .A3(new_n566), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n568), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G57gat), .B(G64gat), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT93), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G71gat), .A2(G78gat), .ZN(new_n581));
  INV_X1    g380(.A(G71gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(new_n424), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT9), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n581), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n578), .A2(new_n579), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n580), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n584), .B1(new_n578), .B2(KEYINPUT91), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n588), .B1(KEYINPUT91), .B2(new_n578), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT92), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n583), .A2(new_n581), .ZN(new_n591));
  AND3_X1   g390(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n590), .B1(new_n589), .B2(new_n591), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n587), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT21), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(G231gat), .A2(G233gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G127gat), .B(G155gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT20), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n598), .B(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n534), .B1(new_n594), .B2(new_n595), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT95), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n601), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G183gat), .B(G211gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n604), .B(new_n607), .Z(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G190gat), .B(G218gat), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT97), .B(G92gat), .ZN(new_n612));
  INV_X1    g411(.A(G85gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(G99gat), .A2(G106gat), .ZN(new_n614));
  AOI22_X1  g413(.A1(new_n612), .A2(new_n613), .B1(KEYINPUT8), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(G85gat), .A2(G92gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT7), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G99gat), .B(G106gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT98), .ZN(new_n620));
  OAI21_X1  g419(.A(KEYINPUT99), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT98), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n619), .B(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT99), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n623), .A2(new_n624), .A3(new_n617), .A4(new_n615), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n618), .A2(new_n620), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n628), .B1(new_n549), .B2(new_n550), .ZN(new_n629));
  AOI22_X1  g428(.A1(new_n621), .A2(new_n625), .B1(new_n620), .B2(new_n618), .ZN(new_n630));
  NAND2_X1  g429(.A1(G232gat), .A2(G233gat), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  AOI22_X1  g431(.A1(new_n630), .A2(new_n526), .B1(KEYINPUT41), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n611), .B1(new_n629), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n632), .A2(KEYINPUT41), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n636), .B(KEYINPUT96), .Z(new_n637));
  XNOR2_X1  g436(.A(G134gat), .B(G162gat), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n637), .B(new_n638), .Z(new_n639));
  NAND3_X1  g438(.A1(new_n629), .A2(new_n611), .A3(new_n633), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n635), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n640), .B1(new_n634), .B2(new_n642), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n629), .A2(KEYINPUT100), .A3(new_n611), .A4(new_n633), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n639), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT101), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI211_X1 g446(.A(KEYINPUT101), .B(new_n639), .C1(new_n643), .C2(new_n644), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n641), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT10), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n628), .A2(new_n594), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n620), .A2(KEYINPUT102), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT102), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n623), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n652), .A2(new_n654), .A3(new_n618), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n626), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n593), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n656), .A2(new_n659), .A3(new_n587), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n594), .A2(new_n630), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g461(.A(KEYINPUT103), .B(KEYINPUT10), .Z(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n651), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(G230gat), .A2(G233gat), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(KEYINPUT106), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n660), .A2(new_n667), .A3(new_n661), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT106), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n663), .B1(new_n660), .B2(new_n661), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n670), .B(new_n666), .C1(new_n671), .C2(new_n651), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n668), .A2(new_n669), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g472(.A(G120gat), .B(G148gat), .Z(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT105), .ZN(new_n675));
  XNOR2_X1  g474(.A(G176gat), .B(G204gat), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n675), .B(new_n676), .Z(new_n677));
  NAND2_X1  g476(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n665), .A2(KEYINPUT104), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT104), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n680), .B1(new_n671), .B2(new_n651), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n679), .A2(new_n666), .A3(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n677), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n682), .A2(new_n669), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n678), .A2(new_n684), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n609), .A2(new_n649), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n577), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(new_n445), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(new_n507), .ZN(G1324gat));
  AND2_X1   g488(.A1(new_n577), .A2(new_n686), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n533), .B1(new_n690), .B2(new_n470), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT16), .B(G8gat), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n687), .A2(new_n365), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT42), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n694), .B1(KEYINPUT42), .B2(new_n693), .ZN(G1325gat));
  INV_X1    g494(.A(G15gat), .ZN(new_n696));
  INV_X1    g495(.A(new_n405), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n690), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n489), .A2(new_n500), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n687), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n698), .B1(new_n696), .B2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT107), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  OAI211_X1 g502(.A(new_n698), .B(KEYINPUT107), .C1(new_n696), .C2(new_n700), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(G1326gat));
  INV_X1    g504(.A(new_n497), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n687), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g506(.A(KEYINPUT43), .B(G22gat), .Z(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(G1327gat));
  XNOR2_X1  g508(.A(new_n685), .B(KEYINPUT109), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n609), .A2(new_n566), .A3(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT111), .ZN(new_n713));
  OAI21_X1  g512(.A(KEYINPUT110), .B1(new_n574), .B2(new_n501), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT110), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n487), .A2(new_n715), .A3(new_n502), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n449), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n649), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n713), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n715), .B1(new_n487), .B2(new_n502), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n574), .A2(KEYINPUT110), .A3(new_n501), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n571), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n719), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n723), .A2(KEYINPUT111), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n720), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n718), .B1(new_n575), .B2(new_n649), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n712), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(G29gat), .B1(new_n730), .B2(new_n445), .ZN(new_n731));
  INV_X1    g530(.A(new_n685), .ZN(new_n732));
  AND4_X1   g531(.A1(KEYINPUT108), .A2(new_n609), .A3(new_n649), .A4(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n608), .A2(new_n685), .ZN(new_n734));
  AOI21_X1  g533(.A(KEYINPUT108), .B1(new_n734), .B2(new_n649), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n736), .B1(new_n568), .B2(new_n576), .ZN(new_n737));
  INV_X1    g536(.A(G29gat), .ZN(new_n738));
  INV_X1    g537(.A(new_n445), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n737), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT45), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OR2_X1    g541(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n731), .A2(new_n742), .A3(new_n743), .ZN(G1328gat));
  INV_X1    g543(.A(KEYINPUT112), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n365), .A2(G36gat), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n737), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n745), .B1(new_n737), .B2(new_n746), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT113), .ZN(new_n749));
  OAI22_X1  g548(.A1(new_n747), .A2(new_n748), .B1(new_n749), .B2(KEYINPUT46), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(KEYINPUT46), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n749), .B(KEYINPUT46), .C1(new_n747), .C2(new_n748), .ZN(new_n753));
  OAI21_X1  g552(.A(G36gat), .B1(new_n730), .B2(new_n365), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(G1329gat));
  INV_X1    g554(.A(KEYINPUT47), .ZN(new_n756));
  INV_X1    g555(.A(G43gat), .ZN(new_n757));
  INV_X1    g556(.A(new_n699), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n757), .B1(new_n729), .B2(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n737), .A2(new_n757), .A3(new_n697), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n756), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT114), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n763), .B1(new_n729), .B2(new_n758), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n727), .B1(new_n720), .B2(new_n725), .ZN(new_n765));
  NOR4_X1   g564(.A1(new_n765), .A2(KEYINPUT114), .A3(new_n699), .A4(new_n712), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n764), .A2(new_n766), .A3(new_n757), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n760), .A2(KEYINPUT47), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n762), .B1(new_n767), .B2(new_n768), .ZN(G1330gat));
  INV_X1    g568(.A(new_n737), .ZN(new_n770));
  INV_X1    g569(.A(G50gat), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n497), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT115), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n765), .A2(new_n432), .A3(new_n712), .ZN(new_n774));
  OAI221_X1 g573(.A(KEYINPUT48), .B1(new_n770), .B2(new_n773), .C1(new_n774), .C2(new_n771), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n770), .A2(new_n773), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n729), .A2(new_n497), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n776), .B1(G50gat), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n775), .B1(new_n778), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g578(.A(new_n649), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n608), .A2(new_n567), .A3(new_n780), .A4(new_n710), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n717), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n739), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(G57gat), .ZN(G1332gat));
  INV_X1    g583(.A(KEYINPUT49), .ZN(new_n785));
  INV_X1    g584(.A(G64gat), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n470), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT116), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n782), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n785), .A2(new_n786), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n789), .B(new_n790), .ZN(G1333gat));
  AOI21_X1  g590(.A(new_n582), .B1(new_n782), .B2(new_n758), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n405), .A2(G71gat), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n792), .B1(new_n782), .B2(new_n793), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g594(.A1(new_n782), .A2(new_n497), .ZN(new_n796));
  XNOR2_X1  g595(.A(KEYINPUT117), .B(G78gat), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n796), .B(new_n797), .ZN(G1335gat));
  NOR2_X1   g597(.A1(new_n608), .A2(new_n566), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n685), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n800), .B1(new_n726), .B2(new_n728), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(G85gat), .B1(new_n802), .B2(new_n445), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n723), .A2(KEYINPUT51), .A3(new_n649), .A4(new_n799), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n799), .A2(new_n649), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n805), .B1(new_n717), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n685), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n739), .A2(new_n613), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n803), .B1(new_n809), .B2(new_n810), .ZN(G1336gat));
  OR2_X1    g610(.A1(KEYINPUT118), .A2(KEYINPUT52), .ZN(new_n812));
  NAND2_X1  g611(.A1(KEYINPUT118), .A2(KEYINPUT52), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n612), .B1(new_n801), .B2(new_n470), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n711), .B1(new_n804), .B2(new_n807), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n365), .A2(G92gat), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n812), .B(new_n813), .C1(new_n814), .C2(new_n818), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n717), .A2(new_n713), .A3(new_n719), .ZN(new_n820));
  AOI21_X1  g619(.A(KEYINPUT111), .B1(new_n723), .B2(new_n724), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n728), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n800), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n822), .A2(new_n470), .A3(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n612), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n826), .A2(KEYINPUT118), .A3(KEYINPUT52), .A4(new_n817), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n819), .A2(new_n827), .ZN(G1337gat));
  OAI21_X1  g627(.A(G99gat), .B1(new_n802), .B2(new_n699), .ZN(new_n829));
  OR2_X1    g628(.A1(new_n405), .A2(G99gat), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n829), .B1(new_n809), .B2(new_n830), .ZN(G1338gat));
  XOR2_X1   g630(.A(KEYINPUT119), .B(G106gat), .Z(new_n832));
  OAI21_X1  g631(.A(new_n832), .B1(new_n802), .B2(new_n432), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n432), .A2(G106gat), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT53), .B1(new_n815), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n801), .A2(new_n497), .ZN(new_n837));
  AOI22_X1  g636(.A1(new_n837), .A2(new_n832), .B1(new_n815), .B2(new_n834), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT53), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n836), .B1(new_n838), .B2(new_n839), .ZN(G1339gat));
  NAND2_X1  g639(.A1(new_n668), .A2(new_n672), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n842), .B1(new_n665), .B2(new_n667), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n682), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n843), .A2(new_n677), .A3(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT55), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n843), .A2(new_n845), .A3(KEYINPUT55), .A4(new_n677), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n848), .A2(new_n566), .A3(new_n684), .A4(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n535), .A2(new_n536), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n540), .A2(new_n541), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n561), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n565), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n685), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n649), .B1(new_n850), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n848), .A2(new_n684), .A3(new_n849), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n649), .A2(new_n854), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n609), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n608), .A2(new_n567), .A3(new_n780), .A4(new_n732), .ZN(new_n861));
  AOI211_X1 g660(.A(new_n497), .B(new_n405), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n470), .A2(new_n445), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n862), .A2(KEYINPUT120), .A3(new_n863), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n868), .A2(new_n214), .A3(new_n567), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n445), .B1(new_n860), .B2(new_n861), .ZN(new_n870));
  AND4_X1   g669(.A1(new_n365), .A2(new_n870), .A3(new_n442), .A4(new_n444), .ZN(new_n871));
  AOI21_X1  g670(.A(G113gat), .B1(new_n871), .B2(new_n566), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n869), .A2(new_n872), .ZN(G1340gat));
  NOR2_X1   g672(.A1(new_n711), .A2(new_n212), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n866), .A2(new_n867), .A3(new_n874), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n871), .A2(new_n685), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n875), .B1(G120gat), .B2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT121), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n877), .B(new_n878), .ZN(G1341gat));
  OAI21_X1  g678(.A(G127gat), .B1(new_n868), .B2(new_n609), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n871), .A2(new_n207), .A3(new_n608), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(G1342gat));
  NAND3_X1  g681(.A1(new_n871), .A2(new_n205), .A3(new_n649), .ZN(new_n883));
  XOR2_X1   g682(.A(new_n883), .B(KEYINPUT56), .Z(new_n884));
  OAI21_X1  g683(.A(G134gat), .B1(new_n868), .B2(new_n780), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(G1343gat));
  NAND2_X1  g685(.A1(new_n699), .A2(new_n863), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n432), .B1(new_n860), .B2(new_n861), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT122), .ZN(new_n891));
  OAI22_X1  g690(.A1(new_n856), .A2(new_n891), .B1(new_n857), .B2(new_n858), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n856), .A2(new_n891), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n609), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n706), .B1(new_n894), .B2(new_n861), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n890), .B1(new_n895), .B2(new_n889), .ZN(new_n896));
  OAI21_X1  g695(.A(G141gat), .B1(new_n896), .B2(new_n567), .ZN(new_n897));
  AND4_X1   g696(.A1(new_n433), .A2(new_n870), .A3(new_n365), .A4(new_n699), .ZN(new_n898));
  INV_X1    g697(.A(G141gat), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n898), .A2(new_n899), .A3(new_n566), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(KEYINPUT58), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT58), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n897), .A2(new_n903), .A3(new_n900), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(G1344gat));
  NAND2_X1  g704(.A1(new_n860), .A2(new_n861), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n433), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n706), .A2(KEYINPUT57), .ZN(new_n908));
  AOI22_X1  g707(.A1(new_n907), .A2(KEYINPUT57), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  AND4_X1   g708(.A1(new_n699), .A2(new_n909), .A3(new_n685), .A4(new_n863), .ZN(new_n910));
  INV_X1    g709(.A(G148gat), .ZN(new_n911));
  OAI21_X1  g710(.A(KEYINPUT59), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n911), .A2(KEYINPUT59), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n913), .B1(new_n896), .B2(new_n732), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n898), .A2(new_n911), .A3(new_n685), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(G1345gat));
  OAI21_X1  g716(.A(G155gat), .B1(new_n896), .B2(new_n609), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n898), .A2(new_n222), .A3(new_n608), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(G1346gat));
  OR3_X1    g719(.A1(new_n896), .A2(new_n223), .A3(new_n780), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(G162gat), .B1(new_n898), .B2(new_n649), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n922), .A2(new_n923), .ZN(G1347gat));
  AOI21_X1  g723(.A(new_n739), .B1(new_n860), .B2(new_n861), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n442), .A2(new_n444), .A3(new_n470), .ZN(new_n926));
  XOR2_X1   g725(.A(new_n926), .B(KEYINPUT123), .Z(new_n927));
  AND2_X1   g726(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n928), .A2(new_n312), .A3(new_n566), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT124), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n739), .A2(new_n365), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n862), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(G169gat), .B1(new_n932), .B2(new_n567), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n930), .A2(new_n933), .ZN(G1348gat));
  OAI21_X1  g733(.A(G176gat), .B1(new_n932), .B2(new_n711), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n928), .A2(new_n313), .A3(new_n685), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1349gat));
  NAND4_X1  g736(.A1(new_n925), .A2(new_n320), .A3(new_n608), .A4(new_n927), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT125), .ZN(new_n939));
  OAI21_X1  g738(.A(G183gat), .B1(new_n932), .B2(new_n609), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g741(.A1(new_n928), .A2(new_n321), .A3(new_n649), .ZN(new_n943));
  OAI21_X1  g742(.A(G190gat), .B1(new_n932), .B2(new_n780), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n944), .A2(KEYINPUT61), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n944), .A2(KEYINPUT61), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n943), .B1(new_n945), .B2(new_n946), .ZN(G1351gat));
  NAND2_X1  g746(.A1(new_n906), .A2(new_n908), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n699), .A2(new_n931), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n948), .B(new_n949), .C1(new_n889), .C2(new_n888), .ZN(new_n950));
  OAI21_X1  g749(.A(KEYINPUT126), .B1(new_n950), .B2(new_n567), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT126), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n909), .A2(new_n952), .A3(new_n566), .A4(new_n949), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n951), .A2(new_n953), .A3(G197gat), .ZN(new_n954));
  AND4_X1   g753(.A1(new_n433), .A2(new_n925), .A3(new_n470), .A4(new_n699), .ZN(new_n955));
  INV_X1    g754(.A(G197gat), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n955), .A2(new_n956), .A3(new_n566), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT127), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n954), .A2(KEYINPUT127), .A3(new_n957), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(G1352gat));
  INV_X1    g761(.A(G204gat), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n955), .A2(new_n963), .A3(new_n685), .ZN(new_n964));
  XOR2_X1   g763(.A(new_n964), .B(KEYINPUT62), .Z(new_n965));
  OAI21_X1  g764(.A(G204gat), .B1(new_n950), .B2(new_n711), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(G1353gat));
  NAND3_X1  g766(.A1(new_n955), .A2(new_n284), .A3(new_n608), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n909), .A2(new_n608), .A3(new_n949), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n969), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g770(.A(KEYINPUT63), .B1(new_n969), .B2(G211gat), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n968), .B1(new_n971), .B2(new_n972), .ZN(G1354gat));
  OAI21_X1  g772(.A(G218gat), .B1(new_n950), .B2(new_n780), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n955), .A2(new_n285), .A3(new_n649), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(G1355gat));
endmodule


