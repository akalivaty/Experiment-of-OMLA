//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 1 0 0 1 1 1 1 0 1 0 0 1 0 0 0 0 0 1 0 0 1 1 0 1 1 0 1 1 0 1 0 0 0 1 0 0 0 0 1 1 1 1 0 1 1 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:14 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078;
  INV_X1    g000(.A(G478), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(KEYINPUT15), .ZN(new_n188));
  INV_X1    g002(.A(G122), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G116), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G122), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  AND3_X1   g007(.A1(new_n190), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G128), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G143), .ZN(new_n199));
  INV_X1    g013(.A(G134), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n197), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n200), .B1(new_n197), .B2(new_n199), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n195), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT14), .ZN(new_n205));
  OAI21_X1  g019(.A(G107), .B1(new_n192), .B2(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(G116), .B(G122), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n206), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  OR2_X1    g022(.A1(new_n204), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT13), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT93), .B1(new_n197), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT93), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n212), .A2(new_n196), .A3(KEYINPUT13), .A4(G128), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n197), .A2(new_n210), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n211), .A2(new_n213), .A3(new_n199), .A4(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G134), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n207), .A2(new_n193), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n216), .B(new_n201), .C1(new_n217), .C2(new_n194), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT9), .B(G234), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n219), .B(KEYINPUT76), .ZN(new_n220));
  INV_X1    g034(.A(G953), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(G217), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n209), .A2(new_n218), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n201), .B1(new_n217), .B2(new_n194), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n225), .B1(G134), .B2(new_n215), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n204), .A2(new_n208), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n222), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT94), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n224), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT70), .B(G902), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n218), .A2(new_n209), .A3(KEYINPUT94), .A4(new_n223), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n188), .B1(new_n233), .B2(KEYINPUT95), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(KEYINPUT95), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT95), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n230), .A2(new_n232), .A3(new_n236), .A4(new_n231), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n234), .B1(new_n238), .B2(new_n188), .ZN(new_n239));
  OR2_X1    g053(.A1(KEYINPUT96), .A2(G952), .ZN(new_n240));
  NAND2_X1  g054(.A1(KEYINPUT96), .A2(G952), .ZN(new_n241));
  AOI21_X1  g055(.A(G953), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G234), .ZN(new_n243));
  INV_X1    g057(.A(G237), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  AOI211_X1 g060(.A(new_n221), .B(new_n231), .C1(G234), .C2(G237), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT21), .B(G898), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n239), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(G237), .A2(G953), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(G143), .A3(G214), .ZN(new_n253));
  INV_X1    g067(.A(G131), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(G143), .B1(new_n252), .B2(G214), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT87), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n253), .ZN(new_n258));
  OAI21_X1  g072(.A(G131), .B1(new_n258), .B2(new_n256), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n252), .A2(G214), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(new_n196), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT87), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n261), .A2(new_n262), .A3(new_n254), .A4(new_n253), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT17), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n257), .A2(new_n259), .A3(new_n263), .A4(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT16), .ZN(new_n266));
  INV_X1    g080(.A(G140), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(new_n267), .A3(G125), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(G125), .ZN(new_n269));
  INV_X1    g083(.A(G125), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G140), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n268), .B1(new_n272), .B2(new_n266), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT72), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n273), .A2(new_n274), .A3(G146), .ZN(new_n275));
  NOR3_X1   g089(.A1(new_n270), .A2(KEYINPUT16), .A3(G140), .ZN(new_n276));
  XNOR2_X1  g090(.A(G125), .B(G140), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n276), .B1(new_n277), .B2(KEYINPUT16), .ZN(new_n278));
  INV_X1    g092(.A(G146), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT72), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n274), .A2(G146), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n278), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n275), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n261), .A2(new_n253), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(KEYINPUT17), .A3(G131), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n265), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(G113), .B(G122), .ZN(new_n287));
  INV_X1    g101(.A(G104), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n287), .B(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT89), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n289), .B(new_n290), .ZN(new_n291));
  AND2_X1   g105(.A1(KEYINPUT64), .A2(G146), .ZN(new_n292));
  NOR2_X1   g106(.A1(KEYINPUT64), .A2(G146), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n277), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n295), .B1(new_n279), .B2(new_n277), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT18), .ZN(new_n297));
  NOR3_X1   g111(.A1(new_n284), .A2(new_n297), .A3(new_n254), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n261), .A2(new_n253), .B1(KEYINPUT18), .B2(G131), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n296), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AND3_X1   g114(.A1(new_n286), .A2(new_n291), .A3(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n257), .A2(new_n259), .A3(new_n263), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n278), .A2(G146), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT19), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n272), .A2(KEYINPUT88), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT88), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT19), .B1(new_n277), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n294), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n302), .A2(new_n303), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n289), .B1(new_n309), .B2(new_n300), .ZN(new_n310));
  OAI21_X1  g124(.A(KEYINPUT90), .B1(new_n301), .B2(new_n310), .ZN(new_n311));
  NOR2_X1   g125(.A1(G475), .A2(G902), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n309), .A2(new_n300), .ZN(new_n313));
  INV_X1    g127(.A(new_n289), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT90), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n286), .A2(new_n291), .A3(new_n300), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n311), .A2(new_n312), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT20), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n315), .A2(new_n317), .ZN(new_n321));
  NOR3_X1   g135(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT92), .ZN(new_n325));
  INV_X1    g139(.A(G902), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n289), .B1(new_n286), .B2(new_n300), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n326), .B1(new_n301), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT91), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT91), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n330), .B(new_n326), .C1(new_n301), .C2(new_n327), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n329), .A2(G475), .A3(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n324), .A2(new_n325), .A3(new_n332), .ZN(new_n333));
  AOI22_X1  g147(.A1(new_n319), .A2(KEYINPUT20), .B1(new_n321), .B2(new_n322), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n329), .A2(G475), .A3(new_n331), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT92), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n251), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  OR2_X1    g151(.A1(KEYINPUT0), .A2(G128), .ZN(new_n338));
  NAND2_X1  g152(.A1(KEYINPUT0), .A2(G128), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n196), .B1(new_n292), .B2(new_n293), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n279), .A2(G143), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT64), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n279), .ZN(new_n345));
  NAND2_X1  g159(.A1(KEYINPUT64), .A2(G146), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n345), .A2(KEYINPUT65), .A3(G143), .A4(new_n346), .ZN(new_n347));
  NOR3_X1   g161(.A1(new_n292), .A2(new_n293), .A3(new_n196), .ZN(new_n348));
  AOI21_X1  g162(.A(KEYINPUT65), .B1(new_n196), .B2(G146), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n347), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n339), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n343), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT82), .B1(new_n353), .B2(new_n270), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT1), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G128), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n351), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(G128), .B1(new_n348), .B2(new_n355), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n341), .A2(new_n342), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n358), .A2(new_n361), .A3(new_n270), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT82), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n345), .A2(G143), .A3(new_n346), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n349), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n339), .B1(new_n365), .B2(new_n347), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n363), .B(G125), .C1(new_n366), .C2(new_n343), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n221), .A2(G224), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n368), .B(KEYINPUT83), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT7), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n354), .A2(new_n362), .A3(new_n367), .A4(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT68), .ZN(new_n373));
  INV_X1    g187(.A(G119), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G116), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n191), .A2(G119), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n373), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(G116), .B(G119), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n373), .ZN(new_n380));
  XNOR2_X1  g194(.A(KEYINPUT2), .B(G113), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n378), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n375), .A2(new_n376), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n383), .A2(new_n381), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(KEYINPUT3), .B1(new_n288), .B2(G107), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT3), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(new_n193), .A3(G104), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n288), .A2(G107), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n387), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT4), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n392), .A3(G101), .ZN(new_n393));
  INV_X1    g207(.A(G101), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n387), .A2(new_n389), .A3(new_n394), .A4(new_n390), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n395), .B(KEYINPUT77), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n392), .B1(new_n391), .B2(G101), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n386), .B(new_n393), .C1(new_n396), .C2(new_n398), .ZN(new_n399));
  NOR3_X1   g213(.A1(new_n288), .A2(KEYINPUT3), .A3(G107), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n193), .A2(G104), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n402), .A2(KEYINPUT77), .A3(new_n394), .A4(new_n387), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT77), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n395), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(G104), .B(G107), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT78), .B1(new_n406), .B2(new_n394), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT78), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n288), .A2(G107), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n408), .B(G101), .C1(new_n409), .C2(new_n401), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n403), .A2(new_n405), .B1(new_n407), .B2(new_n410), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n375), .A2(new_n376), .A3(new_n373), .ZN(new_n412));
  OAI21_X1  g226(.A(KEYINPUT5), .B1(new_n412), .B2(new_n377), .ZN(new_n413));
  OAI21_X1  g227(.A(G113), .B1(new_n375), .B2(KEYINPUT5), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n384), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n411), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(G110), .B(G122), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n399), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n364), .A2(KEYINPUT1), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n420), .A2(G128), .B1(new_n342), .B2(new_n341), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n356), .B1(new_n365), .B2(new_n347), .ZN(new_n422));
  NOR3_X1   g236(.A1(new_n421), .A2(new_n422), .A3(G125), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n351), .A2(new_n352), .ZN(new_n424));
  INV_X1    g238(.A(new_n343), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n270), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n370), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n407), .A2(new_n410), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n395), .A2(new_n404), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n395), .A2(new_n404), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n416), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n379), .A2(KEYINPUT5), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n385), .B1(new_n433), .B2(new_n414), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n411), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n418), .B(KEYINPUT8), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n432), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n372), .A2(new_n419), .A3(new_n427), .A4(new_n437), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n438), .A2(KEYINPUT85), .A3(new_n326), .ZN(new_n439));
  AOI21_X1  g253(.A(KEYINPUT85), .B1(new_n438), .B2(new_n326), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT6), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n418), .B(KEYINPUT81), .ZN(new_n443));
  AOI211_X1 g257(.A(new_n442), .B(new_n443), .C1(new_n399), .C2(new_n417), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n399), .A2(new_n417), .ZN(new_n445));
  INV_X1    g259(.A(new_n443), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n419), .A2(KEYINPUT6), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n444), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT84), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n354), .A2(new_n362), .A3(new_n367), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n369), .ZN(new_n452));
  INV_X1    g266(.A(new_n369), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n354), .A2(new_n453), .A3(new_n362), .A4(new_n367), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NOR3_X1   g269(.A1(new_n449), .A2(new_n450), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n445), .A2(KEYINPUT6), .A3(new_n446), .ZN(new_n457));
  INV_X1    g271(.A(new_n393), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n403), .A2(new_n405), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n458), .B1(new_n459), .B2(new_n397), .ZN(new_n460));
  AOI22_X1  g274(.A1(new_n460), .A2(new_n386), .B1(new_n411), .B2(new_n416), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n442), .B1(new_n461), .B2(new_n418), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n461), .A2(new_n443), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n457), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n455), .ZN(new_n465));
  AOI21_X1  g279(.A(KEYINPUT84), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n441), .B1(new_n456), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(G210), .B1(G237), .B2(G902), .ZN(new_n468));
  XOR2_X1   g282(.A(new_n468), .B(KEYINPUT86), .Z(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(G214), .B1(G237), .B2(G902), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n441), .B(new_n469), .C1(new_n456), .C2(new_n466), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n337), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT10), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n342), .A2(KEYINPUT1), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(G128), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n365), .A2(new_n347), .A3(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n479), .A2(new_n422), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n476), .B1(new_n480), .B2(new_n431), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT11), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n482), .B1(new_n200), .B2(G137), .ZN(new_n483));
  INV_X1    g297(.A(G137), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n484), .A2(KEYINPUT11), .A3(G134), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n200), .A2(G137), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n483), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(G131), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n483), .A2(new_n485), .A3(new_n254), .A4(new_n486), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n358), .A2(new_n361), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(KEYINPUT10), .A3(new_n411), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n353), .B(new_n393), .C1(new_n396), .C2(new_n398), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n481), .A2(new_n491), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(G110), .B(G140), .ZN(new_n496));
  INV_X1    g310(.A(G227), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n497), .A2(G953), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n496), .B(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT79), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n481), .A2(new_n494), .A3(new_n493), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n490), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT79), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n495), .A2(new_n505), .A3(new_n500), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n502), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n411), .B1(new_n422), .B2(new_n479), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n421), .A2(new_n422), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n431), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(KEYINPUT12), .B1(new_n511), .B2(new_n490), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT12), .ZN(new_n513));
  AOI211_X1 g327(.A(new_n513), .B(new_n491), .C1(new_n508), .C2(new_n510), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n495), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n499), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n507), .A2(new_n516), .A3(G469), .ZN(new_n517));
  INV_X1    g331(.A(G469), .ZN(new_n518));
  INV_X1    g332(.A(new_n514), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n511), .A2(new_n490), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n513), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n501), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n500), .B1(new_n504), .B2(new_n495), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n518), .B(new_n231), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n518), .A2(new_n326), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n517), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(G221), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n528), .B1(new_n220), .B2(new_n326), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT80), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n527), .A2(KEYINPUT80), .A3(new_n530), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n475), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(G217), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n537), .B1(new_n231), .B2(G234), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT71), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n540), .B1(new_n374), .B2(G128), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n198), .A2(KEYINPUT71), .A3(G119), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n374), .A2(G128), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT24), .B(G110), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT73), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT23), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n548), .B1(new_n374), .B2(G128), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n198), .A2(KEYINPUT23), .A3(G119), .ZN(new_n550));
  INV_X1    g364(.A(G110), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n549), .A2(new_n550), .A3(new_n551), .A4(new_n543), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n546), .A2(new_n547), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n303), .A2(new_n295), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n547), .B1(new_n546), .B2(new_n552), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n544), .ZN(new_n558));
  INV_X1    g372(.A(new_n545), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n549), .A2(new_n543), .A3(new_n550), .ZN(new_n560));
  AOI22_X1  g374(.A1(new_n558), .A2(new_n559), .B1(new_n560), .B2(G110), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n561), .A2(new_n275), .A3(new_n282), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(KEYINPUT74), .B1(new_n557), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT74), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n546), .A2(new_n552), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT73), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(new_n295), .A3(new_n303), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n565), .B(new_n562), .C1(new_n568), .C2(new_n554), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT22), .B(G137), .ZN(new_n570));
  NOR3_X1   g384(.A1(new_n528), .A2(new_n243), .A3(G953), .ZN(new_n571));
  XOR2_X1   g385(.A(new_n570), .B(new_n571), .Z(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n564), .A2(new_n569), .A3(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n562), .B1(new_n568), .B2(new_n554), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n575), .A2(KEYINPUT74), .A3(new_n572), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n231), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT25), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n577), .A2(KEYINPUT25), .A3(new_n231), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n539), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n538), .A2(G902), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n577), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n486), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n200), .A2(G137), .ZN(new_n587));
  OAI21_X1  g401(.A(G131), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n588), .A2(new_n489), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n589), .B1(new_n421), .B2(new_n422), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(KEYINPUT67), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT67), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n592), .B(new_n589), .C1(new_n421), .C2(new_n422), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n353), .A2(KEYINPUT66), .A3(new_n490), .ZN(new_n594));
  AOI21_X1  g408(.A(KEYINPUT66), .B1(new_n353), .B2(new_n490), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n591), .B(new_n593), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n596), .A2(KEYINPUT69), .A3(new_n386), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n353), .A2(new_n490), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n590), .ZN(new_n599));
  OR2_X1    g413(.A1(new_n599), .A2(new_n386), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(KEYINPUT69), .B1(new_n596), .B2(new_n386), .ZN(new_n602));
  OAI21_X1  g416(.A(KEYINPUT28), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT28), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n252), .A2(G210), .ZN(new_n607));
  XOR2_X1   g421(.A(new_n607), .B(KEYINPUT27), .Z(new_n608));
  XNOR2_X1  g422(.A(KEYINPUT26), .B(G101), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT30), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n596), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n599), .A2(new_n611), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n612), .A2(new_n386), .A3(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n610), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(new_n600), .A3(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT31), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n599), .A2(new_n386), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n613), .B1(new_n596), .B2(new_n611), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n620), .B1(new_n621), .B2(new_n386), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n622), .A2(KEYINPUT31), .A3(new_n616), .ZN(new_n623));
  AOI22_X1  g437(.A1(new_n606), .A2(new_n610), .B1(new_n619), .B2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(G472), .A2(G902), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT32), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n620), .A2(KEYINPUT28), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n630), .A2(new_n610), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(KEYINPUT29), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n599), .A2(new_n386), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n604), .B1(new_n600), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n231), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n603), .A2(new_n631), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n615), .A2(new_n600), .ZN(new_n637));
  AOI21_X1  g451(.A(KEYINPUT29), .B1(new_n637), .B2(new_n610), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n635), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(G472), .ZN(new_n640));
  OAI22_X1  g454(.A1(new_n624), .A2(new_n629), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n596), .A2(new_n386), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT69), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n644), .A2(new_n600), .A3(new_n597), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n630), .B1(new_n645), .B2(KEYINPUT28), .ZN(new_n646));
  AND4_X1   g460(.A1(KEYINPUT31), .A2(new_n615), .A3(new_n600), .A4(new_n616), .ZN(new_n647));
  AOI21_X1  g461(.A(KEYINPUT31), .B1(new_n622), .B2(new_n616), .ZN(new_n648));
  OAI22_X1  g462(.A1(new_n646), .A2(new_n616), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(KEYINPUT32), .B1(new_n649), .B2(new_n625), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n585), .B1(new_n641), .B2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT75), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n231), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n605), .A2(new_n616), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT29), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n634), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n654), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n655), .B1(new_n645), .B2(KEYINPUT28), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n656), .B1(new_n622), .B2(new_n616), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  AOI22_X1  g476(.A1(new_n649), .A2(new_n628), .B1(new_n662), .B2(G472), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n627), .B1(new_n624), .B2(new_n626), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n665), .A2(KEYINPUT75), .A3(new_n585), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n536), .B1(new_n653), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(new_n394), .ZN(G3));
  AOI21_X1  g482(.A(new_n640), .B1(new_n649), .B2(new_n231), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT97), .ZN(new_n670));
  AOI22_X1  g484(.A1(new_n669), .A2(new_n670), .B1(new_n625), .B2(new_n649), .ZN(new_n671));
  INV_X1    g485(.A(new_n585), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n672), .B1(new_n533), .B2(new_n534), .ZN(new_n673));
  OAI21_X1  g487(.A(G472), .B1(new_n624), .B2(new_n654), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(KEYINPUT97), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n671), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n676), .B(KEYINPUT98), .Z(new_n677));
  AOI21_X1  g491(.A(new_n223), .B1(new_n209), .B2(new_n218), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT100), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n678), .B1(new_n679), .B2(new_n224), .ZN(new_n680));
  AOI211_X1 g494(.A(KEYINPUT100), .B(new_n223), .C1(new_n218), .C2(new_n209), .ZN(new_n681));
  OAI21_X1  g495(.A(KEYINPUT33), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n230), .A2(new_n232), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT33), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n654), .A2(new_n187), .ZN(new_n687));
  AOI22_X1  g501(.A1(new_n686), .A2(new_n687), .B1(new_n187), .B2(new_n233), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n688), .B1(new_n336), .B2(new_n333), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT99), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n690), .B1(new_n471), .B2(new_n473), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n469), .A2(KEYINPUT99), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n472), .B1(new_n467), .B2(new_n693), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n691), .A2(new_n249), .A3(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n677), .A2(new_n689), .A3(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT34), .B(G104), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G6));
  INV_X1    g512(.A(KEYINPUT20), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n311), .A2(new_n318), .A3(new_n699), .A4(new_n312), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n320), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n332), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n702), .A2(new_n239), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n677), .A2(new_n695), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT101), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT102), .ZN(new_n706));
  XOR2_X1   g520(.A(KEYINPUT35), .B(G107), .Z(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G9));
  INV_X1    g522(.A(KEYINPUT103), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n573), .A2(KEYINPUT36), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n575), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n583), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n709), .B1(new_n582), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g528(.A(KEYINPUT25), .B1(new_n577), .B2(new_n231), .ZN(new_n715));
  AOI211_X1 g529(.A(new_n579), .B(new_n654), .C1(new_n574), .C2(new_n576), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n538), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(KEYINPUT103), .A3(new_n712), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n475), .A2(new_n535), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n649), .A2(new_n231), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n670), .A3(G472), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n649), .A2(new_n625), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n675), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(KEYINPUT37), .B(G110), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(G12));
  INV_X1    g541(.A(G900), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n246), .B1(new_n247), .B2(new_n728), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n702), .A2(new_n239), .A3(new_n729), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n719), .B(new_n730), .C1(new_n641), .C2(new_n650), .ZN(new_n731));
  INV_X1    g545(.A(new_n473), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n450), .B1(new_n449), .B2(new_n455), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n464), .A2(KEYINPUT84), .A3(new_n465), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n469), .B1(new_n735), .B2(new_n441), .ZN(new_n736));
  OAI21_X1  g550(.A(KEYINPUT99), .B1(new_n732), .B2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n694), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n527), .A2(KEYINPUT80), .A3(new_n530), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT80), .B1(new_n527), .B2(new_n530), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n737), .B(new_n738), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n731), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g556(.A(KEYINPUT104), .B(G128), .Z(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G30));
  XOR2_X1   g558(.A(new_n729), .B(KEYINPUT39), .Z(new_n745));
  NAND2_X1  g559(.A1(new_n535), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(KEYINPUT106), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  OR2_X1    g562(.A1(new_n748), .A2(KEYINPUT40), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(KEYINPUT40), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n471), .A2(new_n473), .ZN(new_n751));
  XOR2_X1   g565(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n752));
  XNOR2_X1  g566(.A(new_n751), .B(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n617), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n616), .B1(new_n600), .B2(new_n633), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n326), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(G472), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n757), .B1(new_n624), .B2(new_n629), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n758), .A2(new_n650), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n239), .B1(new_n336), .B2(new_n333), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n760), .A2(new_n472), .A3(new_n714), .A4(new_n718), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n753), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n749), .A2(new_n750), .A3(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G143), .ZN(G45));
  INV_X1    g578(.A(new_n741), .ZN(new_n765));
  AOI22_X1  g579(.A1(new_n663), .A2(new_n664), .B1(new_n714), .B2(new_n718), .ZN(new_n766));
  AOI211_X1 g580(.A(new_n688), .B(new_n729), .C1(new_n336), .C2(new_n333), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n765), .A2(KEYINPUT107), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT107), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n767), .B(new_n719), .C1(new_n641), .C2(new_n650), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n769), .B1(new_n770), .B2(new_n741), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G146), .ZN(G48));
  NOR2_X1   g587(.A1(new_n522), .A2(new_n523), .ZN(new_n774));
  OAI21_X1  g588(.A(G469), .B1(new_n774), .B2(new_n654), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(new_n530), .A3(new_n524), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n585), .B(new_n777), .C1(new_n641), .C2(new_n650), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n737), .A2(new_n738), .A3(new_n250), .A4(new_n689), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  XOR2_X1   g594(.A(KEYINPUT41), .B(G113), .Z(new_n781));
  XNOR2_X1  g595(.A(new_n780), .B(new_n781), .ZN(G15));
  AOI21_X1  g596(.A(new_n672), .B1(new_n663), .B2(new_n664), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n783), .A2(new_n695), .A3(new_n703), .A4(new_n777), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G116), .ZN(G18));
  INV_X1    g599(.A(new_n337), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n786), .B(new_n719), .C1(new_n641), .C2(new_n650), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n737), .A2(new_n738), .A3(new_n777), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(new_n374), .ZN(G21));
  AND2_X1   g604(.A1(new_n777), .A2(new_n760), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n619), .A2(new_n623), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n610), .B1(new_n634), .B2(new_n630), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n626), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n794), .B1(new_n721), .B2(G472), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n791), .A2(new_n795), .A3(new_n585), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n737), .A2(new_n250), .A3(new_n738), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(new_n189), .ZN(G24));
  INV_X1    g613(.A(new_n794), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n767), .A2(new_n674), .A3(new_n719), .A4(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(KEYINPUT108), .B1(new_n801), .B2(new_n788), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n674), .A2(new_n719), .A3(new_n800), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT108), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n691), .A2(new_n694), .A3(new_n776), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n803), .A2(new_n804), .A3(new_n805), .A4(new_n767), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G125), .ZN(G27));
  INV_X1    g622(.A(KEYINPUT110), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n651), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n665), .A2(KEYINPUT110), .A3(new_n585), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n527), .A2(KEYINPUT109), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT109), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n517), .A2(new_n524), .A3(new_n813), .A4(new_n526), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n812), .A2(new_n530), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n336), .A2(new_n333), .ZN(new_n816));
  INV_X1    g630(.A(new_n688), .ZN(new_n817));
  INV_X1    g631(.A(new_n729), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n472), .B1(new_n732), .B2(new_n736), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n815), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n810), .A2(new_n811), .A3(KEYINPUT42), .A4(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n815), .A2(new_n820), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n783), .A2(new_n767), .A3(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT42), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(G131), .ZN(G33));
  AND3_X1   g642(.A1(new_n783), .A2(new_n730), .A3(new_n823), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(new_n200), .ZN(G36));
  NOR2_X1   g644(.A1(new_n816), .A2(new_n688), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT43), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n832), .A2(new_n719), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n724), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT44), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n472), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n837), .B1(new_n471), .B2(new_n473), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n833), .A2(KEYINPUT44), .A3(new_n724), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n836), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT45), .B1(new_n507), .B2(new_n516), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n518), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n507), .A2(new_n516), .A3(KEYINPUT45), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n526), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT46), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n524), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT111), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI211_X1 g663(.A(KEYINPUT111), .B(new_n524), .C1(new_n845), .C2(new_n846), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT112), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n845), .A2(new_n851), .A3(new_n846), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n845), .A2(new_n846), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT112), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n849), .A2(new_n850), .A3(new_n852), .A4(new_n854), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n855), .A2(new_n530), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n745), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n840), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(new_n484), .ZN(G39));
  AND3_X1   g673(.A1(new_n855), .A2(KEYINPUT47), .A3(new_n530), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT47), .B1(new_n855), .B2(new_n530), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n767), .A2(new_n838), .ZN(new_n863));
  NOR4_X1   g677(.A1(new_n862), .A2(new_n665), .A3(new_n585), .A4(new_n863), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(new_n267), .ZN(G42));
  NAND2_X1  g679(.A1(new_n775), .A2(new_n524), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n866), .A2(KEYINPUT49), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n585), .A2(new_n530), .A3(new_n472), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n866), .A2(KEYINPUT49), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n870), .A2(new_n753), .A3(new_n759), .A4(new_n831), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT118), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n829), .B1(new_n822), .B2(new_n826), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n471), .A2(new_n472), .A3(new_n473), .A4(new_n250), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n816), .A2(new_n817), .ZN(new_n876));
  INV_X1    g690(.A(new_n239), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n336), .A2(new_n333), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n875), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n671), .A2(new_n879), .A3(new_n673), .A4(new_n675), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(new_n784), .ZN(new_n881));
  OAI22_X1  g695(.A1(new_n720), .A2(new_n724), .B1(new_n778), .B2(new_n779), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OAI22_X1  g697(.A1(new_n796), .A2(new_n797), .B1(new_n787), .B2(new_n788), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n667), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n239), .A2(new_n701), .A3(new_n332), .A4(new_n818), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n717), .A2(KEYINPUT103), .A3(new_n712), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT103), .B1(new_n717), .B2(new_n712), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n890), .B1(new_n664), .B2(new_n663), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT113), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n891), .A2(new_n892), .A3(new_n535), .A4(new_n838), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n886), .B1(new_n714), .B2(new_n718), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n894), .B(new_n838), .C1(new_n641), .C2(new_n650), .ZN(new_n895));
  INV_X1    g709(.A(new_n535), .ZN(new_n896));
  OAI21_X1  g710(.A(KEYINPUT113), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI22_X1  g711(.A1(new_n893), .A2(new_n897), .B1(new_n803), .B2(new_n821), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n874), .A2(new_n883), .A3(new_n885), .A4(new_n898), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n582), .A2(new_n713), .A3(new_n729), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n900), .B1(new_n758), .B2(new_n650), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n737), .A2(new_n738), .A3(new_n760), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n901), .A2(new_n902), .A3(new_n815), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n903), .A2(new_n742), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n772), .A2(new_n904), .A3(new_n807), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT52), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n772), .A2(new_n904), .A3(KEYINPUT52), .A4(new_n807), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n899), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  XOR2_X1   g723(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n873), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(KEYINPUT52), .B1(new_n905), .B2(KEYINPUT114), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  AND4_X1   g728(.A1(new_n874), .A2(new_n883), .A3(new_n885), .A4(new_n898), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n905), .A2(KEYINPUT114), .A3(KEYINPUT52), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n914), .A2(KEYINPUT53), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n812), .A2(new_n530), .A3(new_n814), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n918), .B(new_n900), .C1(new_n650), .C2(new_n758), .ZN(new_n919));
  OAI22_X1  g733(.A1(new_n919), .A2(new_n902), .B1(new_n731), .B2(new_n741), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n920), .B1(new_n771), .B2(new_n768), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT52), .B1(new_n921), .B2(new_n807), .ZN(new_n922));
  AND4_X1   g736(.A1(KEYINPUT52), .A2(new_n772), .A3(new_n807), .A4(new_n904), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI211_X1 g738(.A(KEYINPUT118), .B(new_n910), .C1(new_n924), .C2(new_n899), .ZN(new_n925));
  AND4_X1   g739(.A1(new_n872), .A2(new_n912), .A3(new_n917), .A4(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n907), .A2(new_n908), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n927), .A2(new_n911), .A3(new_n915), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT117), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n909), .A2(KEYINPUT117), .A3(new_n911), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n905), .A2(KEYINPUT114), .A3(KEYINPUT52), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n933), .A2(new_n913), .A3(new_n899), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n934), .A2(KEYINPUT115), .A3(KEYINPUT53), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT115), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT53), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n932), .B1(new_n935), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n926), .B1(new_n940), .B2(KEYINPUT54), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n810), .A2(new_n811), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n820), .A2(new_n245), .A3(new_n776), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n942), .A2(new_n832), .A3(new_n943), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT48), .ZN(new_n945));
  NOR4_X1   g759(.A1(new_n669), .A2(new_n672), .A3(new_n245), .A4(new_n794), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n832), .A2(new_n805), .A3(new_n946), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n943), .A2(new_n585), .A3(new_n759), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(new_n689), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n945), .A2(new_n242), .A3(new_n947), .A4(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n776), .A2(new_n472), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n832), .A2(new_n946), .A3(new_n753), .A4(new_n951), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n952), .A2(KEYINPUT119), .A3(KEYINPUT50), .ZN(new_n953));
  AOI21_X1  g767(.A(KEYINPUT50), .B1(new_n952), .B2(KEYINPUT119), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n832), .A2(new_n803), .A3(new_n943), .ZN(new_n955));
  INV_X1    g769(.A(new_n948), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n336), .A2(new_n333), .A3(new_n688), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n953), .A2(new_n954), .A3(new_n958), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n866), .A2(new_n530), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n860), .A2(new_n861), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n832), .A2(new_n838), .A3(new_n946), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(KEYINPUT51), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT51), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n959), .B(new_n965), .C1(new_n961), .C2(new_n962), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n950), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT120), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n941), .A2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(G952), .A2(G953), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n871), .B1(new_n971), .B2(new_n972), .ZN(G75));
  XNOR2_X1  g787(.A(new_n464), .B(new_n465), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT55), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n911), .B1(new_n927), .B2(new_n915), .ZN(new_n977));
  AOI22_X1  g791(.A1(KEYINPUT53), .A2(new_n934), .B1(new_n977), .B2(KEYINPUT118), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n231), .B1(new_n978), .B2(new_n912), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(new_n469), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT56), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n976), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  AOI211_X1 g796(.A(KEYINPUT56), .B(new_n975), .C1(new_n979), .C2(new_n469), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n221), .A2(G952), .ZN(new_n984));
  NOR3_X1   g798(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(G51));
  XNOR2_X1  g799(.A(new_n525), .B(KEYINPUT57), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n872), .B1(new_n978), .B2(new_n912), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n986), .B1(new_n987), .B2(new_n926), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n774), .B(KEYINPUT121), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n979), .A2(new_n843), .A3(new_n842), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n984), .B1(new_n990), .B2(new_n991), .ZN(G54));
  NAND3_X1  g806(.A1(new_n979), .A2(KEYINPUT58), .A3(G475), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n311), .A2(new_n318), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n993), .A2(new_n994), .ZN(new_n996));
  NOR3_X1   g810(.A1(new_n995), .A2(new_n996), .A3(new_n984), .ZN(G60));
  INV_X1    g811(.A(new_n686), .ZN(new_n998));
  NAND2_X1  g812(.A1(G478), .A2(G902), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT59), .Z(new_n1000));
  OAI21_X1  g814(.A(new_n998), .B1(new_n941), .B2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n998), .A2(new_n1000), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1002), .B1(new_n987), .B2(new_n926), .ZN(new_n1003));
  INV_X1    g817(.A(new_n984), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n1003), .A2(KEYINPUT122), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT122), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1002), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n925), .A2(new_n917), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n977), .A2(KEYINPUT118), .ZN(new_n1009));
  OAI21_X1  g823(.A(KEYINPUT54), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n912), .A2(new_n925), .A3(new_n872), .A4(new_n917), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1007), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1006), .B1(new_n1012), .B2(new_n984), .ZN(new_n1013));
  AND3_X1   g827(.A1(new_n1001), .A2(new_n1005), .A3(new_n1013), .ZN(G63));
  NAND2_X1  g828(.A1(G217), .A2(G902), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n1015), .B(KEYINPUT60), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1016), .ZN(new_n1017));
  OAI211_X1 g831(.A(new_n711), .B(new_n1017), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1018));
  AOI21_X1  g832(.A(KEYINPUT61), .B1(new_n1018), .B2(KEYINPUT123), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n978), .A2(new_n912), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n577), .B1(new_n1020), .B2(new_n1017), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1018), .A2(new_n1004), .ZN(new_n1022));
  OR3_X1    g836(.A1(new_n1019), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1019), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1023), .A2(new_n1024), .ZN(G66));
  INV_X1    g839(.A(G224), .ZN(new_n1026));
  OAI21_X1  g840(.A(G953), .B1(new_n248), .B2(new_n1026), .ZN(new_n1027));
  AND2_X1   g841(.A1(new_n883), .A2(new_n885), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1027), .B1(new_n1028), .B2(G953), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n449), .B1(G898), .B2(new_n221), .ZN(new_n1030));
  XNOR2_X1  g844(.A(new_n1029), .B(new_n1030), .ZN(G69));
  NOR2_X1   g845(.A1(new_n305), .A2(new_n307), .ZN(new_n1032));
  XNOR2_X1  g846(.A(new_n621), .B(new_n1032), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1033), .B1(new_n497), .B2(G953), .ZN(new_n1034));
  INV_X1    g848(.A(new_n858), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n742), .B1(new_n768), .B2(new_n771), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1036), .A2(new_n807), .ZN(new_n1037));
  INV_X1    g851(.A(new_n1037), .ZN(new_n1038));
  AOI21_X1  g852(.A(KEYINPUT126), .B1(new_n1035), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g853(.A(KEYINPUT126), .ZN(new_n1040));
  NOR3_X1   g854(.A1(new_n858), .A2(new_n1037), .A3(new_n1040), .ZN(new_n1041));
  NOR2_X1   g855(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g856(.A(new_n902), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n942), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g858(.A(new_n874), .B1(new_n857), .B2(new_n1044), .ZN(new_n1045));
  NOR3_X1   g859(.A1(new_n1042), .A2(new_n864), .A3(new_n1045), .ZN(new_n1046));
  OAI21_X1  g860(.A(new_n1034), .B1(new_n1046), .B2(G953), .ZN(new_n1047));
  AND2_X1   g861(.A1(new_n1033), .A2(new_n497), .ZN(new_n1048));
  OAI21_X1  g862(.A(G953), .B1(new_n1048), .B2(new_n728), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n653), .A2(new_n666), .ZN(new_n1050));
  AOI21_X1  g864(.A(new_n820), .B1(new_n876), .B2(new_n878), .ZN(new_n1051));
  NAND3_X1  g865(.A1(new_n747), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g866(.A(new_n1052), .B(KEYINPUT124), .ZN(new_n1053));
  OR3_X1    g867(.A1(new_n858), .A2(new_n1053), .A3(KEYINPUT125), .ZN(new_n1054));
  OAI21_X1  g868(.A(KEYINPUT125), .B1(new_n858), .B2(new_n1053), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g870(.A1(new_n763), .A2(new_n1038), .ZN(new_n1057));
  INV_X1    g871(.A(KEYINPUT62), .ZN(new_n1058));
  NAND2_X1  g872(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g873(.A1(new_n763), .A2(KEYINPUT62), .A3(new_n1038), .ZN(new_n1060));
  AOI21_X1  g874(.A(new_n864), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g875(.A1(new_n1056), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g876(.A1(new_n1062), .A2(new_n221), .A3(new_n1033), .ZN(new_n1063));
  NAND3_X1  g877(.A1(new_n1047), .A2(new_n1049), .A3(new_n1063), .ZN(G72));
  NAND3_X1  g878(.A1(new_n1056), .A2(new_n1061), .A3(new_n1028), .ZN(new_n1065));
  NAND2_X1  g879(.A1(G472), .A2(G902), .ZN(new_n1066));
  XOR2_X1   g880(.A(new_n1066), .B(KEYINPUT63), .Z(new_n1067));
  NAND2_X1  g881(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g882(.A(new_n637), .B(KEYINPUT127), .ZN(new_n1069));
  NAND3_X1  g883(.A1(new_n1068), .A2(new_n616), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g884(.A1(new_n637), .A2(new_n610), .ZN(new_n1071));
  NAND2_X1  g885(.A1(new_n1071), .A2(new_n617), .ZN(new_n1072));
  NAND3_X1  g886(.A1(new_n940), .A2(new_n1067), .A3(new_n1072), .ZN(new_n1073));
  NOR2_X1   g887(.A1(new_n864), .A2(new_n1045), .ZN(new_n1074));
  OAI211_X1 g888(.A(new_n1074), .B(new_n1028), .C1(new_n1039), .C2(new_n1041), .ZN(new_n1075));
  NAND2_X1  g889(.A1(new_n1075), .A2(new_n1067), .ZN(new_n1076));
  NOR2_X1   g890(.A1(new_n1069), .A2(new_n616), .ZN(new_n1077));
  AOI21_X1  g891(.A(new_n984), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  AND3_X1   g892(.A1(new_n1070), .A2(new_n1073), .A3(new_n1078), .ZN(G57));
endmodule


