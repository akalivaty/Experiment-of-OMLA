//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 0 0 0 1 0 1 0 1 0 1 1 1 0 1 0 0 0 0 1 1 0 0 1 1 0 1 1 0 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994;
  INV_X1    g000(.A(KEYINPUT15), .ZN(new_n187));
  AND2_X1   g001(.A1(new_n187), .A2(KEYINPUT97), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n187), .A2(KEYINPUT97), .ZN(new_n189));
  OAI21_X1  g003(.A(G478), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT9), .B(G234), .ZN(new_n191));
  INV_X1    g005(.A(G217), .ZN(new_n192));
  NOR3_X1   g006(.A1(new_n191), .A2(new_n192), .A3(G953), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G107), .ZN(new_n195));
  INV_X1    g009(.A(G116), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G122), .ZN(new_n197));
  XNOR2_X1  g011(.A(new_n197), .B(KEYINPUT95), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT96), .ZN(new_n199));
  AND2_X1   g013(.A1(KEYINPUT94), .A2(G122), .ZN(new_n200));
  NOR2_X1   g014(.A1(KEYINPUT94), .A2(G122), .ZN(new_n201));
  OAI21_X1  g015(.A(G116), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n198), .A2(new_n199), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n199), .B1(new_n198), .B2(new_n202), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n195), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n198), .A2(KEYINPUT14), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(new_n202), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n198), .A2(KEYINPUT14), .ZN(new_n209));
  OAI21_X1  g023(.A(G107), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G128), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(G143), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT65), .B(G128), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n212), .B1(new_n213), .B2(G143), .ZN(new_n214));
  INV_X1    g028(.A(G134), .ZN(new_n215));
  XNOR2_X1  g029(.A(new_n214), .B(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n206), .A2(new_n210), .A3(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n214), .A2(KEYINPUT13), .ZN(new_n219));
  INV_X1    g033(.A(new_n212), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n219), .B(G134), .C1(KEYINPUT13), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n214), .A2(new_n215), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n205), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n224), .A2(G107), .A3(new_n203), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n223), .B1(new_n206), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n194), .B1(new_n218), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n206), .A2(new_n225), .ZN(new_n228));
  INV_X1    g042(.A(new_n223), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n230), .A2(new_n217), .A3(new_n193), .ZN(new_n231));
  AOI21_X1  g045(.A(G902), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT98), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n190), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n233), .ZN(new_n235));
  XOR2_X1   g049(.A(new_n234), .B(new_n235), .Z(new_n236));
  INV_X1    g050(.A(G902), .ZN(new_n237));
  XNOR2_X1  g051(.A(G113), .B(G122), .ZN(new_n238));
  INV_X1    g052(.A(G104), .ZN(new_n239));
  XNOR2_X1  g053(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(G125), .B(G140), .ZN(new_n241));
  INV_X1    g055(.A(G146), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n243), .B(KEYINPUT90), .ZN(new_n244));
  INV_X1    g058(.A(G237), .ZN(new_n245));
  INV_X1    g059(.A(G953), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n245), .A2(new_n246), .A3(G214), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n247), .B(G143), .ZN(new_n248));
  INV_X1    g062(.A(G131), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT18), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT18), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n248), .B1(new_n252), .B2(new_n249), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n244), .A2(new_n251), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G140), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G125), .ZN(new_n256));
  INV_X1    g070(.A(G125), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G140), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n256), .A2(new_n258), .A3(KEYINPUT16), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT73), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT73), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n256), .A2(new_n258), .A3(new_n261), .A4(KEYINPUT16), .ZN(new_n262));
  OR3_X1    g076(.A1(new_n257), .A2(KEYINPUT16), .A3(G140), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n260), .A2(G146), .A3(new_n262), .A4(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT74), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n262), .A2(new_n263), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n267), .A2(KEYINPUT74), .A3(G146), .A4(new_n260), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n262), .A2(new_n263), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n261), .B1(new_n241), .B2(KEYINPUT16), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n242), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n266), .A2(new_n268), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT91), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n266), .A2(new_n268), .A3(KEYINPUT91), .A4(new_n271), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n250), .A2(KEYINPUT17), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n274), .A2(KEYINPUT92), .A3(new_n275), .A4(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n248), .B(new_n249), .ZN(new_n278));
  OR2_X1    g092(.A1(new_n278), .A2(KEYINPUT17), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n272), .A2(new_n273), .B1(KEYINPUT17), .B2(new_n250), .ZN(new_n281));
  AOI21_X1  g095(.A(KEYINPUT92), .B1(new_n281), .B2(new_n275), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n240), .B(new_n254), .C1(new_n280), .C2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT93), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT92), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(new_n277), .A3(new_n279), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n240), .B1(new_n289), .B2(new_n254), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n237), .B1(new_n285), .B2(new_n290), .ZN(new_n291));
  AOI211_X1 g105(.A(new_n284), .B(new_n240), .C1(new_n289), .C2(new_n254), .ZN(new_n292));
  OAI21_X1  g106(.A(G475), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  XOR2_X1   g107(.A(new_n241), .B(KEYINPUT19), .Z(new_n294));
  OAI211_X1 g108(.A(new_n278), .B(new_n264), .C1(G146), .C2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n254), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n240), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n283), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(G475), .A2(G902), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT20), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT20), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n299), .A2(new_n303), .A3(new_n300), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n236), .A2(new_n293), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n246), .A2(G952), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n307), .B1(G234), .B2(G237), .ZN(new_n308));
  NAND2_X1  g122(.A1(G234), .A2(G237), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(G902), .A3(G953), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT21), .B(G898), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n308), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n306), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT76), .B(KEYINPUT25), .ZN(new_n315));
  XOR2_X1   g129(.A(KEYINPUT22), .B(G137), .Z(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(KEYINPUT75), .ZN(new_n317));
  AND3_X1   g131(.A1(new_n246), .A2(G221), .A3(G234), .ZN(new_n318));
  XOR2_X1   g132(.A(new_n317), .B(new_n318), .Z(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G119), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G128), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT23), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n323), .B1(new_n321), .B2(G128), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n213), .A2(G119), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT23), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G110), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n325), .A2(new_n322), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT72), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT72), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n325), .A2(new_n331), .A3(new_n322), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT24), .B(G110), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n330), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n272), .A2(new_n328), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n241), .A2(new_n242), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n334), .B1(new_n330), .B2(new_n332), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n327), .A2(G110), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n264), .B(new_n337), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n320), .A2(new_n336), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n320), .B1(new_n336), .B2(new_n340), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI211_X1 g158(.A(KEYINPUT77), .B(new_n315), .C1(new_n344), .C2(G902), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT77), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n336), .A2(new_n340), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n319), .ZN(new_n348));
  AOI21_X1  g162(.A(G902), .B1(new_n348), .B2(new_n341), .ZN(new_n349));
  INV_X1    g163(.A(new_n315), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n346), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(KEYINPUT25), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n345), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n192), .B1(G234), .B2(new_n237), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n344), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n354), .A2(G902), .ZN(new_n357));
  XOR2_X1   g171(.A(new_n357), .B(KEYINPUT78), .Z(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT31), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT11), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n362), .B1(new_n215), .B2(G137), .ZN(new_n363));
  INV_X1    g177(.A(G137), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n364), .A2(KEYINPUT11), .A3(G134), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n215), .A2(G137), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n363), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G131), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n363), .A2(new_n365), .A3(new_n249), .A4(new_n366), .ZN(new_n369));
  INV_X1    g183(.A(G143), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n370), .A2(G146), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n242), .A2(G143), .ZN(new_n372));
  NOR2_X1   g186(.A1(KEYINPUT0), .A2(G128), .ZN(new_n373));
  AND2_X1   g187(.A1(KEYINPUT0), .A2(G128), .ZN(new_n374));
  OAI22_X1  g188(.A1(new_n371), .A2(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n242), .A2(G143), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n370), .A2(G146), .ZN(new_n377));
  NAND2_X1  g191(.A1(KEYINPUT0), .A2(G128), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  AOI22_X1  g193(.A1(new_n368), .A2(new_n369), .B1(new_n375), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n215), .A2(G137), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n364), .A2(G134), .ZN(new_n383));
  OAI21_X1  g197(.A(G131), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n369), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n376), .A2(new_n377), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT1), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n387), .B1(G143), .B2(new_n242), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n386), .B1(new_n213), .B2(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(G143), .B(G146), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(new_n387), .A3(G128), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n385), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n381), .A2(new_n393), .ZN(new_n394));
  XOR2_X1   g208(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n368), .A2(new_n369), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n374), .A2(new_n373), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n379), .B(KEYINPUT67), .C1(new_n398), .C2(new_n390), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(KEYINPUT67), .B1(new_n375), .B2(new_n379), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n397), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(KEYINPUT30), .A3(new_n393), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT2), .ZN(new_n404));
  INV_X1    g218(.A(G113), .ZN(new_n405));
  OAI21_X1  g219(.A(KEYINPUT66), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT66), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(KEYINPUT2), .A3(G113), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n404), .A2(new_n405), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(G116), .B(G119), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n409), .A2(new_n410), .A3(new_n412), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n396), .A2(new_n403), .A3(new_n416), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n409), .A2(new_n410), .A3(new_n412), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n412), .B1(new_n409), .B2(new_n410), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n402), .A2(new_n420), .A3(new_n393), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n417), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n245), .A2(new_n246), .A3(G210), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n423), .B(KEYINPUT27), .ZN(new_n424));
  XNOR2_X1  g238(.A(KEYINPUT26), .B(G101), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n424), .B(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n361), .B1(new_n422), .B2(new_n427), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n417), .A2(KEYINPUT31), .A3(new_n426), .A4(new_n421), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n369), .A2(new_n384), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n431), .B1(new_n389), .B2(new_n391), .ZN(new_n432));
  OAI211_X1 g246(.A(KEYINPUT68), .B(new_n416), .C1(new_n432), .C2(new_n380), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n421), .ZN(new_n434));
  AOI21_X1  g248(.A(KEYINPUT68), .B1(new_n394), .B2(new_n416), .ZN(new_n435));
  OAI21_X1  g249(.A(KEYINPUT28), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT28), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n421), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(KEYINPUT69), .B1(new_n440), .B2(new_n427), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT68), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n375), .A2(new_n379), .ZN(new_n443));
  AOI22_X1  g257(.A1(new_n397), .A2(new_n443), .B1(new_n385), .B2(new_n392), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n442), .B1(new_n444), .B2(new_n420), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n445), .A2(new_n421), .A3(new_n433), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n438), .B1(new_n446), .B2(KEYINPUT28), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT69), .ZN(new_n448));
  NOR3_X1   g262(.A1(new_n447), .A2(new_n448), .A3(new_n426), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n430), .B1(new_n441), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(G472), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n450), .A2(new_n451), .A3(new_n237), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT32), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n448), .B1(new_n447), .B2(new_n426), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n433), .A2(new_n421), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n437), .B1(new_n455), .B2(new_n445), .ZN(new_n456));
  OAI211_X1 g270(.A(KEYINPUT69), .B(new_n427), .C1(new_n456), .C2(new_n438), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(G902), .B1(new_n458), .B2(new_n430), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT32), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n460), .A3(new_n451), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n453), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT70), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n421), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n402), .A2(new_n393), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n416), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n466), .A2(KEYINPUT70), .ZN(new_n468));
  OAI21_X1  g282(.A(KEYINPUT28), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n426), .A2(KEYINPUT29), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n469), .A2(new_n439), .A3(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT71), .ZN(new_n472));
  OR2_X1    g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n426), .B1(new_n417), .B2(new_n421), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(KEYINPUT29), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n447), .A2(new_n426), .ZN(new_n476));
  AOI21_X1  g290(.A(G902), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n471), .A2(new_n472), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n473), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G472), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n360), .B1(new_n462), .B2(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(G110), .B(G122), .ZN(new_n482));
  OAI21_X1  g296(.A(KEYINPUT3), .B1(new_n239), .B2(G107), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT3), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n484), .A2(new_n195), .A3(G104), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n239), .A2(G107), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n483), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT4), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(new_n488), .A3(G101), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(G101), .ZN(new_n490));
  INV_X1    g304(.A(G101), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n483), .A2(new_n485), .A3(new_n491), .A4(new_n486), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n490), .A2(KEYINPUT4), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n416), .A2(new_n489), .A3(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n239), .A2(G107), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n195), .A2(G104), .ZN(new_n496));
  OAI21_X1  g310(.A(G101), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n321), .A2(G116), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT5), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n405), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n196), .A2(G119), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n500), .A2(new_n504), .A3(KEYINPUT5), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n499), .A2(new_n415), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n482), .B1(new_n494), .B2(new_n507), .ZN(new_n508));
  OR2_X1    g322(.A1(new_n508), .A2(KEYINPUT6), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n493), .A2(new_n489), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n507), .B(new_n482), .C1(new_n510), .C2(new_n420), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT84), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n494), .A2(KEYINPUT84), .A3(new_n507), .A4(new_n482), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n508), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT6), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n509), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n375), .A2(G125), .A3(new_n379), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n518), .B1(new_n392), .B2(G125), .ZN(new_n519));
  XOR2_X1   g333(.A(KEYINPUT85), .B(G224), .Z(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n246), .ZN(new_n521));
  XOR2_X1   g335(.A(new_n519), .B(new_n521), .Z(new_n522));
  NAND2_X1  g336(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT89), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT7), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n525), .B1(new_n520), .B2(new_n246), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT88), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n526), .B1(new_n518), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n519), .A2(new_n528), .ZN(new_n529));
  OAI221_X1 g343(.A(new_n518), .B1(new_n526), .B2(new_n527), .C1(new_n392), .C2(G125), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n506), .A2(new_n498), .A3(new_n415), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT86), .B(KEYINPUT8), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n482), .B(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT87), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n505), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n412), .A2(KEYINPUT87), .A3(KEYINPUT5), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(new_n538), .A3(new_n503), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n498), .B1(new_n539), .B2(new_n415), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n524), .B1(new_n531), .B2(new_n541), .ZN(new_n542));
  AND2_X1   g356(.A1(new_n539), .A2(new_n415), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n532), .B(new_n534), .C1(new_n543), .C2(new_n498), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n544), .A2(KEYINPUT89), .A3(new_n529), .A4(new_n530), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n513), .A2(new_n514), .ZN(new_n547));
  AOI21_X1  g361(.A(G902), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(G210), .B1(G237), .B2(G902), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n523), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n549), .B1(new_n523), .B2(new_n548), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(G214), .B1(G237), .B2(G902), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(KEYINPUT83), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(G221), .B1(new_n191), .B2(G902), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n376), .A2(KEYINPUT1), .ZN(new_n558));
  AOI22_X1  g372(.A1(new_n558), .A2(G128), .B1(new_n376), .B2(new_n377), .ZN(new_n559));
  AND4_X1   g373(.A1(new_n387), .A2(new_n376), .A3(new_n377), .A4(G128), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n492), .B(new_n497), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT10), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n562), .B1(new_n389), .B2(new_n391), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n561), .A2(new_n562), .B1(new_n563), .B2(new_n499), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n493), .B(new_n489), .C1(new_n400), .C2(new_n401), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(KEYINPUT80), .A3(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(KEYINPUT80), .B1(new_n564), .B2(new_n565), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n397), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n397), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n561), .A2(new_n562), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n563), .A2(new_n499), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n565), .A2(new_n570), .A3(new_n571), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(KEYINPUT79), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT79), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n564), .A2(new_n575), .A3(new_n565), .A4(new_n570), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n569), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(G110), .B(G140), .ZN(new_n579));
  INV_X1    g393(.A(G227), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(G953), .ZN(new_n581));
  XOR2_X1   g395(.A(new_n579), .B(new_n581), .Z(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT81), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n577), .A2(new_n585), .A3(new_n582), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n561), .B1(new_n392), .B2(new_n499), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n397), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT12), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n583), .B1(new_n574), .B2(new_n576), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n592), .A2(new_n585), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n584), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(G469), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n595), .A3(new_n237), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(KEYINPUT82), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n577), .A2(new_n582), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT81), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n588), .B(KEYINPUT12), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n592), .B2(new_n585), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(G902), .B1(new_n602), .B2(new_n584), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT82), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n603), .A2(new_n604), .A3(new_n595), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n597), .A2(new_n605), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n592), .A2(new_n569), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n582), .B1(new_n590), .B2(new_n577), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(G469), .B1(new_n609), .B2(G902), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n557), .B1(new_n606), .B2(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n314), .A2(new_n481), .A3(new_n555), .A4(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(G101), .ZN(G3));
  AOI22_X1  g427(.A1(new_n454), .A2(new_n457), .B1(new_n428), .B2(new_n429), .ZN(new_n614));
  OAI21_X1  g428(.A(G472), .B1(new_n614), .B2(G902), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n452), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n360), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n611), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n313), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n523), .A2(new_n548), .A3(new_n549), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n620), .B1(new_n551), .B2(KEYINPUT99), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT99), .ZN(new_n622));
  AOI211_X1 g436(.A(new_n622), .B(new_n549), .C1(new_n523), .C2(new_n548), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n619), .B(new_n553), .C1(new_n621), .C2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n218), .A2(new_n226), .A3(new_n194), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n193), .B1(new_n230), .B2(new_n217), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT100), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n628), .B1(new_n230), .B2(new_n217), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT33), .ZN(new_n630));
  OAI22_X1  g444(.A1(new_n626), .A2(new_n627), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(KEYINPUT100), .B1(new_n218), .B2(new_n226), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n227), .A2(new_n632), .A3(new_n231), .A4(KEYINPUT33), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n631), .A2(new_n633), .A3(new_n237), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(G478), .ZN(new_n635));
  INV_X1    g449(.A(G478), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n232), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n293), .B2(new_n305), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n625), .A2(KEYINPUT101), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(KEYINPUT101), .B1(new_n625), .B2(new_n639), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n618), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT34), .B(G104), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  XNOR2_X1  g458(.A(new_n234), .B(new_n235), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n293), .A2(new_n305), .A3(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n647), .A2(KEYINPUT102), .A3(new_n625), .ZN(new_n648));
  AOI21_X1  g462(.A(KEYINPUT102), .B1(new_n647), .B2(new_n625), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n618), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(new_n650), .B(KEYINPUT103), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT35), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G107), .ZN(G9));
  NOR2_X1   g467(.A1(new_n320), .A2(KEYINPUT36), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(new_n347), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n358), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n657), .B1(new_n353), .B2(new_n354), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n616), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n314), .A2(new_n659), .A3(new_n555), .A4(new_n611), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT37), .B(G110), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G12));
  AOI21_X1  g476(.A(new_n658), .B1(new_n462), .B2(new_n480), .ZN(new_n663));
  INV_X1    g477(.A(new_n308), .ZN(new_n664));
  INV_X1    g478(.A(G900), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n311), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n646), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n553), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n523), .A2(new_n548), .ZN(new_n671));
  INV_X1    g485(.A(new_n549), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n550), .B1(new_n673), .B2(new_n622), .ZN(new_n674));
  INV_X1    g488(.A(new_n623), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n670), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n663), .A2(new_n669), .A3(new_n611), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G128), .ZN(G30));
  XNOR2_X1  g492(.A(new_n667), .B(KEYINPUT39), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n611), .A2(new_n679), .ZN(new_n680));
  OR2_X1    g494(.A1(new_n680), .A2(KEYINPUT40), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n467), .A2(new_n468), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n682), .A2(new_n426), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n422), .A2(new_n427), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n237), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(G472), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n460), .B1(new_n459), .B2(new_n451), .ZN(new_n687));
  NOR4_X1   g501(.A1(new_n614), .A2(KEYINPUT32), .A3(G472), .A4(G902), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n686), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n552), .B(KEYINPUT38), .ZN(new_n691));
  INV_X1    g505(.A(new_n658), .ZN(new_n692));
  NOR4_X1   g506(.A1(new_n690), .A2(new_n691), .A3(new_n670), .A4(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n680), .A2(KEYINPUT40), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n289), .A2(new_n254), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n297), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n696), .A2(new_n284), .A3(new_n283), .ZN(new_n697));
  INV_X1    g511(.A(new_n292), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n697), .A2(new_n698), .A3(new_n237), .ZN(new_n699));
  AOI22_X1  g513(.A1(new_n699), .A2(G475), .B1(new_n302), .B2(new_n304), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n700), .A2(new_n236), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n681), .A2(new_n693), .A3(new_n694), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G143), .ZN(G45));
  AOI211_X1 g517(.A(new_n668), .B(new_n638), .C1(new_n293), .C2(new_n305), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n663), .A2(new_n704), .A3(new_n611), .A4(new_n676), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G146), .ZN(G48));
  AND3_X1   g520(.A1(new_n594), .A2(KEYINPUT104), .A3(new_n237), .ZN(new_n707));
  AOI21_X1  g521(.A(KEYINPUT104), .B1(new_n594), .B2(new_n237), .ZN(new_n708));
  OAI21_X1  g522(.A(G469), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n709), .A2(new_n606), .A3(new_n556), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  AND2_X1   g525(.A1(new_n711), .A2(new_n481), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n712), .B1(new_n640), .B2(new_n641), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT41), .B(G113), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G15));
  OAI21_X1  g529(.A(new_n712), .B1(new_n649), .B2(new_n648), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G116), .ZN(G18));
  NAND4_X1  g531(.A1(new_n676), .A2(new_n556), .A3(new_n606), .A4(new_n709), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n480), .B1(new_n687), .B2(new_n688), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n692), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n314), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G119), .ZN(G21));
  AOI22_X1  g537(.A1(new_n353), .A2(new_n354), .B1(new_n356), .B2(new_n358), .ZN(new_n724));
  NOR2_X1   g538(.A1(G472), .A2(G902), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(KEYINPUT105), .ZN(new_n726));
  INV_X1    g540(.A(new_n430), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n426), .B1(new_n469), .B2(new_n439), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n724), .A2(new_n615), .A3(new_n619), .A4(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n710), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n553), .B1(new_n621), .B2(new_n623), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n700), .A2(new_n732), .A3(new_n236), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G122), .ZN(G24));
  NAND2_X1  g549(.A1(new_n615), .A2(new_n729), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n658), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n711), .A2(new_n676), .A3(new_n704), .A4(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G125), .ZN(G27));
  NAND2_X1  g553(.A1(new_n673), .A2(new_n620), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n670), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n481), .A2(new_n704), .A3(new_n611), .A4(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT42), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n604), .B1(new_n603), .B2(new_n595), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n582), .B1(new_n569), .B2(new_n577), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n746), .B1(new_n599), .B2(new_n601), .ZN(new_n747));
  NOR4_X1   g561(.A1(new_n747), .A2(KEYINPUT82), .A3(G469), .A4(G902), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n610), .B1(new_n745), .B2(new_n748), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n749), .A2(new_n556), .A3(new_n741), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n750), .A2(KEYINPUT42), .A3(new_n481), .A4(new_n704), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n744), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G131), .ZN(G33));
  NAND3_X1  g567(.A1(new_n750), .A2(new_n481), .A3(new_n669), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G134), .ZN(G36));
  OR3_X1    g569(.A1(new_n607), .A2(new_n608), .A3(KEYINPUT45), .ZN(new_n756));
  OAI21_X1  g570(.A(KEYINPUT45), .B1(new_n607), .B2(new_n608), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n758), .A2(KEYINPUT106), .A3(G469), .ZN(new_n759));
  AOI21_X1  g573(.A(KEYINPUT106), .B1(new_n758), .B2(G469), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(G469), .A2(G902), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(KEYINPUT46), .A3(new_n762), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n762), .B1(new_n759), .B2(new_n760), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT46), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n763), .A2(new_n606), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n556), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n293), .A2(new_n305), .ZN(new_n770));
  OR3_X1    g584(.A1(new_n770), .A2(KEYINPUT43), .A3(new_n638), .ZN(new_n771));
  OAI21_X1  g585(.A(KEYINPUT43), .B1(new_n770), .B2(new_n638), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n658), .B1(new_n615), .B2(new_n452), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(KEYINPUT44), .A3(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n769), .A2(new_n679), .A3(new_n775), .A4(new_n741), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT44), .B1(new_n773), .B2(new_n774), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(new_n364), .ZN(G39));
  INV_X1    g593(.A(new_n741), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n719), .A2(new_n780), .A3(new_n724), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n767), .A2(KEYINPUT47), .A3(new_n556), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(KEYINPUT47), .B1(new_n767), .B2(new_n556), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n704), .B(new_n781), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT107), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n785), .B(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G140), .ZN(G42));
  OR2_X1    g602(.A1(G952), .A2(G953), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT119), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n360), .A2(new_n736), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n771), .A2(new_n308), .A3(new_n791), .A4(new_n772), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n711), .A2(new_n670), .A3(new_n691), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT50), .ZN(new_n794));
  OR3_X1    g608(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n794), .B1(new_n792), .B2(new_n793), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n690), .A2(new_n724), .A3(new_n308), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n710), .A2(new_n780), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT115), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n799), .A2(new_n803), .A3(new_n800), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n802), .A2(new_n700), .A3(new_n638), .A4(new_n804), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n773), .A2(new_n308), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(new_n737), .A3(new_n800), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n797), .A2(new_n805), .A3(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n792), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n809), .A2(KEYINPUT113), .A3(new_n741), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT113), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n811), .B1(new_n792), .B2(new_n780), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n784), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n782), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n709), .A2(new_n606), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n817), .A2(new_n556), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n814), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n808), .A2(new_n819), .A3(KEYINPUT51), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT116), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n808), .A2(new_n819), .A3(KEYINPUT116), .A4(KEYINPUT51), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n802), .A2(new_n639), .A3(new_n804), .ZN(new_n825));
  XOR2_X1   g639(.A(new_n307), .B(KEYINPUT117), .Z(new_n826));
  OAI211_X1 g640(.A(new_n825), .B(new_n826), .C1(new_n718), .C2(new_n792), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n806), .A2(new_n481), .A3(new_n800), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT48), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(KEYINPUT118), .ZN(new_n830));
  XOR2_X1   g644(.A(new_n828), .B(new_n830), .Z(new_n831));
  OR2_X1    g645(.A1(new_n829), .A2(KEYINPUT118), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n827), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n797), .A2(new_n805), .A3(new_n807), .ZN(new_n834));
  OAI21_X1  g648(.A(KEYINPUT114), .B1(new_n783), .B2(new_n784), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT114), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n815), .A2(new_n836), .A3(new_n782), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n835), .B(new_n837), .C1(new_n556), .C2(new_n817), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n834), .B1(new_n838), .B2(new_n814), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n833), .B1(new_n839), .B2(KEYINPUT51), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n790), .B1(new_n824), .B2(new_n840), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n839), .A2(KEYINPUT51), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n822), .A2(new_n823), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n842), .A2(new_n843), .A3(KEYINPUT119), .A4(new_n833), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n721), .A2(new_n314), .B1(new_n733), .B2(new_n731), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n752), .A2(new_n713), .A3(new_n716), .A4(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT108), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n552), .A2(new_n553), .A3(new_n667), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n849), .B1(new_n306), .B2(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n740), .A2(new_n670), .A3(new_n668), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n700), .A2(KEYINPUT108), .A3(new_n852), .A4(new_n236), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n851), .A2(new_n853), .A3(new_n663), .A4(new_n611), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n750), .A2(new_n704), .A3(new_n737), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n854), .A2(new_n754), .A3(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n646), .B1(new_n700), .B2(new_n638), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n555), .A2(new_n619), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n857), .A2(new_n617), .A3(new_n611), .A4(new_n859), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n612), .A2(new_n660), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n856), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n848), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n738), .A2(new_n677), .A3(new_n705), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT109), .ZN(new_n866));
  AOI211_X1 g680(.A(new_n668), .B(new_n657), .C1(new_n353), .C2(new_n354), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n689), .A2(new_n556), .A3(new_n749), .A4(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n676), .A2(new_n770), .A3(new_n645), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n866), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n355), .A2(new_n656), .A3(new_n667), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n871), .B1(new_n462), .B2(new_n686), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n733), .A2(new_n872), .A3(KEYINPUT109), .A4(new_n611), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT52), .B1(new_n865), .B2(new_n874), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n875), .A2(KEYINPUT110), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n677), .A2(new_n705), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n877), .A2(new_n874), .A3(KEYINPUT52), .A4(new_n738), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n878), .B1(new_n875), .B2(KEYINPUT110), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n846), .B(new_n863), .C1(new_n876), .C2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT52), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n870), .A2(new_n873), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n881), .B1(new_n882), .B2(new_n864), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(new_n878), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n863), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT53), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n880), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(KEYINPUT54), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n856), .A2(new_n861), .A3(KEYINPUT53), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT112), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n889), .B1(new_n890), .B2(new_n848), .ZN(new_n891));
  OR2_X1    g705(.A1(new_n848), .A2(new_n890), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n891), .B(new_n892), .C1(new_n876), .C2(new_n879), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT111), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n894), .B1(new_n885), .B2(new_n846), .ZN(new_n895));
  AOI211_X1 g709(.A(KEYINPUT111), .B(KEYINPUT53), .C1(new_n863), .C2(new_n884), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n893), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n888), .B1(KEYINPUT54), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n789), .B1(new_n845), .B2(new_n898), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n817), .B(KEYINPUT49), .Z(new_n900));
  NOR2_X1   g714(.A1(new_n557), .A2(new_n554), .ZN(new_n901));
  AND4_X1   g715(.A1(new_n724), .A2(new_n690), .A3(new_n691), .A4(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n638), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n900), .A2(new_n902), .A3(new_n700), .A4(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n899), .A2(new_n904), .ZN(G75));
  NAND3_X1  g719(.A1(new_n897), .A2(G210), .A3(G902), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT56), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n517), .B(KEYINPUT120), .Z(new_n909));
  XOR2_X1   g723(.A(new_n522), .B(KEYINPUT55), .Z(new_n910));
  XNOR2_X1  g724(.A(new_n909), .B(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n908), .A2(KEYINPUT121), .A3(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n246), .A2(G952), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT121), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n916), .B1(new_n906), .B2(new_n907), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n906), .A2(new_n916), .A3(new_n907), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n917), .B1(new_n911), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n915), .A2(new_n919), .ZN(G51));
  INV_X1    g734(.A(KEYINPUT54), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n897), .B(new_n921), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n762), .B(KEYINPUT57), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n594), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n761), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n897), .A2(G902), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n913), .B1(new_n924), .B2(new_n926), .ZN(G54));
  NAND4_X1  g741(.A1(new_n897), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n928));
  INV_X1    g742(.A(new_n299), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n928), .A2(new_n929), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n930), .A2(new_n931), .A3(new_n913), .ZN(G60));
  AND2_X1   g746(.A1(new_n631), .A2(new_n633), .ZN(new_n933));
  NAND2_X1  g747(.A1(G478), .A2(G902), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT59), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n914), .B1(new_n922), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n933), .B1(new_n898), .B2(new_n935), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(G63));
  OAI21_X1  g753(.A(KEYINPUT60), .B1(new_n192), .B2(new_n237), .ZN(new_n940));
  OR3_X1    g754(.A1(new_n192), .A2(new_n237), .A3(KEYINPUT60), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n897), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n344), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n897), .A2(new_n655), .A3(new_n940), .A4(new_n941), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n943), .A2(new_n914), .A3(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT61), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n943), .A2(KEYINPUT61), .A3(new_n914), .A4(new_n944), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(G66));
  INV_X1    g763(.A(new_n520), .ZN(new_n950));
  OAI21_X1  g764(.A(G953), .B1(new_n950), .B2(new_n312), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n713), .A2(new_n716), .A3(new_n847), .ZN(new_n952));
  INV_X1    g766(.A(new_n861), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n951), .B1(new_n954), .B2(G953), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n909), .B1(G898), .B2(new_n246), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(G69));
  NAND2_X1  g771(.A1(new_n396), .A2(new_n403), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n294), .B(KEYINPUT122), .Z(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(G900), .B2(G953), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n865), .B1(new_n776), .B2(new_n777), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT124), .Z(new_n963));
  NAND4_X1  g777(.A1(new_n769), .A2(new_n481), .A3(new_n679), .A4(new_n733), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n964), .A2(new_n752), .A3(new_n754), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n963), .A2(new_n787), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n961), .B1(new_n966), .B2(G953), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n857), .B(KEYINPUT123), .Z(new_n968));
  AND3_X1   g782(.A1(new_n750), .A2(new_n481), .A3(new_n679), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n778), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n702), .A2(new_n865), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT62), .Z(new_n972));
  NAND3_X1  g786(.A1(new_n787), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n246), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n960), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n967), .A2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT125), .ZN(new_n977));
  OAI221_X1 g791(.A(G953), .B1(new_n580), .B2(new_n665), .C1(new_n960), .C2(new_n977), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT126), .Z(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n976), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n967), .A2(new_n975), .A3(new_n979), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(G72));
  NAND2_X1  g797(.A1(G472), .A2(G902), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT63), .Z(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT127), .Z(new_n986));
  INV_X1    g800(.A(new_n954), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n986), .B1(new_n973), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n427), .B1(new_n417), .B2(new_n421), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n887), .B(new_n985), .C1(new_n474), .C2(new_n684), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n990), .A2(new_n914), .A3(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n986), .B1(new_n966), .B2(new_n987), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n422), .A2(new_n426), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(G57));
endmodule


