//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 0 0 1 0 0 0 0 1 1 1 0 1 1 1 1 1 0 1 0 0 1 1 0 0 0 0 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1193, new_n1194, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1244, new_n1245,
    new_n1246, new_n1247;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT64), .Z(G355));
  AOI22_X1  g0007(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n208));
  INV_X1    g0008(.A(G116), .ZN(new_n209));
  INV_X1    g0009(.A(G270), .ZN(new_n210));
  OAI21_X1  g0010(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  INV_X1    g0013(.A(G97), .ZN(new_n214));
  INV_X1    g0014(.A(G257), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n212), .B1(new_n203), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n211), .B(new_n216), .C1(G58), .C2(G232), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n217), .B1(G1), .B2(G20), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT1), .Z(new_n219));
  NAND2_X1  g0019(.A1(new_n202), .A2(new_n203), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(G50), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  NOR3_X1   g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G1), .ZN(new_n225));
  NOR3_X1   g0025(.A1(new_n225), .A2(new_n222), .A3(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT0), .Z(new_n228));
  NOR3_X1   g0028(.A1(new_n219), .A2(new_n224), .A3(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT2), .ZN(new_n233));
  INV_X1    g0033(.A(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G264), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(new_n210), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G58), .ZN(new_n241));
  INV_X1    g0041(.A(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n243), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(KEYINPUT18), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n222), .A2(G1), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G13), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT8), .B(G58), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n223), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n256), .A2(new_n250), .ZN(new_n257));
  INV_X1    g0057(.A(new_n253), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(new_n254), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n256), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G58), .A2(G68), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n220), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G20), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT72), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(G20), .A2(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G159), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n264), .A2(KEYINPUT72), .A3(G20), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n267), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT3), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT3), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(KEYINPUT7), .A3(new_n222), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n274), .A2(G33), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n272), .A2(KEYINPUT3), .ZN(new_n279));
  OAI21_X1  g0079(.A(KEYINPUT71), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT71), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n273), .A2(new_n275), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(G20), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n277), .B1(new_n283), .B2(KEYINPUT7), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n271), .B1(new_n284), .B2(G68), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n262), .B1(new_n285), .B2(KEYINPUT16), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT7), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT3), .B(G33), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n287), .B1(new_n288), .B2(G20), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n289), .A2(new_n277), .A3(KEYINPUT73), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT73), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n276), .A2(new_n291), .A3(KEYINPUT7), .A4(new_n222), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n290), .A2(G68), .A3(new_n292), .ZN(new_n293));
  AND3_X1   g0093(.A1(new_n267), .A2(new_n269), .A3(new_n270), .ZN(new_n294));
  AOI21_X1  g0094(.A(KEYINPUT16), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n261), .B1(new_n286), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n225), .B1(G41), .B2(G45), .ZN(new_n298));
  INV_X1    g0098(.A(G274), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G41), .ZN(new_n301));
  OAI211_X1 g0101(.A(G1), .B(G13), .C1(new_n272), .C2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n298), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n303), .A2(new_n231), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n288), .A2(G226), .A3(G1698), .ZN(new_n305));
  INV_X1    g0105(.A(G1698), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n288), .A2(G223), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(G33), .A2(G87), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n305), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n302), .ZN(new_n310));
  AOI211_X1 g0110(.A(new_n300), .B(new_n304), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G179), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n309), .A2(new_n310), .ZN(new_n313));
  INV_X1    g0113(.A(new_n304), .ZN(new_n314));
  INV_X1    g0114(.A(new_n300), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G169), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n249), .B1(new_n297), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n277), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n273), .A2(new_n275), .A3(new_n281), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n281), .B1(new_n273), .B2(new_n275), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n222), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n321), .B1(new_n324), .B2(new_n287), .ZN(new_n325));
  OAI211_X1 g0125(.A(KEYINPUT16), .B(new_n294), .C1(new_n325), .C2(new_n203), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n296), .A2(new_n256), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n260), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n328), .A2(KEYINPUT18), .A3(new_n318), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n320), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT17), .ZN(new_n331));
  INV_X1    g0131(.A(G190), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n313), .A2(new_n332), .A3(new_n314), .A4(new_n315), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(new_n311), .B2(G200), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n326), .A2(new_n256), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n260), .B(new_n334), .C1(new_n335), .C2(new_n295), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT74), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT74), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n327), .A2(new_n338), .A3(new_n260), .A4(new_n334), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n331), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n336), .A2(KEYINPUT17), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n330), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(KEYINPUT75), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n250), .A2(new_n201), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT66), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n346), .A2(new_n251), .A3(new_n262), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n204), .A2(G20), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT65), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n348), .A2(new_n349), .B1(G150), .B2(new_n268), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n349), .B2(new_n348), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n272), .A2(G20), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n351), .B1(new_n352), .B2(new_n258), .ZN(new_n353));
  OAI221_X1 g0153(.A(new_n347), .B1(G50), .B2(new_n251), .C1(new_n353), .C2(new_n262), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT9), .ZN(new_n355));
  OR2_X1    g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n355), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n288), .A2(G223), .A3(G1698), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n288), .A2(new_n306), .ZN(new_n359));
  INV_X1    g0159(.A(G222), .ZN(new_n360));
  OAI221_X1 g0160(.A(new_n358), .B1(new_n242), .B2(new_n288), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n310), .ZN(new_n362));
  INV_X1    g0162(.A(new_n303), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(G226), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n362), .A2(new_n315), .A3(new_n364), .ZN(new_n365));
  XOR2_X1   g0165(.A(KEYINPUT69), .B(G200), .Z(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n365), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(G190), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n356), .A2(new_n357), .A3(new_n367), .A4(new_n369), .ZN(new_n370));
  XNOR2_X1  g0170(.A(new_n370), .B(KEYINPUT10), .ZN(new_n371));
  INV_X1    g0171(.A(G179), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n373), .B(new_n354), .C1(G169), .C2(new_n368), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n268), .ZN(new_n376));
  OAI22_X1  g0176(.A1(new_n253), .A2(new_n376), .B1(new_n222), .B2(new_n242), .ZN(new_n377));
  XNOR2_X1  g0177(.A(KEYINPUT15), .B(G87), .ZN(new_n378));
  INV_X1    g0178(.A(new_n352), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n256), .B1(new_n377), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT67), .ZN(new_n382));
  XNOR2_X1  g0182(.A(new_n381), .B(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n252), .A2(new_n242), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n257), .A2(G77), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  OR2_X1    g0186(.A1(new_n386), .A2(KEYINPUT68), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(KEYINPUT68), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n288), .A2(G1698), .ZN(new_n390));
  INV_X1    g0190(.A(G107), .ZN(new_n391));
  OAI22_X1  g0191(.A1(new_n390), .A2(new_n213), .B1(new_n391), .B2(new_n288), .ZN(new_n392));
  NOR3_X1   g0192(.A1(new_n276), .A2(new_n231), .A3(G1698), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n310), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G244), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n394), .B(new_n315), .C1(new_n395), .C2(new_n303), .ZN(new_n396));
  INV_X1    g0196(.A(G169), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OR2_X1    g0198(.A1(new_n396), .A2(G179), .ZN(new_n399));
  AND3_X1   g0199(.A1(new_n389), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n389), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n396), .A2(new_n366), .ZN(new_n402));
  OR2_X1    g0202(.A1(new_n396), .A2(new_n332), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NOR3_X1   g0205(.A1(new_n375), .A2(new_n400), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n288), .A2(G232), .A3(G1698), .ZN(new_n407));
  NAND2_X1  g0207(.A1(G33), .A2(G97), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n407), .B(new_n408), .C1(new_n359), .C2(new_n234), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n300), .B1(new_n409), .B2(new_n310), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n363), .A2(G238), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT13), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT13), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n410), .A2(new_n414), .A3(new_n411), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(G200), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n352), .A2(G77), .B1(new_n268), .B2(G50), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n222), .B2(G68), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n419), .A2(KEYINPUT11), .A3(new_n256), .ZN(new_n420));
  INV_X1    g0220(.A(new_n257), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n420), .B1(new_n203), .B2(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n251), .A2(G68), .ZN(new_n423));
  XNOR2_X1  g0223(.A(new_n423), .B(KEYINPUT12), .ZN(new_n424));
  AOI21_X1  g0224(.A(KEYINPUT11), .B1(new_n419), .B2(new_n256), .ZN(new_n425));
  NOR3_X1   g0225(.A1(new_n422), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n413), .A2(G190), .A3(new_n415), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n417), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n416), .A2(G169), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT70), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n430), .B1(new_n431), .B2(KEYINPUT14), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(KEYINPUT14), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n431), .A2(KEYINPUT14), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n416), .A2(G169), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n413), .A2(G179), .A3(new_n415), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n432), .A2(new_n433), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n426), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n429), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OR2_X1    g0239(.A1(new_n343), .A2(KEYINPUT75), .ZN(new_n440));
  AND4_X1   g0240(.A1(new_n344), .A2(new_n406), .A3(new_n439), .A4(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(G33), .A2(G116), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n442), .A2(G20), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n288), .A2(new_n222), .A3(G87), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n444), .A2(KEYINPUT83), .A3(KEYINPUT22), .ZN(new_n445));
  NAND2_X1  g0245(.A1(KEYINPUT83), .A2(KEYINPUT22), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n288), .A2(new_n222), .A3(G87), .A4(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n443), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT24), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n222), .A2(G107), .ZN(new_n450));
  XNOR2_X1  g0250(.A(new_n450), .B(KEYINPUT23), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n448), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n449), .B1(new_n448), .B2(new_n451), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n256), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT84), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n448), .A2(new_n451), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT24), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n448), .A2(new_n449), .A3(new_n451), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT84), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n459), .A2(new_n460), .A3(new_n256), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n262), .B(new_n251), .C1(G1), .C2(new_n272), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(new_n391), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n251), .A2(G107), .ZN(new_n466));
  XNOR2_X1  g0266(.A(new_n466), .B(KEYINPUT25), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n462), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n288), .A2(G250), .A3(new_n306), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G294), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n469), .B(new_n470), .C1(new_n390), .C2(new_n215), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n310), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT79), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n473), .A2(new_n301), .A3(KEYINPUT5), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT5), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n475), .B1(KEYINPUT79), .B2(G41), .ZN(new_n476));
  INV_X1    g0276(.A(G45), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n477), .A2(G1), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n474), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  OR2_X1    g0279(.A1(new_n479), .A2(new_n299), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n302), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G264), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n472), .A2(new_n480), .A3(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT85), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n471), .A2(new_n310), .B1(new_n482), .B2(G264), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n487), .A2(KEYINPUT85), .A3(new_n480), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G169), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n484), .A2(new_n372), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n490), .A2(KEYINPUT86), .A3(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT86), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n397), .B1(new_n486), .B2(new_n488), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n494), .B1(new_n495), .B2(new_n491), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n468), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n464), .B1(new_n455), .B2(new_n461), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n489), .A2(G190), .ZN(new_n500));
  INV_X1    g0300(.A(new_n484), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(G200), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n499), .B(new_n467), .C1(new_n500), .C2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n288), .A2(G244), .A3(G1698), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n505), .B(new_n442), .C1(new_n359), .C2(new_n213), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n310), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n478), .A2(G274), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n302), .B(G250), .C1(G1), .C2(new_n477), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G190), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n252), .A2(new_n378), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n352), .A2(G97), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT19), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n222), .B1(new_n408), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(G87), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n516), .A2(new_n214), .A3(new_n391), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n288), .A2(new_n222), .A3(G68), .ZN(new_n519));
  AND2_X1   g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n512), .B1(new_n520), .B2(new_n262), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n463), .A2(new_n516), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n366), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n511), .B(new_n523), .C1(new_n510), .C2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n463), .A2(new_n378), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n509), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n528), .B1(new_n506), .B2(new_n310), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n529), .A2(G179), .A3(new_n508), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n397), .B1(new_n529), .B2(new_n508), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n525), .B1(new_n527), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT80), .ZN(new_n535));
  INV_X1    g0335(.A(new_n480), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n481), .A2(new_n215), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT78), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(new_n359), .B2(new_n395), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT4), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n288), .A2(G250), .A3(G1698), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT4), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n538), .B(new_n542), .C1(new_n359), .C2(new_n395), .ZN(new_n543));
  NAND2_X1  g0343(.A1(G33), .A2(G283), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n540), .A2(new_n541), .A3(new_n543), .A4(new_n544), .ZN(new_n545));
  AOI211_X1 g0345(.A(new_n536), .B(new_n537), .C1(new_n545), .C2(new_n310), .ZN(new_n546));
  INV_X1    g0346(.A(G200), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n535), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n252), .A2(new_n214), .ZN(new_n549));
  OAI22_X1  g0349(.A1(new_n463), .A2(new_n214), .B1(new_n549), .B2(KEYINPUT77), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n290), .A2(G107), .A3(new_n292), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n268), .A2(G77), .ZN(new_n552));
  XOR2_X1   g0352(.A(KEYINPUT76), .B(KEYINPUT6), .Z(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(new_n214), .B2(G107), .ZN(new_n554));
  XNOR2_X1  g0354(.A(G97), .B(G107), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n554), .B1(new_n555), .B2(new_n553), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n551), .B(new_n552), .C1(new_n222), .C2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n550), .B1(new_n557), .B2(new_n256), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n549), .A2(KEYINPUT77), .ZN(new_n559));
  AND2_X1   g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n546), .A2(G190), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n545), .A2(new_n310), .ZN(new_n562));
  INV_X1    g0362(.A(new_n537), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n562), .A2(new_n480), .A3(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n564), .A2(KEYINPUT80), .A3(G200), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n548), .A2(new_n560), .A3(new_n561), .A4(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n546), .A2(new_n372), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n564), .A2(new_n397), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n558), .A2(new_n559), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n534), .A2(new_n566), .A3(new_n570), .ZN(new_n571));
  OR2_X1    g0371(.A1(new_n463), .A2(new_n209), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n544), .B(new_n222), .C1(G33), .C2(new_n214), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n573), .B(new_n256), .C1(new_n222), .C2(G116), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT20), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n574), .A2(new_n575), .ZN(new_n577));
  OAI221_X1 g0377(.A(new_n572), .B1(G116), .B2(new_n251), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n480), .B1(new_n210), .B2(new_n481), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(KEYINPUT81), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT81), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n480), .B(new_n582), .C1(new_n210), .C2(new_n481), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n288), .A2(G257), .A3(new_n306), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n288), .A2(G264), .A3(G1698), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n276), .A2(G303), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT82), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT82), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n585), .A2(new_n586), .A3(new_n590), .A4(new_n587), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n310), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n584), .A2(new_n592), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n579), .A2(new_n593), .A3(new_n372), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n593), .A2(G200), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n596), .B(new_n579), .C1(new_n332), .C2(new_n593), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n397), .B1(new_n584), .B2(new_n592), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT21), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n598), .A2(new_n599), .A3(new_n578), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n599), .B1(new_n598), .B2(new_n578), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n595), .B(new_n597), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  NOR3_X1   g0402(.A1(new_n504), .A2(new_n571), .A3(new_n602), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n441), .A2(new_n603), .ZN(G372));
  INV_X1    g0404(.A(new_n374), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n400), .A2(new_n428), .B1(new_n437), .B2(new_n438), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n340), .A2(new_n341), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n330), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n605), .B1(new_n608), .B2(new_n371), .ZN(new_n609));
  INV_X1    g0409(.A(new_n441), .ZN(new_n610));
  OAI21_X1  g0410(.A(KEYINPUT87), .B1(new_n530), .B2(new_n531), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT87), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n529), .A2(G179), .A3(new_n508), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n612), .B(new_n613), .C1(new_n510), .C2(new_n397), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n527), .B1(new_n611), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n525), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n570), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT26), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n615), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(KEYINPUT26), .B1(new_n533), .B2(new_n570), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n495), .A2(new_n491), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n621), .B1(new_n499), .B2(new_n467), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n595), .B1(new_n600), .B2(new_n601), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n503), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n566), .A2(new_n570), .A3(new_n525), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n619), .B(new_n620), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n609), .B1(new_n610), .B2(new_n627), .ZN(new_n628));
  XOR2_X1   g0428(.A(new_n628), .B(KEYINPUT88), .Z(G369));
  INV_X1    g0429(.A(G330), .ZN(new_n630));
  INV_X1    g0430(.A(new_n623), .ZN(new_n631));
  INV_X1    g0431(.A(G13), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n632), .A2(G20), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n225), .ZN(new_n634));
  OR2_X1    g0434(.A1(new_n634), .A2(KEYINPUT27), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(KEYINPUT27), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(G213), .A3(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(G343), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n631), .B(new_n597), .C1(new_n579), .C2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n623), .A2(new_n578), .A3(new_n639), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n630), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n640), .B1(new_n499), .B2(new_n467), .ZN(new_n644));
  OAI22_X1  g0444(.A1(new_n504), .A2(new_n644), .B1(new_n498), .B2(new_n640), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n622), .A2(new_n640), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n631), .A2(new_n639), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n648), .A2(new_n503), .A3(new_n498), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n646), .A2(new_n647), .A3(new_n649), .ZN(G399));
  INV_X1    g0450(.A(new_n226), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n651), .A2(G41), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n517), .A2(G116), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(G1), .A3(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n655), .B1(new_n221), .B2(new_n653), .ZN(new_n656));
  XNOR2_X1  g0456(.A(new_n656), .B(KEYINPUT28), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n627), .A2(new_n639), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT29), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n566), .A2(new_n570), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT92), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n566), .A2(KEYINPUT92), .A3(new_n570), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n615), .A2(new_n616), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n631), .A2(new_n498), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n665), .A2(new_n503), .A3(new_n666), .A4(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n615), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n669), .B1(new_n617), .B2(new_n618), .ZN(new_n670));
  NOR3_X1   g0470(.A1(new_n533), .A2(new_n570), .A3(KEYINPUT26), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n639), .B1(new_n668), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n660), .B1(new_n659), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n603), .A2(new_n640), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n530), .A2(new_n562), .A3(new_n480), .A4(new_n563), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n584), .A2(new_n487), .A3(new_n592), .ZN(new_n677));
  OAI21_X1  g0477(.A(KEYINPUT89), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n584), .A2(new_n592), .A3(new_n487), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT89), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n679), .A2(new_n546), .A3(new_n680), .A4(new_n530), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT30), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n678), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n679), .A2(new_n546), .A3(KEYINPUT30), .A4(new_n530), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n510), .A2(G179), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n564), .A2(new_n685), .A3(new_n484), .A4(new_n593), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n683), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT91), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT91), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n683), .A2(new_n684), .A3(new_n689), .A4(new_n686), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n688), .A2(new_n639), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT31), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n683), .A2(new_n686), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT90), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n683), .A2(KEYINPUT90), .A3(new_n686), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(new_n684), .A3(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n698), .A2(KEYINPUT31), .A3(new_n639), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n675), .A2(new_n693), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n674), .B1(G330), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n657), .B1(new_n701), .B2(G1), .ZN(G364));
  AOI21_X1  g0502(.A(new_n223), .B1(G20), .B2(new_n397), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n222), .A2(G179), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n366), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G190), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(new_n391), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n705), .A2(new_n332), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(G190), .A2(G200), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n704), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G159), .ZN(new_n714));
  OAI22_X1  g0514(.A1(new_n710), .A2(new_n516), .B1(KEYINPUT32), .B2(new_n714), .ZN(new_n715));
  AOI211_X1 g0515(.A(new_n708), .B(new_n715), .C1(KEYINPUT32), .C2(new_n714), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n222), .A2(new_n372), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G200), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(G190), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n288), .B1(new_n720), .B2(new_n203), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n718), .A2(new_n332), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n332), .A2(G179), .A3(G200), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n222), .ZN(new_n725));
  OAI22_X1  g0525(.A1(new_n723), .A2(new_n201), .B1(new_n214), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n717), .A2(G190), .A3(new_n547), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT94), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n727), .A2(new_n728), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  AOI211_X1 g0533(.A(new_n721), .B(new_n726), .C1(new_n733), .C2(G58), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n717), .A2(new_n711), .ZN(new_n735));
  OAI211_X1 g0535(.A(new_n716), .B(new_n734), .C1(new_n242), .C2(new_n735), .ZN(new_n736));
  XNOR2_X1  g0536(.A(new_n736), .B(KEYINPUT95), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n733), .A2(G322), .ZN(new_n738));
  INV_X1    g0538(.A(G326), .ZN(new_n739));
  INV_X1    g0539(.A(G294), .ZN(new_n740));
  OAI22_X1  g0540(.A1(new_n723), .A2(new_n739), .B1(new_n740), .B2(new_n725), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n288), .B1(new_n713), .B2(G329), .ZN(new_n742));
  XOR2_X1   g0542(.A(KEYINPUT33), .B(G317), .Z(new_n743));
  OAI21_X1  g0543(.A(new_n742), .B1(new_n720), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  AOI22_X1  g0545(.A1(G283), .A2(new_n706), .B1(new_n709), .B2(G303), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n738), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n735), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n747), .B1(G311), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n703), .B1(new_n737), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G13), .A2(G33), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n703), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n322), .A2(new_n323), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n651), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n220), .A2(new_n477), .A3(G50), .ZN(new_n758));
  OAI211_X1 g0558(.A(new_n757), .B(new_n758), .C1(new_n243), .C2(new_n477), .ZN(new_n759));
  NAND3_X1  g0559(.A1(G355), .A2(new_n226), .A3(new_n288), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n759), .B(new_n760), .C1(G116), .C2(new_n226), .ZN(new_n761));
  XOR2_X1   g0561(.A(new_n761), .B(KEYINPUT93), .Z(new_n762));
  NAND2_X1  g0562(.A1(new_n641), .A2(new_n642), .ZN(new_n763));
  XOR2_X1   g0563(.A(new_n753), .B(KEYINPUT96), .Z(new_n764));
  OAI221_X1 g0564(.A(new_n750), .B1(new_n755), .B2(new_n762), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n225), .B1(new_n633), .B2(G45), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n652), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n768), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n763), .A2(G330), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n770), .B1(new_n771), .B2(new_n643), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT97), .Z(G396));
  INV_X1    g0574(.A(G283), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n720), .A2(new_n775), .B1(new_n735), .B2(new_n209), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n776), .A2(KEYINPUT98), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(KEYINPUT98), .ZN(new_n778));
  INV_X1    g0578(.A(G303), .ZN(new_n779));
  OAI211_X1 g0579(.A(new_n777), .B(new_n778), .C1(new_n779), .C2(new_n723), .ZN(new_n780));
  OR2_X1    g0580(.A1(new_n780), .A2(KEYINPUT99), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(KEYINPUT99), .ZN(new_n782));
  INV_X1    g0582(.A(G311), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n276), .B1(new_n783), .B2(new_n712), .C1(new_n710), .C2(new_n391), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n784), .B1(G87), .B2(new_n706), .ZN(new_n785));
  INV_X1    g0585(.A(new_n725), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n733), .A2(G294), .B1(G97), .B2(new_n786), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n781), .A2(new_n782), .A3(new_n785), .A4(new_n787), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n722), .A2(G137), .B1(new_n748), .B2(G159), .ZN(new_n789));
  INV_X1    g0589(.A(G150), .ZN(new_n790));
  INV_X1    g0590(.A(G143), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n789), .B1(new_n790), .B2(new_n720), .C1(new_n732), .C2(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT100), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n793), .B(KEYINPUT34), .Z(new_n794));
  AOI22_X1  g0594(.A1(G50), .A2(new_n709), .B1(new_n706), .B2(G68), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n756), .B1(new_n202), .B2(new_n725), .C1(new_n795), .C2(KEYINPUT101), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n796), .B1(KEYINPUT101), .B2(new_n795), .ZN(new_n797));
  INV_X1    g0597(.A(G132), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n797), .B1(new_n798), .B2(new_n712), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n788), .B1(new_n794), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n703), .A2(new_n751), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n800), .A2(new_n703), .B1(new_n242), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n389), .A2(new_n639), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n389), .A2(new_n398), .A3(new_n399), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(KEYINPUT102), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT102), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n387), .A2(new_n388), .B1(new_n397), .B2(new_n396), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n806), .B1(new_n807), .B2(new_n399), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n404), .B(new_n803), .C1(new_n805), .C2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n400), .A2(new_n639), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n768), .B(new_n802), .C1(new_n811), .C2(new_n752), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n400), .A2(new_n806), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n804), .A2(KEYINPUT102), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n405), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n626), .A2(new_n640), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n658), .B2(new_n811), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n700), .A2(G330), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n817), .B(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n812), .B1(new_n819), .B2(new_n768), .ZN(G384));
  NAND2_X1  g0620(.A1(new_n437), .A2(new_n438), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n821), .B(new_n428), .C1(new_n426), .C2(new_n640), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n438), .B(new_n639), .C1(new_n437), .C2(new_n429), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n811), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT108), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n826), .A2(KEYINPUT31), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n688), .A2(new_n639), .A3(new_n690), .A4(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n826), .B1(KEYINPUT107), .B2(KEYINPUT31), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n603), .A2(new_n640), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n830), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n688), .A2(new_n639), .A3(new_n690), .A4(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n825), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n337), .A2(new_n339), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT37), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n328), .A2(new_n318), .ZN(new_n837));
  INV_X1    g0637(.A(new_n637), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n328), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n835), .A2(new_n836), .A3(new_n837), .A4(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n286), .B1(KEYINPUT16), .B2(new_n285), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n260), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n319), .A2(new_n637), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n337), .A2(new_n339), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n840), .B1(new_n836), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n637), .B1(new_n841), .B2(new_n260), .ZN(new_n846));
  AND3_X1   g0646(.A1(new_n342), .A2(KEYINPUT104), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(KEYINPUT104), .B1(new_n342), .B2(new_n846), .ZN(new_n848));
  OAI211_X1 g0648(.A(KEYINPUT38), .B(new_n845), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  AND3_X1   g0649(.A1(new_n837), .A2(new_n839), .A3(new_n336), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n840), .B1(new_n850), .B2(new_n836), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n343), .B2(new_n839), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT38), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n849), .A2(new_n854), .ZN(new_n855));
  AND3_X1   g0655(.A1(new_n834), .A2(KEYINPUT40), .A3(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT40), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT105), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n342), .A2(new_n846), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT104), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n342), .A2(KEYINPUT104), .A3(new_n846), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(KEYINPUT38), .B1(new_n863), .B2(new_n845), .ZN(new_n864));
  INV_X1    g0664(.A(new_n849), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n858), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n845), .B1(new_n847), .B2(new_n848), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n853), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n868), .A2(KEYINPUT105), .A3(new_n849), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n866), .A2(new_n869), .A3(new_n834), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n856), .B1(new_n857), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n829), .A2(new_n830), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n675), .A2(new_n872), .A3(new_n833), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n441), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n871), .B(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(G330), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n674), .A2(new_n441), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n609), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n876), .B(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n821), .A2(new_n639), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT39), .B1(new_n864), .B2(new_n865), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT106), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT39), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n849), .A2(new_n854), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n882), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n884), .B1(new_n868), .B2(new_n849), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n849), .A2(new_n854), .A3(new_n884), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT106), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n881), .B1(new_n886), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n813), .A2(new_n640), .A3(new_n814), .ZN(new_n891));
  OR2_X1    g0691(.A1(new_n891), .A2(KEYINPUT103), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(KEYINPUT103), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n816), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n894), .A2(new_n824), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n895), .A2(new_n866), .A3(new_n869), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n330), .A2(new_n838), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n890), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n879), .B(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n225), .B2(new_n633), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT35), .ZN(new_n903));
  AOI211_X1 g0703(.A(new_n222), .B(new_n223), .C1(new_n556), .C2(new_n903), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n904), .B(G116), .C1(new_n903), .C2(new_n556), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT36), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n263), .A2(G77), .ZN(new_n907));
  OAI22_X1  g0707(.A1(new_n221), .A2(new_n907), .B1(G50), .B2(new_n203), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n908), .A2(G1), .A3(new_n632), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n902), .A2(new_n906), .A3(new_n909), .ZN(G367));
  NOR2_X1   g0710(.A1(new_n523), .A2(new_n640), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n669), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n666), .B2(new_n911), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(KEYINPUT109), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(KEYINPUT43), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n569), .A2(new_n639), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n665), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n917), .A2(new_n649), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n918), .B(KEYINPUT42), .Z(new_n919));
  OR2_X1    g0719(.A1(new_n917), .A2(new_n498), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n639), .B1(new_n920), .B2(new_n570), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n915), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n570), .A2(new_n640), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(new_n665), .B2(new_n916), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n646), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n922), .B(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n914), .A2(KEYINPUT43), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n926), .B(new_n927), .ZN(new_n928));
  XOR2_X1   g0728(.A(KEYINPUT110), .B(KEYINPUT41), .Z(new_n929));
  XOR2_X1   g0729(.A(new_n652), .B(new_n929), .Z(new_n930));
  NAND2_X1  g0730(.A1(new_n649), .A2(new_n647), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n931), .A2(new_n924), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT111), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n933), .A2(KEYINPUT45), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(KEYINPUT45), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n931), .A2(new_n924), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n936), .B(KEYINPUT44), .Z(new_n937));
  NAND3_X1  g0737(.A1(new_n934), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(new_n646), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n649), .B1(new_n645), .B2(new_n648), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(new_n643), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n939), .A2(new_n701), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n930), .B1(new_n942), .B2(new_n701), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n928), .B1(new_n943), .B2(new_n767), .ZN(new_n944));
  INV_X1    g0744(.A(new_n757), .ZN(new_n945));
  OAI221_X1 g0745(.A(new_n754), .B1(new_n226), .B2(new_n378), .C1(new_n238), .C2(new_n945), .ZN(new_n946));
  OAI22_X1  g0746(.A1(new_n202), .A2(new_n710), .B1(new_n707), .B2(new_n242), .ZN(new_n947));
  OAI22_X1  g0747(.A1(new_n723), .A2(new_n791), .B1(new_n203), .B2(new_n725), .ZN(new_n948));
  INV_X1    g0748(.A(G137), .ZN(new_n949));
  OAI221_X1 g0749(.A(new_n288), .B1(new_n712), .B2(new_n949), .C1(new_n201), .C2(new_n735), .ZN(new_n950));
  NOR3_X1   g0750(.A1(new_n947), .A2(new_n948), .A3(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(G159), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n951), .B1(new_n790), .B2(new_n732), .C1(new_n952), .C2(new_n720), .ZN(new_n953));
  XOR2_X1   g0753(.A(KEYINPUT113), .B(G317), .Z(new_n954));
  OAI22_X1  g0754(.A1(new_n720), .A2(new_n740), .B1(new_n954), .B2(new_n712), .ZN(new_n955));
  INV_X1    g0755(.A(new_n756), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n391), .B2(new_n725), .ZN(new_n957));
  AOI211_X1 g0757(.A(new_n955), .B(new_n957), .C1(G97), .C2(new_n706), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n732), .A2(new_n779), .B1(new_n783), .B2(new_n723), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT112), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n959), .A2(new_n960), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n709), .A2(G116), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT46), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n958), .A2(new_n961), .A3(new_n962), .A4(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n735), .A2(new_n775), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n953), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT47), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n770), .B1(new_n968), .B2(new_n703), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n946), .B(new_n969), .C1(new_n914), .C2(new_n764), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n944), .A2(new_n970), .ZN(G387));
  OR2_X1    g0771(.A1(new_n701), .A2(new_n941), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n701), .A2(new_n941), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n972), .A2(new_n652), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n941), .A2(new_n767), .ZN(new_n975));
  INV_X1    g0775(.A(new_n654), .ZN(new_n976));
  AOI211_X1 g0776(.A(G45), .B(new_n976), .C1(G68), .C2(G77), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n978), .A2(KEYINPUT114), .ZN(new_n979));
  OR3_X1    g0779(.A1(new_n253), .A2(KEYINPUT50), .A3(G50), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n978), .A2(KEYINPUT114), .ZN(new_n981));
  OAI21_X1  g0781(.A(KEYINPUT50), .B1(new_n253), .B2(G50), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n979), .A2(new_n980), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  AND2_X1   g0783(.A1(new_n983), .A2(new_n757), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n235), .A2(new_n477), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n984), .A2(new_n985), .B1(new_n391), .B2(new_n651), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n976), .A2(new_n226), .A3(new_n288), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n755), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AOI22_X1  g0788(.A1(G68), .A2(new_n748), .B1(new_n713), .B2(G150), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n253), .B2(new_n720), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(G77), .B2(new_n709), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n725), .A2(new_n378), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(new_n733), .B2(G50), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n706), .A2(G97), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n956), .B1(G159), .B2(new_n722), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n991), .A2(new_n993), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n719), .A2(G311), .B1(new_n722), .B2(G322), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n997), .B1(new_n779), .B2(new_n735), .C1(new_n732), .C2(new_n954), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT48), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n999), .B1(new_n775), .B2(new_n725), .C1(new_n740), .C2(new_n710), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT49), .Z(new_n1001));
  OAI221_X1 g0801(.A(new_n956), .B1(new_n739), .B2(new_n712), .C1(new_n707), .C2(new_n209), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT115), .Z(new_n1003));
  OAI21_X1  g0803(.A(new_n996), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n988), .B1(new_n1004), .B2(new_n703), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n1005), .B(new_n768), .C1(new_n645), .C2(new_n764), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n974), .A2(new_n975), .A3(new_n1006), .ZN(G393));
  INV_X1    g0807(.A(new_n973), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n939), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1009), .A2(new_n652), .A3(new_n942), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n754), .B1(new_n214), .B2(new_n226), .C1(new_n945), .C2(new_n247), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n924), .A2(new_n753), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT116), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n924), .A2(KEYINPUT116), .A3(new_n753), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n203), .A2(new_n710), .B1(new_n707), .B2(new_n516), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n720), .A2(new_n201), .B1(new_n712), .B2(new_n791), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n725), .A2(new_n242), .ZN(new_n1018));
  OR3_X1    g0818(.A1(new_n1017), .A2(new_n956), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT51), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n732), .A2(new_n952), .B1(new_n790), .B2(new_n723), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n1016), .B(new_n1019), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1022), .B1(new_n1020), .B2(new_n1021), .C1(new_n253), .C2(new_n735), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n733), .A2(G311), .B1(G317), .B2(new_n722), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT52), .Z(new_n1025));
  AOI22_X1  g0825(.A1(new_n786), .A2(G116), .B1(new_n748), .B2(G294), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n779), .B2(new_n720), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT117), .Z(new_n1028));
  AOI21_X1  g0828(.A(new_n288), .B1(new_n713), .B2(G322), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n708), .B1(G283), .B2(new_n709), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1025), .A2(new_n1028), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1023), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n770), .B1(new_n1032), .B2(new_n703), .ZN(new_n1033));
  AND4_X1   g0833(.A1(new_n1011), .A2(new_n1014), .A3(new_n1015), .A4(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n939), .B2(new_n767), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1010), .A2(new_n1035), .ZN(G390));
  NAND3_X1  g0836(.A1(new_n441), .A2(G330), .A3(new_n873), .ZN(new_n1037));
  AND3_X1   g0837(.A1(new_n877), .A2(new_n609), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n811), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1039), .A2(new_n630), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n873), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n824), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1041), .A2(KEYINPUT119), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT118), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n891), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1044), .B(new_n1045), .C1(new_n673), .C2(new_n815), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n668), .A2(new_n672), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1047), .A2(new_n640), .A3(new_n815), .ZN(new_n1048));
  AOI21_X1  g0848(.A(KEYINPUT118), .B1(new_n1048), .B2(new_n891), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1043), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n824), .B1(new_n1040), .B2(new_n873), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n700), .A2(G330), .A3(new_n811), .A4(new_n824), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1051), .B1(KEYINPUT119), .B2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1050), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n894), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1042), .B1(new_n818), .B2(new_n1039), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1040), .A2(new_n873), .A3(new_n824), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1055), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1038), .B1(new_n1054), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1057), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n813), .A2(new_n814), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n404), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n639), .B(new_n1062), .C1(new_n668), .C2(new_n672), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1044), .B1(new_n1063), .B2(new_n1045), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1048), .A2(KEYINPUT118), .A3(new_n891), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1064), .A2(new_n824), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n880), .B1(new_n849), .B2(new_n854), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n881), .B1(new_n1055), .B2(new_n1042), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n886), .A2(new_n889), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1060), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1052), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1068), .A2(new_n1070), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1059), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1075), .A2(new_n653), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n877), .A2(new_n609), .A3(new_n1037), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n1052), .A2(KEYINPUT119), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1079), .B(new_n1043), .C1(new_n1080), .C2(new_n1051), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1058), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1078), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1076), .B1(new_n1077), .B2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n886), .A2(new_n889), .A3(new_n751), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n203), .A2(new_n707), .B1(new_n710), .B2(new_n516), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n276), .B1(new_n712), .B2(new_n740), .C1(new_n720), .C2(new_n391), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n723), .A2(new_n775), .ZN(new_n1088));
  NOR4_X1   g0888(.A1(new_n1086), .A2(new_n1087), .A3(new_n1018), .A4(new_n1088), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1089), .B1(new_n214), .B2(new_n735), .C1(new_n209), .C2(new_n732), .ZN(new_n1090));
  INV_X1    g0890(.A(G125), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n712), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(G128), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n723), .A2(new_n1093), .B1(new_n952), .B2(new_n725), .ZN(new_n1094));
  XOR2_X1   g0894(.A(KEYINPUT54), .B(G143), .Z(new_n1095));
  NAND2_X1  g0895(.A1(new_n748), .A2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n288), .B(new_n1096), .C1(new_n720), .C2(new_n949), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n1094), .B(new_n1097), .C1(G50), .C2(new_n706), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n709), .A2(G150), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n1099), .B(KEYINPUT53), .Z(new_n1100));
  OAI211_X1 g0900(.A(new_n1098), .B(new_n1100), .C1(new_n798), .C2(new_n732), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1090), .B1(new_n1092), .B2(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n1102), .A2(new_n703), .B1(new_n253), .B2(new_n801), .ZN(new_n1103));
  AND3_X1   g0903(.A1(new_n1085), .A2(new_n768), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n1077), .B2(new_n767), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1084), .A2(new_n1105), .ZN(G378));
  INV_X1    g0906(.A(KEYINPUT122), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n870), .A2(new_n857), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n856), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1108), .A2(G330), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n883), .B1(new_n882), .B2(new_n885), .ZN(new_n1111));
  NOR3_X1   g0911(.A1(new_n887), .A2(new_n888), .A3(KEYINPUT106), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n880), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n896), .A2(new_n898), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1110), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  OAI211_X1 g0915(.A(G330), .B(new_n871), .C1(new_n890), .C2(new_n899), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n354), .A2(new_n838), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n375), .B(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT55), .ZN(new_n1120));
  XOR2_X1   g0920(.A(new_n1120), .B(KEYINPUT56), .Z(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1117), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1115), .A2(new_n1116), .A3(new_n1121), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1068), .A2(new_n1070), .A3(new_n1073), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1083), .B1(new_n1125), .B2(new_n1071), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1123), .A2(new_n1124), .B1(new_n1038), .B2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1107), .B1(new_n1127), .B2(KEYINPUT57), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n653), .B1(new_n1127), .B2(KEYINPUT57), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1124), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1121), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n1130), .A2(new_n1131), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT57), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1132), .A2(KEYINPUT122), .A3(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1128), .A2(new_n1129), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n766), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n725), .A2(new_n790), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n723), .A2(new_n1091), .B1(new_n735), .B2(new_n949), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n1137), .B(new_n1138), .C1(new_n709), .C2(new_n1095), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n1139), .B1(new_n1093), .B2(new_n732), .C1(new_n798), .C2(new_n720), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n1141));
  OR2_X1    g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1143));
  AOI21_X1  g0943(.A(G33), .B1(new_n713), .B2(G124), .ZN(new_n1144));
  AOI21_X1  g0944(.A(G41), .B1(new_n706), .B2(G159), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n706), .A2(G58), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n710), .B2(new_n242), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n732), .A2(new_n391), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n301), .B1(new_n712), .B2(new_n775), .C1(new_n378), .C2(new_n735), .ZN(new_n1150));
  NOR4_X1   g0950(.A1(new_n1148), .A2(new_n1149), .A3(new_n756), .A4(new_n1150), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(G68), .A2(new_n786), .B1(new_n722), .B2(G116), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT120), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1151), .B(new_n1153), .C1(new_n214), .C2(new_n720), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT58), .ZN(new_n1155));
  AOI21_X1  g0955(.A(G41), .B1(new_n756), .B2(G33), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1146), .B(new_n1155), .C1(G50), .C2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n770), .B1(new_n1157), .B2(new_n703), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n1122), .B2(new_n752), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n201), .B2(new_n801), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1136), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1135), .A2(new_n1161), .ZN(G375));
  NOR2_X1   g0962(.A1(new_n1054), .A2(new_n1058), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n1078), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n930), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1164), .A2(new_n1165), .A3(new_n1059), .ZN(new_n1166));
  XOR2_X1   g0966(.A(new_n1166), .B(KEYINPUT123), .Z(new_n1167));
  NAND2_X1  g0967(.A1(new_n1042), .A2(new_n751), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n242), .A2(new_n707), .B1(new_n710), .B2(new_n214), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n276), .B1(new_n391), .B2(new_n735), .C1(new_n720), .C2(new_n209), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n723), .A2(new_n740), .ZN(new_n1171));
  NOR4_X1   g0971(.A1(new_n1169), .A2(new_n1170), .A3(new_n992), .A4(new_n1171), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n1172), .B1(new_n775), .B2(new_n732), .C1(new_n779), .C2(new_n712), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(G150), .A2(new_n748), .B1(new_n713), .B2(G128), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1147), .B(new_n1174), .C1(new_n710), .C2(new_n952), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n719), .B2(new_n1095), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n756), .B1(new_n201), .B2(new_n725), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n733), .B2(G137), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1176), .B(new_n1178), .C1(new_n798), .C2(new_n723), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1173), .A2(new_n1179), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n1180), .A2(new_n703), .B1(new_n203), .B2(new_n801), .ZN(new_n1181));
  AND3_X1   g0981(.A1(new_n1168), .A2(new_n768), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1163), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1182), .B1(new_n1183), .B2(new_n767), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1167), .A2(new_n1184), .ZN(G381));
  INV_X1    g0985(.A(KEYINPUT124), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(G378), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1084), .A2(new_n1105), .A3(KEYINPUT124), .ZN(new_n1188));
  AOI21_X1  g0988(.A(G375), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(G387), .A2(G390), .A3(G384), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(G381), .A2(G396), .A3(G393), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(G407));
  INV_X1    g0992(.A(G213), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n1189), .B2(new_n638), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(G407), .ZN(G409));
  NOR2_X1   g0995(.A1(new_n1193), .A2(G343), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1135), .A2(G378), .A3(new_n1161), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT125), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1135), .A2(KEYINPUT125), .A3(G378), .A4(new_n1161), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1127), .A2(new_n1165), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1187), .A2(new_n1188), .B1(new_n1161), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1196), .B1(new_n1201), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT126), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT60), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n653), .B1(new_n1164), .B2(new_n1207), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1208), .B(new_n1059), .C1(new_n1207), .C2(new_n1164), .ZN(new_n1209));
  AND3_X1   g1009(.A1(new_n1209), .A2(G384), .A3(new_n1184), .ZN(new_n1210));
  AOI21_X1  g1010(.A(G384), .B1(new_n1209), .B2(new_n1184), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1206), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n1210), .A2(new_n1211), .A3(new_n1206), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1196), .A2(G2897), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1212), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n1214), .B2(new_n1212), .ZN(new_n1216));
  OAI21_X1  g1016(.A(KEYINPUT63), .B1(new_n1205), .B2(new_n1216), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1205), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1217), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT61), .ZN(new_n1222));
  INV_X1    g1022(.A(G390), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(G387), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  XOR2_X1   g1025(.A(G393), .B(G396), .Z(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(G387), .A2(new_n1223), .ZN(new_n1228));
  OR3_X1    g1028(.A1(new_n1225), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1227), .B1(new_n1225), .B2(new_n1228), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1203), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(new_n1232), .A2(new_n1218), .A3(new_n1196), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1231), .B1(new_n1233), .B2(KEYINPUT63), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1221), .A2(new_n1222), .A3(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1222), .B1(new_n1205), .B2(new_n1216), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT62), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n1205), .B2(new_n1219), .ZN(new_n1238));
  NOR4_X1   g1038(.A1(new_n1232), .A2(KEYINPUT62), .A3(new_n1218), .A4(new_n1196), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(new_n1236), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT127), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1231), .B(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1235), .B1(new_n1240), .B2(new_n1242), .ZN(G405));
  NAND2_X1  g1043(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(G375), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1201), .A2(new_n1245), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1246), .B(new_n1219), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(new_n1231), .ZN(G402));
endmodule


