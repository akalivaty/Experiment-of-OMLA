//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 0 1 0 0 1 1 0 0 0 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 0 1 1 1 1 0 1 0 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1268, new_n1269, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(new_n202), .A2(G50), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G13), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(new_n208), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(KEYINPUT64), .B(G77), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n220), .B1(G244), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(KEYINPUT65), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n223), .A2(KEYINPUT65), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n213), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n210), .B(new_n216), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G226), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  NAND2_X1  g0047(.A1(G33), .A2(G41), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n248), .A2(G1), .A3(G13), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT3), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G33), .ZN(new_n254));
  NAND4_X1  g0054(.A1(new_n252), .A2(new_n254), .A3(G264), .A4(G1698), .ZN(new_n255));
  INV_X1    g0055(.A(G303), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT3), .B(G33), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  AND3_X1   g0059(.A1(new_n257), .A2(G257), .A3(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n250), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G45), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(G1), .ZN(new_n263));
  AND2_X1   g0063(.A1(KEYINPUT5), .A2(G41), .ZN(new_n264));
  NOR2_X1   g0064(.A1(KEYINPUT5), .A2(G41), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AND2_X1   g0066(.A1(G33), .A2(G41), .ZN(new_n267));
  OAI21_X1  g0067(.A(G274), .B1(new_n267), .B2(new_n207), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT5), .B(G41), .ZN(new_n270));
  INV_X1    g0070(.A(new_n207), .ZN(new_n271));
  AOI22_X1  g0071(.A1(new_n270), .A2(new_n263), .B1(new_n271), .B2(new_n248), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n269), .B1(G270), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n261), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT82), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G13), .ZN(new_n277));
  NOR3_X1   g0077(.A1(new_n277), .A2(new_n208), .A3(G1), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n207), .ZN(new_n280));
  OR3_X1    g0080(.A1(new_n278), .A2(new_n280), .A3(KEYINPUT71), .ZN(new_n281));
  OAI21_X1  g0081(.A(KEYINPUT71), .B1(new_n278), .B2(new_n280), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n211), .A2(G33), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n281), .A2(G116), .A3(new_n282), .A4(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT80), .B(G116), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G20), .ZN(new_n286));
  NOR3_X1   g0086(.A1(new_n286), .A2(G1), .A3(new_n277), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n280), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n289), .B1(G20), .B2(new_n285), .ZN(new_n290));
  NAND2_X1  g0090(.A1(G33), .A2(G283), .ZN(new_n291));
  INV_X1    g0091(.A(G97), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n291), .B(new_n208), .C1(G33), .C2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(KEYINPUT20), .B1(new_n290), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n286), .A2(new_n280), .A3(new_n293), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT20), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n284), .B(new_n288), .C1(new_n294), .C2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n261), .A2(new_n273), .A3(KEYINPUT82), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n276), .A2(new_n298), .A3(G169), .A4(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT21), .ZN(new_n301));
  OAI21_X1  g0101(.A(KEYINPUT83), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  AND3_X1   g0102(.A1(new_n261), .A2(new_n273), .A3(KEYINPUT82), .ZN(new_n303));
  AOI21_X1  g0103(.A(KEYINPUT82), .B1(new_n261), .B2(new_n273), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G169), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n290), .A2(KEYINPUT20), .A3(new_n293), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n295), .A2(new_n296), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n287), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n306), .B1(new_n309), .B2(new_n284), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT83), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n305), .A2(new_n310), .A3(new_n311), .A4(KEYINPUT21), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n302), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(KEYINPUT21), .B1(new_n305), .B2(new_n310), .ZN(new_n314));
  INV_X1    g0114(.A(G179), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n274), .A2(new_n315), .ZN(new_n316));
  AND2_X1   g0116(.A1(new_n316), .A2(new_n298), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  AND2_X1   g0118(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(G190), .B1(new_n303), .B2(new_n304), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n276), .A2(G200), .A3(new_n299), .ZN(new_n321));
  INV_X1    g0121(.A(new_n298), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT84), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n323), .B(new_n324), .ZN(new_n325));
  XNOR2_X1  g0125(.A(G97), .B(G107), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT6), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NOR3_X1   g0128(.A1(new_n327), .A2(new_n292), .A3(G107), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NOR2_X1   g0131(.A1(G20), .A2(G33), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n331), .A2(G20), .B1(G77), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT7), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n334), .B1(new_n257), .B2(G20), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n252), .A2(new_n254), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g0138(.A(KEYINPUT69), .B(G107), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n289), .B1(new_n333), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n278), .A2(new_n292), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n278), .A2(new_n280), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n283), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n342), .B1(new_n344), .B2(new_n292), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n266), .A2(G257), .A3(new_n249), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n270), .A2(new_n249), .A3(G274), .A4(new_n263), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n252), .A2(new_n254), .A3(G244), .A4(new_n259), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT4), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n257), .A2(KEYINPUT4), .A3(G244), .A4(new_n259), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n257), .A2(G250), .A3(G1698), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n351), .A2(new_n352), .A3(new_n291), .A4(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n348), .B1(new_n354), .B2(new_n250), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n341), .A2(new_n345), .B1(new_n355), .B2(G169), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n250), .ZN(new_n357));
  INV_X1    g0157(.A(new_n348), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n357), .A2(new_n315), .A3(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT78), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n355), .A2(KEYINPUT78), .A3(new_n315), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n356), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n355), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(G200), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n341), .A2(new_n345), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n355), .A2(G190), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT77), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT77), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n365), .A2(new_n366), .A3(new_n370), .A4(new_n367), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n363), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  AND2_X1   g0172(.A1(KEYINPUT69), .A2(G107), .ZN(new_n373));
  NOR2_X1   g0173(.A1(KEYINPUT69), .A2(G107), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(G87), .A2(G97), .ZN(new_n376));
  NAND3_X1  g0176(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n375), .A2(new_n376), .B1(new_n208), .B2(new_n377), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n252), .A2(new_n254), .A3(new_n208), .A4(G68), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT19), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n208), .A2(G33), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n380), .B1(new_n381), .B2(new_n292), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n280), .B1(new_n378), .B2(new_n383), .ZN(new_n384));
  XNOR2_X1  g0184(.A(KEYINPUT15), .B(G87), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n278), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n343), .A2(new_n386), .A3(new_n283), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n384), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT81), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT81), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n384), .A2(new_n393), .A3(new_n389), .A4(new_n390), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n211), .A2(G45), .ZN(new_n396));
  AND3_X1   g0196(.A1(new_n249), .A2(G250), .A3(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT79), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n398), .B1(new_n268), .B2(new_n396), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n249), .A2(KEYINPUT79), .A3(G274), .A4(new_n263), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n397), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n252), .A2(new_n254), .A3(G244), .A4(G1698), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n252), .A2(new_n254), .A3(G238), .A4(new_n259), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n402), .B(new_n403), .C1(new_n251), .C2(new_n285), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n250), .ZN(new_n405));
  AND3_X1   g0205(.A1(new_n401), .A2(new_n405), .A3(new_n315), .ZN(new_n406));
  AOI21_X1  g0206(.A(G169), .B1(new_n401), .B2(new_n405), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n343), .A2(G87), .A3(new_n283), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n384), .A2(new_n389), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n401), .A2(new_n405), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n410), .B1(G200), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n411), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(G190), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n395), .A2(new_n408), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n319), .A2(new_n325), .A3(new_n372), .A4(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n278), .A2(new_n218), .ZN(new_n417));
  XNOR2_X1  g0217(.A(new_n417), .B(KEYINPUT12), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n332), .A2(G50), .B1(G20), .B2(new_n218), .ZN(new_n419));
  INV_X1    g0219(.A(G77), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n419), .B1(new_n420), .B2(new_n381), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n421), .A2(KEYINPUT11), .A3(new_n280), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(KEYINPUT11), .B1(new_n421), .B2(new_n280), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n281), .A2(new_n282), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n426), .B(G68), .C1(G1), .C2(new_n208), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT67), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n211), .B(KEYINPUT67), .C1(G41), .C2(G45), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n431), .A2(G238), .A3(new_n249), .A4(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n429), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n434), .A2(new_n249), .A3(G274), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n252), .A2(new_n254), .A3(G232), .A4(G1698), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n252), .A2(new_n254), .A3(G226), .A4(new_n259), .ZN(new_n438));
  NAND2_X1  g0238(.A1(G33), .A2(G97), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n250), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT13), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n436), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n442), .B1(new_n436), .B2(new_n441), .ZN(new_n445));
  OAI21_X1  g0245(.A(G169), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT14), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n436), .A2(new_n441), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT13), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n443), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n451), .A2(KEYINPUT14), .A3(G169), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT73), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n443), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n436), .A2(new_n441), .A3(KEYINPUT73), .A4(new_n442), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n455), .A2(new_n450), .A3(G179), .A4(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n428), .B1(new_n453), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  AND3_X1   g0259(.A1(new_n455), .A2(new_n456), .A3(new_n450), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G190), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n451), .A2(G200), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n461), .A2(new_n428), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n431), .A2(new_n249), .A3(new_n432), .ZN(new_n465));
  INV_X1    g0265(.A(G226), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n435), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n257), .A2(G222), .A3(new_n259), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n257), .A2(G1698), .ZN(new_n469));
  INV_X1    g0269(.A(G223), .ZN(new_n470));
  OAI221_X1 g0270(.A(new_n468), .B1(new_n221), .B2(new_n257), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n467), .B1(new_n471), .B2(new_n250), .ZN(new_n472));
  INV_X1    g0272(.A(G200), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n474), .B1(G190), .B2(new_n472), .ZN(new_n475));
  OAI21_X1  g0275(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n476));
  INV_X1    g0276(.A(G150), .ZN(new_n477));
  INV_X1    g0277(.A(new_n332), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  XNOR2_X1  g0279(.A(KEYINPUT8), .B(G58), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT68), .ZN(new_n481));
  XNOR2_X1  g0281(.A(new_n480), .B(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n381), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n479), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(new_n289), .ZN(new_n485));
  INV_X1    g0285(.A(G50), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n278), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n289), .B1(G1), .B2(new_n208), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n487), .B1(new_n488), .B2(new_n486), .ZN(new_n489));
  OAI21_X1  g0289(.A(KEYINPUT9), .B1(new_n485), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT9), .ZN(new_n491));
  INV_X1    g0291(.A(new_n489), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n491), .B(new_n492), .C1(new_n484), .C2(new_n289), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n475), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT10), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n472), .A2(G190), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n497), .B(KEYINPUT72), .C1(new_n473), .C2(new_n472), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n495), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n475), .B(new_n494), .C1(KEYINPUT72), .C2(KEYINPUT10), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n485), .A2(new_n489), .ZN(new_n502));
  INV_X1    g0302(.A(new_n472), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n502), .B1(new_n306), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n472), .A2(new_n315), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n426), .B(G77), .C1(G1), .C2(new_n208), .ZN(new_n508));
  XNOR2_X1  g0308(.A(new_n480), .B(KEYINPUT70), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n509), .A2(new_n478), .ZN(new_n510));
  OAI22_X1  g0310(.A1(new_n208), .A2(new_n221), .B1(new_n385), .B2(new_n381), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n280), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n508), .B(new_n512), .C1(new_n222), .C2(new_n387), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n257), .A2(G232), .A3(new_n259), .ZN(new_n514));
  OAI221_X1 g0314(.A(new_n514), .B1(new_n257), .B2(new_n375), .C1(new_n469), .C2(new_n219), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n250), .ZN(new_n516));
  INV_X1    g0316(.A(new_n435), .ZN(new_n517));
  INV_X1    g0317(.A(new_n465), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n517), .B1(new_n518), .B2(G244), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(G190), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n473), .B1(new_n516), .B2(new_n519), .ZN(new_n523));
  OR3_X1    g0323(.A1(new_n513), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n516), .A2(new_n315), .A3(new_n519), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n520), .A2(new_n306), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n513), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  NOR4_X1   g0328(.A1(new_n464), .A2(new_n501), .A3(new_n507), .A4(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(G87), .ZN(new_n530));
  OAI22_X1  g0330(.A1(new_n469), .A2(new_n466), .B1(new_n251), .B2(new_n530), .ZN(new_n531));
  NOR3_X1   g0331(.A1(new_n336), .A2(new_n470), .A3(G1698), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n250), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n517), .B1(new_n518), .B2(G232), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G169), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(new_n315), .B2(new_n535), .ZN(new_n537));
  INV_X1    g0337(.A(G58), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n538), .A2(new_n218), .ZN(new_n539));
  OAI21_X1  g0339(.A(G20), .B1(new_n539), .B2(new_n201), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n332), .A2(G159), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n542), .B1(new_n338), .B2(G68), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n280), .B1(new_n543), .B2(KEYINPUT16), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT74), .ZN(new_n545));
  AND3_X1   g0345(.A1(new_n252), .A2(new_n254), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n545), .B1(new_n252), .B2(new_n254), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(KEYINPUT7), .B1(new_n548), .B2(new_n208), .ZN(new_n549));
  NOR3_X1   g0349(.A1(new_n257), .A2(new_n334), .A3(G20), .ZN(new_n550));
  OAI21_X1  g0350(.A(G68), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n542), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n551), .A2(KEYINPUT75), .A3(KEYINPUT16), .A4(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n253), .A2(G33), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n555));
  OAI21_X1  g0355(.A(KEYINPUT74), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n252), .A2(new_n254), .A3(new_n545), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n556), .A2(new_n208), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n550), .B1(new_n558), .B2(new_n334), .ZN(new_n559));
  OAI211_X1 g0359(.A(KEYINPUT16), .B(new_n552), .C1(new_n559), .C2(new_n218), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT75), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n544), .B1(new_n553), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n482), .A2(new_n488), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n278), .B2(new_n482), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n537), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT18), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT18), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n537), .B(new_n569), .C1(new_n563), .C2(new_n566), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n544), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n560), .A2(new_n561), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n560), .A2(new_n561), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n533), .A2(G190), .A3(new_n534), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n565), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n473), .B1(new_n533), .B2(new_n534), .ZN(new_n578));
  NOR3_X1   g0378(.A1(new_n577), .A2(KEYINPUT17), .A3(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n575), .A2(KEYINPUT76), .A3(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT76), .ZN(new_n581));
  INV_X1    g0381(.A(new_n578), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT17), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n582), .A2(new_n583), .A3(new_n565), .A4(new_n576), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n581), .B1(new_n563), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n582), .A2(new_n565), .A3(new_n576), .ZN(new_n586));
  OAI21_X1  g0386(.A(KEYINPUT17), .B1(new_n563), .B2(new_n586), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n580), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n571), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n529), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n252), .A2(new_n254), .A3(G257), .A4(G1698), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n252), .A2(new_n254), .A3(G250), .A4(new_n259), .ZN(new_n592));
  NAND2_X1  g0392(.A1(G33), .A2(G294), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n594), .A2(new_n250), .B1(new_n272), .B2(G264), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n595), .A2(new_n315), .A3(new_n347), .ZN(new_n596));
  AOI21_X1  g0396(.A(G169), .B1(new_n595), .B2(new_n347), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(G107), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n278), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT86), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n600), .A2(new_n601), .A3(KEYINPUT25), .ZN(new_n602));
  XOR2_X1   g0402(.A(KEYINPUT86), .B(KEYINPUT25), .Z(new_n603));
  OAI221_X1 g0403(.A(new_n602), .B1(new_n600), .B2(new_n603), .C1(new_n344), .C2(new_n599), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(G116), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT80), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT80), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(G116), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n381), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT23), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n611), .A2(new_n599), .A3(G20), .ZN(new_n612));
  NAND2_X1  g0412(.A1(KEYINPUT85), .A2(KEYINPUT24), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n252), .A2(new_n254), .A3(new_n208), .A4(G87), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT22), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n257), .A2(KEYINPUT22), .A3(new_n208), .A4(G87), .ZN(new_n619));
  OAI21_X1  g0419(.A(KEYINPUT23), .B1(new_n339), .B2(new_n208), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n615), .A2(new_n618), .A3(new_n619), .A4(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(KEYINPUT85), .A2(KEYINPUT24), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n280), .B1(new_n621), .B2(new_n622), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n605), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n598), .A2(new_n626), .A3(KEYINPUT87), .ZN(new_n627));
  AOI21_X1  g0427(.A(KEYINPUT87), .B1(new_n598), .B2(new_n626), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT88), .ZN(new_n630));
  INV_X1    g0430(.A(new_n625), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n604), .B1(new_n631), .B2(new_n623), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n595), .A2(G190), .A3(new_n347), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n595), .A2(new_n347), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(G200), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n632), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n629), .A2(new_n630), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n598), .A2(new_n626), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT87), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n598), .A2(new_n626), .A3(KEYINPUT87), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(new_n641), .A3(new_n636), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(KEYINPUT88), .ZN(new_n643));
  AOI211_X1 g0443(.A(new_n416), .B(new_n590), .C1(new_n637), .C2(new_n643), .ZN(G372));
  INV_X1    g0444(.A(new_n590), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n313), .A2(new_n638), .A3(new_n318), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n646), .A2(new_n636), .A3(new_n372), .A4(new_n415), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n395), .A2(new_n408), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(KEYINPUT26), .B1(new_n363), .B2(new_n415), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n363), .A2(new_n415), .A3(KEYINPUT26), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n649), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n647), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n645), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n588), .ZN(new_n656));
  INV_X1    g0456(.A(new_n527), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n463), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n459), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n660), .A2(new_n568), .A3(new_n570), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT89), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n501), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n499), .A2(KEYINPUT89), .A3(new_n500), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n507), .B1(new_n661), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n655), .A2(new_n666), .ZN(G369));
  XNOR2_X1  g0467(.A(new_n323), .B(KEYINPUT84), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n313), .A2(new_n318), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n211), .A2(new_n208), .A3(G13), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n672), .A2(G213), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G343), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n298), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT90), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n670), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n319), .B2(new_n678), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(G330), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n637), .A2(new_n643), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n632), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n630), .B1(new_n629), .B2(new_n636), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n642), .A2(KEYINPUT88), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n675), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n638), .A2(new_n675), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n683), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n681), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n682), .A2(new_n669), .A3(new_n675), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n598), .A2(new_n626), .A3(new_n675), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n692), .A2(new_n695), .ZN(G399));
  INV_X1    g0496(.A(new_n214), .ZN(new_n697));
  OR3_X1    g0497(.A1(new_n697), .A2(KEYINPUT91), .A3(G41), .ZN(new_n698));
  OAI21_X1  g0498(.A(KEYINPUT91), .B1(new_n697), .B2(G41), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n376), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n339), .A2(G116), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n700), .A2(G1), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n205), .B2(new_n700), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT28), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n676), .B1(new_n647), .B2(new_n653), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT29), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n372), .A2(new_n415), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n629), .A2(new_n313), .A3(new_n318), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(new_n636), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n652), .B1(new_n650), .B2(KEYINPUT92), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n361), .A2(new_n362), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n412), .A2(new_n414), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n329), .B1(new_n327), .B2(new_n326), .ZN(new_n715));
  OAI22_X1  g0515(.A1(new_n715), .A2(new_n208), .B1(new_n420), .B2(new_n478), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n375), .B1(new_n335), .B2(new_n337), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n280), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n345), .ZN(new_n719));
  AOI22_X1  g0519(.A1(new_n364), .A2(new_n306), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n648), .A2(new_n713), .A3(new_n714), .A4(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT26), .ZN(new_n722));
  OR3_X1    g0522(.A1(new_n721), .A2(KEYINPUT92), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n649), .B1(new_n712), .B2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT93), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n711), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  AOI211_X1 g0526(.A(KEYINPUT93), .B(new_n649), .C1(new_n712), .C2(new_n723), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n675), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n708), .B1(new_n728), .B2(KEYINPUT29), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n316), .A2(new_n595), .A3(new_n355), .A4(new_n413), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT30), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n413), .A2(new_n595), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n733), .A2(KEYINPUT30), .A3(new_n355), .A4(new_n316), .ZN(new_n734));
  INV_X1    g0534(.A(new_n305), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n364), .A2(new_n315), .A3(new_n634), .A4(new_n411), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n732), .B(new_n734), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n737), .A2(KEYINPUT31), .A3(new_n676), .ZN(new_n738));
  AOI21_X1  g0538(.A(KEYINPUT31), .B1(new_n737), .B2(new_n676), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(new_n686), .B2(new_n416), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G330), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n729), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n705), .B1(new_n744), .B2(G1), .ZN(G364));
  INV_X1    g0545(.A(new_n700), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n277), .A2(G20), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G45), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n211), .B1(new_n749), .B2(KEYINPUT94), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(KEYINPUT94), .B2(new_n749), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n746), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n752), .B1(new_n680), .B2(G330), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(G330), .B2(new_n680), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT95), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n697), .A2(new_n336), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G355), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n758), .B1(G116), .B2(new_n214), .ZN(new_n759));
  INV_X1    g0559(.A(new_n548), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n697), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n762), .B1(new_n262), .B2(new_n206), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n243), .A2(new_n262), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n759), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G13), .A2(G33), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n207), .B1(G20), .B2(new_n306), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n752), .B1(new_n765), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n208), .A2(new_n315), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n773), .A2(G190), .A3(new_n473), .ZN(new_n774));
  INV_X1    g0574(.A(G322), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G190), .A2(G200), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n773), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G311), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n336), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n208), .A2(G179), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(new_n777), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n776), .B(new_n780), .C1(G329), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n773), .A2(G200), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G190), .ZN(new_n786));
  INV_X1    g0586(.A(G317), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(KEYINPUT33), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n787), .A2(KEYINPUT33), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n786), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n781), .A2(G190), .A3(G200), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n315), .A2(new_n473), .A3(G190), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G20), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n792), .A2(G303), .B1(new_n794), .B2(G294), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n785), .A2(new_n521), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n781), .A2(new_n521), .A3(G200), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n796), .A2(G326), .B1(new_n798), .B2(G283), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n784), .A2(new_n790), .A3(new_n795), .A4(new_n799), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n794), .B(KEYINPUT98), .Z(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n292), .ZN(new_n803));
  INV_X1    g0603(.A(new_n774), .ZN(new_n804));
  INV_X1    g0604(.A(new_n778), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n804), .A2(G58), .B1(new_n805), .B2(new_n222), .ZN(new_n806));
  INV_X1    g0606(.A(new_n796), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n806), .B1(new_n486), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G159), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n782), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g0610(.A(KEYINPUT96), .B(KEYINPUT32), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  INV_X1    g0613(.A(new_n786), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n814), .B2(new_n218), .ZN(new_n815));
  OR4_X1    g0615(.A1(new_n803), .A2(new_n808), .A3(new_n812), .A4(new_n815), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n257), .B1(new_n797), .B2(new_n599), .C1(new_n530), .C2(new_n791), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT97), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n800), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT99), .ZN(new_n820));
  OR2_X1    g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n769), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(new_n819), .B2(new_n820), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n772), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n768), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n824), .B1(new_n680), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n756), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT100), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n827), .B(new_n828), .ZN(G396));
  NOR2_X1   g0629(.A1(new_n527), .A2(new_n676), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n513), .A2(new_n676), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n524), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n830), .B1(new_n832), .B2(new_n527), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n706), .A2(new_n833), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT102), .Z(new_n835));
  NOR2_X1   g0635(.A1(new_n528), .A2(new_n676), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n654), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n752), .B1(new_n838), .B2(new_n742), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n742), .B2(new_n838), .ZN(new_n840));
  INV_X1    g0640(.A(new_n752), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n769), .A2(new_n766), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n841), .B1(new_n420), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n285), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n796), .A2(G303), .B1(new_n805), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(G283), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n845), .B1(new_n846), .B2(new_n814), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n847), .B(KEYINPUT101), .Z(new_n848));
  INV_X1    g0648(.A(G294), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n336), .B1(new_n782), .B2(new_n779), .C1(new_n774), .C2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n791), .A2(new_n599), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n797), .A2(new_n530), .ZN(new_n852));
  NOR4_X1   g0652(.A1(new_n803), .A2(new_n850), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n548), .B1(G132), .B2(new_n783), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n798), .A2(G68), .B1(new_n794), .B2(G58), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n854), .B(new_n855), .C1(new_n486), .C2(new_n791), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT34), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n804), .A2(G143), .B1(new_n805), .B2(G159), .ZN(new_n858));
  INV_X1    g0658(.A(G137), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n858), .B1(new_n807), .B2(new_n859), .C1(new_n477), .C2(new_n814), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n856), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  OR2_X1    g0661(.A1(new_n860), .A2(new_n857), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n848), .A2(new_n853), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n843), .B1(new_n822), .B2(new_n863), .C1(new_n833), .C2(new_n767), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n840), .A2(new_n864), .ZN(G384));
  NOR3_X1   g0665(.A1(new_n205), .A2(new_n221), .A3(new_n539), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(new_n486), .B2(G68), .ZN(new_n867));
  NOR3_X1   g0667(.A1(new_n867), .A2(new_n211), .A3(G13), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n868), .B(KEYINPUT104), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n331), .A2(KEYINPUT35), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n331), .A2(KEYINPUT35), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n870), .A2(G116), .A3(new_n209), .A4(new_n871), .ZN(new_n872));
  XOR2_X1   g0672(.A(new_n872), .B(KEYINPUT36), .Z(new_n873));
  INV_X1    g0673(.A(KEYINPUT103), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n869), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(new_n874), .B2(new_n873), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT106), .ZN(new_n877));
  AOI22_X1  g0677(.A1(new_n448), .A2(new_n452), .B1(new_n460), .B2(G179), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n463), .B(new_n877), .C1(new_n878), .C2(new_n428), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n675), .B1(new_n425), .B2(new_n427), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT14), .B1(new_n451), .B2(G169), .ZN(new_n883));
  AOI211_X1 g0683(.A(new_n447), .B(new_n306), .C1(new_n450), .C2(new_n443), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n457), .B(new_n880), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n886), .B(new_n463), .C1(new_n458), .C2(new_n877), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n882), .A2(new_n887), .A3(new_n833), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n682), .A2(new_n670), .A3(new_n709), .A4(new_n675), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n888), .B1(new_n889), .B2(new_n740), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n553), .A2(new_n562), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n552), .B1(new_n559), .B2(new_n218), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT16), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n289), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n566), .B1(new_n891), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n674), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n571), .B2(new_n588), .ZN(new_n898));
  OAI22_X1  g0698(.A1(new_n895), .A2(new_n896), .B1(new_n563), .B2(new_n586), .ZN(new_n899));
  INV_X1    g0699(.A(new_n537), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n895), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(KEYINPUT37), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n563), .A2(new_n586), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n674), .B1(new_n563), .B2(new_n566), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT37), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n903), .A2(new_n567), .A3(new_n904), .A4(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n898), .A2(new_n907), .A3(KEYINPUT38), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT38), .B1(new_n898), .B2(new_n907), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n890), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  XNOR2_X1  g0710(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(KEYINPUT109), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT109), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n910), .A2(new_n915), .A3(new_n912), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n898), .A2(new_n907), .A3(KEYINPUT38), .ZN(new_n917));
  INV_X1    g0717(.A(new_n904), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n571), .B2(new_n588), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n903), .A2(new_n567), .A3(new_n904), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(KEYINPUT37), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n906), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n917), .B1(new_n923), .B2(KEYINPUT38), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n890), .A2(KEYINPUT40), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n914), .A2(new_n916), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n645), .A2(new_n741), .ZN(new_n928));
  OAI21_X1  g0728(.A(G330), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(new_n928), .B2(new_n927), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT38), .B1(new_n919), .B2(new_n922), .ZN(new_n931));
  NOR3_X1   g0731(.A1(new_n908), .A2(new_n931), .A3(KEYINPUT39), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT39), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n898), .A2(new_n907), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT38), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n933), .B1(new_n936), .B2(new_n917), .ZN(new_n937));
  OAI21_X1  g0737(.A(KEYINPUT107), .B1(new_n932), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n459), .A2(new_n676), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n917), .B(new_n933), .C1(new_n923), .C2(KEYINPUT38), .ZN(new_n940));
  OAI21_X1  g0740(.A(KEYINPUT39), .B1(new_n908), .B2(new_n909), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT107), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n938), .A2(new_n939), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n882), .A2(new_n887), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT105), .ZN(new_n946));
  INV_X1    g0746(.A(new_n830), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n837), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n836), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(new_n647), .B2(new_n653), .ZN(new_n950));
  OAI21_X1  g0750(.A(KEYINPUT105), .B1(new_n950), .B2(new_n830), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n945), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n936), .A2(new_n917), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n952), .A2(new_n953), .B1(new_n571), .B2(new_n896), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n944), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(KEYINPUT92), .B1(new_n721), .B2(new_n722), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n721), .A2(new_n722), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR3_X1   g0758(.A1(new_n721), .A2(KEYINPUT92), .A3(new_n722), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n648), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(KEYINPUT93), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n724), .A2(new_n725), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n961), .A2(new_n962), .A3(new_n711), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n707), .B1(new_n963), .B2(new_n675), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n645), .B1(new_n964), .B2(new_n708), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n666), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n955), .B(new_n966), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n930), .A2(new_n967), .B1(new_n211), .B2(new_n747), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n930), .A2(new_n967), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n876), .B1(new_n968), .B2(new_n969), .ZN(G367));
  OAI21_X1  g0770(.A(new_n372), .B1(new_n366), .B2(new_n675), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n363), .A2(new_n676), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n693), .A2(new_n974), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n975), .A2(KEYINPUT42), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n971), .A2(new_n629), .ZN(new_n977));
  INV_X1    g0777(.A(new_n363), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n676), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(new_n975), .B2(KEYINPUT42), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n676), .A2(new_n410), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n415), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n648), .B2(new_n981), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n976), .A2(new_n980), .B1(KEYINPUT43), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n983), .A2(KEYINPUT43), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n984), .B(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n691), .A2(new_n973), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n986), .B(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n700), .B(KEYINPUT41), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT44), .ZN(new_n990));
  NOR3_X1   g0790(.A1(new_n695), .A2(new_n990), .A3(new_n973), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n991), .A2(KEYINPUT110), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n990), .B1(new_n695), .B2(new_n973), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(KEYINPUT111), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT111), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n995), .B(new_n990), .C1(new_n695), .C2(new_n973), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n991), .A2(KEYINPUT110), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n992), .A2(new_n994), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n695), .A2(new_n973), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT45), .Z(new_n1000));
  NAND2_X1  g0800(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n691), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n319), .A2(new_n676), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n693), .B1(new_n689), .B2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(new_n681), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n743), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n998), .A2(new_n692), .A3(new_n1000), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1002), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n989), .B1(new_n1008), .B2(new_n744), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n751), .B(KEYINPUT112), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n988), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n770), .B1(new_n214), .B2(new_n385), .C1(new_n762), .C2(new_n239), .ZN(new_n1012));
  AND2_X1   g0812(.A1(new_n752), .A2(new_n1012), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n814), .A2(new_n809), .B1(new_n778), .B2(new_n486), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1014), .A2(KEYINPUT113), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n801), .A2(G68), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1014), .A2(KEYINPUT113), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n257), .B1(new_n774), .B2(new_n477), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(G137), .B2(new_n783), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n796), .A2(G143), .B1(new_n798), .B2(new_n222), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1020), .B(new_n1021), .C1(new_n538), .C2(new_n791), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n798), .A2(G97), .B1(new_n339), .B2(new_n794), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n807), .B2(new_n779), .C1(new_n849), .C2(new_n814), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n778), .A2(new_n846), .B1(new_n782), .B2(new_n787), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(G303), .B2(new_n804), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT46), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n791), .B2(new_n285), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n792), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1026), .A2(new_n548), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n1018), .A2(new_n1022), .B1(new_n1024), .B2(new_n1030), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT47), .Z(new_n1032));
  OAI221_X1 g0832(.A(new_n1013), .B1(new_n825), .B2(new_n983), .C1(new_n1032), .C2(new_n822), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1011), .A2(new_n1033), .ZN(G387));
  AOI22_X1  g0834(.A1(new_n804), .A2(G317), .B1(new_n805), .B2(G303), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n807), .B2(new_n775), .C1(new_n779), .C2(new_n814), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT48), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n792), .A2(G294), .B1(new_n794), .B2(G283), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT49), .Z(new_n1042));
  AOI21_X1  g0842(.A(new_n760), .B1(G326), .B2(new_n783), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n285), .B2(new_n797), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n774), .A2(new_n486), .B1(new_n782), .B2(new_n477), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(G68), .B2(new_n805), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n548), .B1(G97), .B2(new_n798), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n791), .A2(new_n221), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(G159), .B2(new_n796), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n482), .A2(new_n786), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1047), .A2(new_n1048), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n802), .A2(new_n385), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n769), .B1(new_n1045), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n702), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n757), .A2(new_n1056), .B1(new_n599), .B2(new_n697), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n509), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n486), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT50), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n262), .B1(new_n218), .B2(new_n420), .ZN(new_n1061));
  NOR3_X1   g0861(.A1(new_n1060), .A2(new_n1056), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n236), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n761), .B1(new_n1063), .B2(new_n262), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1057), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n841), .B1(new_n1065), .B2(new_n770), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1055), .B(new_n1066), .C1(new_n689), .C2(new_n825), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1010), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n746), .B1(new_n743), .B2(new_n1005), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n743), .A2(new_n1005), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1067), .B1(new_n1005), .B2(new_n1068), .C1(new_n1069), .C2(new_n1070), .ZN(G393));
  AND2_X1   g0871(.A1(new_n1008), .A2(new_n746), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n1002), .A2(new_n1007), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1072), .B1(new_n1006), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n974), .A2(new_n768), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n770), .B1(new_n292), .B2(new_n214), .C1(new_n762), .C2(new_n246), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT114), .ZN(new_n1077));
  OR2_X1    g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1078), .A2(new_n752), .A3(new_n1079), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n807), .A2(new_n787), .B1(new_n779), .B2(new_n774), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT52), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n336), .B1(new_n782), .B2(new_n775), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(G294), .B2(new_n805), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n786), .A2(G303), .B1(new_n798), .B2(G107), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n792), .A2(G283), .B1(new_n844), .B2(new_n794), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1082), .A2(new_n1084), .A3(new_n1085), .A4(new_n1086), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(G150), .A2(new_n796), .B1(new_n804), .B2(G159), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT51), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n791), .A2(new_n218), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n852), .B(new_n1090), .C1(G50), .C2(new_n786), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n801), .A2(G77), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n548), .B1(G143), .B2(new_n783), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1058), .A2(new_n805), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1087), .B1(new_n1089), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1080), .B1(new_n1096), .B2(new_n769), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1073), .A2(new_n1010), .B1(new_n1075), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1074), .A2(new_n1098), .ZN(G390));
  AND2_X1   g0899(.A1(new_n741), .A2(G330), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n945), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1100), .A2(new_n833), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n948), .A2(new_n951), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n939), .B1(new_n1103), .B2(new_n1101), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n938), .B2(new_n943), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n939), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n924), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n832), .A2(new_n527), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n947), .B1(new_n728), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1107), .B1(new_n1110), .B2(new_n1101), .ZN(new_n1111));
  OAI211_X1 g0911(.A(KEYINPUT115), .B(new_n1102), .C1(new_n1105), .C2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1103), .A2(new_n1101), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n1106), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n942), .B1(new_n940), .B2(new_n941), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1114), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1111), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1102), .A2(KEYINPUT115), .ZN(new_n1119));
  OR2_X1    g0919(.A1(new_n1102), .A2(KEYINPUT115), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1112), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1100), .A2(new_n645), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n666), .B(new_n1123), .C1(new_n729), .C2(new_n590), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT116), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n965), .A2(KEYINPUT116), .A3(new_n666), .A4(new_n1123), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1101), .B1(new_n1100), .B2(new_n833), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n833), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n742), .A2(new_n1129), .A3(new_n945), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1103), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n963), .A2(new_n675), .A3(new_n1108), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n945), .B1(new_n742), .B2(new_n1129), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1102), .A2(new_n1132), .A3(new_n1133), .A4(new_n947), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1126), .A2(new_n1127), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1122), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT117), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1138), .A2(new_n1139), .A3(new_n746), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1136), .B1(new_n1112), .B2(new_n1121), .ZN(new_n1141));
  OAI21_X1  g0941(.A(KEYINPUT117), .B1(new_n1141), .B2(new_n700), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1112), .A2(new_n1121), .A3(new_n1136), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1140), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n766), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n842), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n752), .B1(new_n482), .B2(new_n1146), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n778), .A2(new_n292), .B1(new_n782), .B2(new_n849), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n257), .B(new_n1148), .C1(G116), .C2(new_n804), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n792), .A2(G87), .B1(new_n798), .B2(G68), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n339), .A2(new_n786), .B1(new_n796), .B2(G283), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1149), .A2(new_n1092), .A3(new_n1150), .A4(new_n1151), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n786), .A2(G137), .B1(new_n796), .B2(G128), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT54), .B(G143), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n336), .B1(new_n805), .B2(new_n1155), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n804), .A2(G132), .B1(new_n783), .B2(G125), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n798), .A2(G50), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1153), .A2(new_n1156), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n791), .A2(new_n477), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT53), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n802), .B2(new_n809), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1152), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1147), .B1(new_n769), .B2(new_n1163), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n1122), .A2(new_n1010), .B1(new_n1145), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1144), .A2(new_n1165), .ZN(G378));
  INV_X1    g0966(.A(KEYINPUT121), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(new_n944), .B2(new_n954), .ZN(new_n1168));
  XOR2_X1   g0968(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1169));
  INV_X1    g0969(.A(new_n664), .ZN(new_n1170));
  AOI21_X1  g0970(.A(KEYINPUT89), .B1(new_n499), .B2(new_n500), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n506), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1172), .A2(KEYINPUT119), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT119), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n665), .B2(new_n506), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1169), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n502), .A2(new_n896), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1172), .A2(KEYINPUT119), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n665), .A2(new_n1174), .A3(new_n506), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1169), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  AND3_X1   g0981(.A1(new_n1176), .A2(new_n1177), .A3(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1177), .B1(new_n1176), .B2(new_n1181), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n926), .B2(G330), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n925), .A2(new_n924), .ZN(new_n1186));
  AND3_X1   g0986(.A1(new_n910), .A2(new_n915), .A3(new_n912), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n915), .B1(new_n910), .B2(new_n912), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1186), .B(G330), .C1(new_n1187), .C2(new_n1188), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1168), .B1(new_n1185), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n914), .A2(new_n916), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1193), .A2(new_n1184), .A3(G330), .A4(new_n1186), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1194), .B(new_n1195), .C1(new_n955), .C2(new_n1167), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1068), .B1(new_n1192), .B2(new_n1196), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n774), .A2(new_n599), .B1(new_n778), .B2(new_n385), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n760), .A2(G41), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1198), .B(new_n1200), .C1(G283), .C2(new_n783), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1049), .B1(G58), .B2(new_n798), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n786), .A2(G97), .B1(new_n796), .B2(G116), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1201), .A2(new_n1016), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT58), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n486), .B1(G33), .B2(G41), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1207), .B1(new_n1199), .B2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(G128), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n774), .A2(new_n1210), .B1(new_n778), .B2(new_n859), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(G132), .B2(new_n786), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n796), .A2(G125), .B1(new_n792), .B2(new_n1155), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(new_n802), .C2(new_n477), .ZN(new_n1214));
  XOR2_X1   g1014(.A(new_n1214), .B(KEYINPUT118), .Z(new_n1215));
  OR2_X1    g1015(.A1(new_n1215), .A2(KEYINPUT59), .ZN(new_n1216));
  AOI211_X1 g1016(.A(G33), .B(G41), .C1(new_n783), .C2(G124), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n809), .B2(new_n797), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n1215), .B2(KEYINPUT59), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1206), .B(new_n1209), .C1(new_n1216), .C2(new_n1219), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n752), .B1(G50), .B2(new_n1146), .C1(new_n1220), .C2(new_n822), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(new_n1190), .B2(new_n766), .ZN(new_n1222));
  XOR2_X1   g1022(.A(new_n1222), .B(KEYINPUT120), .Z(new_n1223));
  NOR2_X1   g1023(.A1(new_n1197), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n944), .A2(new_n954), .ZN(new_n1225));
  AND3_X1   g1025(.A1(new_n1195), .A2(new_n1194), .A3(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1225), .B1(new_n1195), .B2(new_n1194), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT57), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1138), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT122), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1229), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n955), .B1(new_n1185), .B2(new_n1191), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1195), .A2(new_n1194), .A3(new_n1225), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1235), .A2(KEYINPUT57), .A3(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1230), .B1(new_n1122), .B2(new_n1135), .ZN(new_n1238));
  OAI21_X1  g1038(.A(KEYINPUT122), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1234), .A2(new_n1239), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1138), .A2(new_n1231), .B1(new_n1192), .B2(new_n1196), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n746), .B1(new_n1241), .B2(KEYINPUT57), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1224), .B1(new_n1240), .B2(new_n1242), .ZN(G375));
  INV_X1    g1043(.A(new_n1053), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n774), .A2(new_n846), .B1(new_n778), .B2(new_n375), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n257), .B(new_n1245), .C1(G303), .C2(new_n783), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n796), .A2(G294), .B1(new_n798), .B2(G77), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n786), .A2(new_n844), .B1(new_n792), .B2(G97), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1244), .A2(new_n1246), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n796), .A2(G132), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(new_n809), .B2(new_n791), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n786), .B2(new_n1155), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n801), .A2(G50), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n548), .B1(G58), .B2(new_n798), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n778), .A2(new_n477), .B1(new_n782), .B2(new_n1210), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(G137), .B2(new_n804), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1252), .A2(new_n1253), .A3(new_n1254), .A4(new_n1256), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1249), .A2(new_n1257), .ZN(new_n1258));
  OAI221_X1 g1058(.A(new_n752), .B1(G68), .B2(new_n1146), .C1(new_n1258), .C2(new_n822), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(new_n945), .B2(new_n766), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(new_n1135), .B2(new_n1010), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1135), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1230), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n989), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1136), .A2(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1261), .B1(new_n1264), .B2(new_n1266), .ZN(G381));
  OR2_X1    g1067(.A1(G375), .A2(G378), .ZN(new_n1268));
  OR4_X1    g1068(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1269));
  OR4_X1    g1069(.A1(G387), .A2(new_n1268), .A3(new_n1269), .A4(G381), .ZN(G407));
  OAI211_X1 g1070(.A(G407), .B(G213), .C1(G343), .C2(new_n1268), .ZN(G409));
  INV_X1    g1071(.A(G390), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(G396), .B(G393), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT124), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1274), .B1(G387), .B2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1273), .B1(new_n1011), .B2(new_n1033), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1272), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(G387), .A2(new_n1274), .ZN(new_n1279));
  AOI21_X1  g1079(.A(KEYINPUT124), .B1(new_n1011), .B2(new_n1033), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1279), .B(G390), .C1(new_n1274), .C2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1278), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(G343), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(G213), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  OAI211_X1 g1086(.A(G378), .B(new_n1224), .C1(new_n1240), .C2(new_n1242), .ZN(new_n1287));
  AND2_X1   g1087(.A1(new_n1241), .A2(new_n1265), .ZN(new_n1288));
  NOR3_X1   g1088(.A1(new_n1226), .A2(new_n1227), .A3(new_n1068), .ZN(new_n1289));
  OR2_X1    g1089(.A1(new_n1289), .A2(new_n1223), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1144), .B(new_n1165), .C1(new_n1288), .C2(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1286), .B1(new_n1287), .B2(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1264), .B1(KEYINPUT60), .B2(new_n1136), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1230), .A2(KEYINPUT60), .A3(new_n1262), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n746), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1261), .B1(new_n1293), .B2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1296), .A2(new_n840), .A3(new_n864), .ZN(new_n1297));
  OAI211_X1 g1097(.A(G384), .B(new_n1261), .C1(new_n1293), .C2(new_n1295), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  AND3_X1   g1100(.A1(new_n1292), .A2(KEYINPUT62), .A3(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT62), .B1(new_n1292), .B2(new_n1300), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT125), .ZN(new_n1303));
  NOR3_X1   g1103(.A1(new_n1301), .A2(new_n1302), .A3(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1292), .A2(new_n1300), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT62), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1305), .A2(new_n1303), .A3(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1287), .A2(new_n1291), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(new_n1285), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1286), .A2(G2897), .ZN(new_n1310));
  AND3_X1   g1110(.A1(new_n1297), .A2(new_n1298), .A3(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1310), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(KEYINPUT61), .B1(new_n1309), .B2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1307), .A2(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1283), .B1(new_n1304), .B2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT61), .ZN(new_n1317));
  OR2_X1    g1117(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1318));
  OAI211_X1 g1118(.A(new_n1282), .B(new_n1317), .C1(new_n1318), .C2(new_n1292), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1292), .A2(KEYINPUT63), .A3(new_n1300), .ZN(new_n1321));
  AOI211_X1 g1121(.A(KEYINPUT123), .B(KEYINPUT63), .C1(new_n1292), .C2(new_n1300), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT123), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT63), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1323), .B1(new_n1305), .B2(new_n1324), .ZN(new_n1325));
  OAI211_X1 g1125(.A(new_n1320), .B(new_n1321), .C1(new_n1322), .C2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1316), .A2(new_n1326), .ZN(G405));
  INV_X1    g1127(.A(G378), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(G375), .A2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(new_n1299), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1300), .A2(G375), .A3(new_n1328), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1332), .A2(KEYINPUT126), .A3(new_n1287), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1287), .A2(KEYINPUT126), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1330), .A2(new_n1331), .A3(new_n1334), .ZN(new_n1335));
  AND3_X1   g1135(.A1(new_n1333), .A2(new_n1335), .A3(new_n1283), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1283), .B1(new_n1333), .B2(new_n1335), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1336), .A2(new_n1337), .ZN(G402));
endmodule


