//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 1 1 0 1 1 1 0 0 1 0 0 0 0 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 1 1 0 0 0 1 1 1 1 0 1 1 0 1 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(G353));
  NOR2_X1   g0006(.A1(G97), .A2(G107), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n214), .B1(new_n203), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G107), .ZN(new_n222));
  INV_X1    g0022(.A(G264), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n213), .B1(new_n218), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT65), .Z(new_n227));
  NOR2_X1   g0027(.A1(new_n213), .A2(G13), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT0), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n202), .A2(new_n203), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G50), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(G1), .A2(G13), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n234), .A2(new_n211), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  OAI211_X1 g0036(.A(new_n230), .B(new_n236), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n227), .A2(new_n237), .ZN(G361));
  XOR2_X1   g0038(.A(G238), .B(G244), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XOR2_X1   g0040(.A(KEYINPUT2), .B(G226), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT66), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n242), .B(new_n246), .ZN(G358));
  XNOR2_X1  g0047(.A(G68), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(new_n202), .ZN(new_n249));
  XOR2_X1   g0049(.A(KEYINPUT67), .B(G50), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(KEYINPUT69), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G87), .B(G97), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(KEYINPUT68), .ZN(new_n254));
  XOR2_X1   g0054(.A(G107), .B(G116), .Z(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n252), .B(new_n256), .ZN(G351));
  INV_X1    g0057(.A(G200), .ZN(new_n258));
  AND2_X1   g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G77), .ZN(new_n262));
  OR2_X1    g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G1698), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G222), .ZN(new_n268));
  INV_X1    g0068(.A(G223), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n265), .A2(G1698), .ZN(new_n270));
  OAI221_X1 g0070(.A(new_n262), .B1(new_n267), .B2(new_n268), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n272), .A2(G1), .A3(G13), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n210), .A2(G274), .ZN(new_n276));
  AND2_X1   g0076(.A1(KEYINPUT70), .A2(G41), .ZN(new_n277));
  NOR2_X1   g0077(.A1(KEYINPUT70), .A2(G41), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G45), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n276), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n282));
  AND2_X1   g0082(.A1(new_n273), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n281), .B1(G226), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n258), .B1(new_n275), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n275), .A2(new_n284), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n285), .B1(new_n287), .B2(G190), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT10), .B1(new_n285), .B2(KEYINPUT73), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT8), .B(G58), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n211), .A2(G33), .ZN(new_n291));
  INV_X1    g0091(.A(G150), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G20), .A2(G33), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  OAI22_X1  g0094(.A1(new_n290), .A2(new_n291), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n295), .B1(G20), .B2(new_n204), .ZN(new_n296));
  NAND3_X1  g0096(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n234), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G13), .ZN(new_n301));
  NOR3_X1   g0101(.A1(new_n301), .A2(new_n211), .A3(G1), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(new_n298), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n210), .A2(G20), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n303), .A2(G50), .A3(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n302), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n305), .B1(G50), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(KEYINPUT9), .B1(new_n300), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NOR3_X1   g0109(.A1(new_n300), .A2(KEYINPUT9), .A3(new_n307), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n288), .B(new_n289), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n285), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n275), .A2(G190), .A3(new_n284), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n312), .B(new_n313), .C1(new_n309), .C2(new_n310), .ZN(new_n314));
  INV_X1    g0114(.A(new_n289), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n303), .A2(KEYINPUT72), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT72), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(new_n302), .B2(new_n298), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n321), .A2(G77), .A3(new_n304), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(G77), .B2(new_n306), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n290), .A2(new_n294), .B1(new_n211), .B2(new_n220), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT15), .B(G87), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n325), .A2(new_n291), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n298), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  XOR2_X1   g0127(.A(new_n327), .B(KEYINPUT71), .Z(new_n328));
  OR2_X1    g0128(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n265), .A2(G232), .A3(new_n266), .ZN(new_n330));
  OAI221_X1 g0130(.A(new_n330), .B1(new_n222), .B2(new_n265), .C1(new_n270), .C2(new_n215), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n274), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n281), .B1(G244), .B2(new_n283), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G200), .ZN(new_n335));
  INV_X1    g0135(.A(G190), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n335), .B1(new_n336), .B2(new_n334), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n329), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n323), .A2(new_n328), .ZN(new_n339));
  INV_X1    g0139(.A(G169), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n334), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G179), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n332), .A2(new_n342), .A3(new_n333), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n338), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n287), .A2(new_n342), .ZN(new_n347));
  OAI221_X1 g0147(.A(new_n347), .B1(G169), .B2(new_n287), .C1(new_n300), .C2(new_n307), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n317), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT74), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT74), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n317), .A2(new_n346), .A3(new_n351), .A4(new_n348), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT14), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n265), .A2(G232), .A3(G1698), .ZN(new_n355));
  NAND2_X1  g0155(.A1(G33), .A2(G97), .ZN(new_n356));
  INV_X1    g0156(.A(G226), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n355), .B(new_n356), .C1(new_n267), .C2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n274), .ZN(new_n359));
  XOR2_X1   g0159(.A(KEYINPUT75), .B(KEYINPUT13), .Z(new_n360));
  AOI21_X1  g0160(.A(new_n281), .B1(G238), .B2(new_n283), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n360), .B1(new_n359), .B2(new_n361), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n354), .B(G169), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n359), .A2(new_n361), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT13), .ZN(new_n368));
  OAI211_X1 g0168(.A(G179), .B(new_n362), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n365), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n364), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n340), .B1(new_n371), .B2(new_n362), .ZN(new_n372));
  OAI21_X1  g0172(.A(KEYINPUT78), .B1(new_n372), .B2(new_n354), .ZN(new_n373));
  OAI21_X1  g0173(.A(G169), .B1(new_n363), .B2(new_n364), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT78), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n374), .A2(new_n375), .A3(KEYINPUT14), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n370), .B1(new_n373), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n294), .A2(new_n201), .ZN(new_n378));
  OAI22_X1  g0178(.A1(new_n291), .A2(new_n220), .B1(new_n211), .B2(G68), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n298), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  XNOR2_X1  g0180(.A(new_n380), .B(KEYINPUT11), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT77), .B1(new_n302), .B2(new_n203), .ZN(new_n382));
  XNOR2_X1  g0182(.A(new_n382), .B(KEYINPUT12), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  AND3_X1   g0184(.A1(new_n321), .A2(G68), .A3(new_n304), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n377), .A2(new_n386), .ZN(new_n387));
  OAI211_X1 g0187(.A(G190), .B(new_n362), .C1(new_n367), .C2(new_n368), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n386), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n258), .B1(new_n371), .B2(new_n362), .ZN(new_n390));
  OR2_X1    g0190(.A1(new_n390), .A2(KEYINPUT76), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(KEYINPUT76), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n389), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n387), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT16), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n263), .A2(new_n211), .A3(new_n264), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n263), .A2(KEYINPUT7), .A3(new_n211), .A4(new_n264), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n203), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(G58), .A2(G68), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT79), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(KEYINPUT79), .A2(G58), .A3(G68), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n403), .A2(new_n231), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(G20), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n293), .A2(G159), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n395), .B1(new_n400), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(KEYINPUT7), .B1(new_n261), .B2(new_n211), .ZN(new_n410));
  NOR4_X1   g0210(.A1(new_n259), .A2(new_n260), .A3(new_n397), .A4(G20), .ZN(new_n411));
  OAI21_X1  g0211(.A(G68), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n405), .A2(G20), .B1(G159), .B2(new_n293), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(KEYINPUT16), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n409), .A2(new_n414), .A3(new_n298), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n269), .A2(new_n266), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n357), .A2(G1698), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n416), .B(new_n417), .C1(new_n259), .C2(new_n260), .ZN(new_n418));
  NAND2_X1  g0218(.A1(G33), .A2(G87), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(G190), .B1(new_n420), .B2(new_n274), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT80), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n273), .A2(G232), .A3(new_n282), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n422), .B1(new_n281), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g0224(.A(KEYINPUT70), .B(G41), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n210), .B(G274), .C1(new_n425), .C2(G45), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n273), .A2(G232), .A3(new_n282), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n426), .A2(KEYINPUT80), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n421), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n426), .A2(new_n427), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n273), .B1(new_n418), .B2(new_n419), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n258), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n290), .B1(new_n210), .B2(G20), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n434), .A2(new_n303), .B1(new_n302), .B2(new_n290), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n415), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT17), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT82), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n415), .A2(new_n433), .A3(KEYINPUT82), .A4(new_n435), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n438), .B1(new_n442), .B2(KEYINPUT17), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT18), .ZN(new_n444));
  AOI21_X1  g0244(.A(G179), .B1(new_n420), .B2(new_n274), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n445), .A2(new_n424), .A3(new_n428), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT81), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n340), .B1(new_n430), .B2(new_n431), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n447), .B1(new_n446), .B2(new_n448), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n415), .A2(new_n435), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n444), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n446), .A2(new_n448), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT81), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n456));
  AND4_X1   g0256(.A1(new_n444), .A2(new_n452), .A3(new_n455), .A4(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n443), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n353), .A2(new_n394), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(KEYINPUT23), .B1(new_n211), .B2(G107), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT23), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n463), .A2(new_n222), .A3(G20), .ZN(new_n464));
  INV_X1    g0264(.A(G116), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n462), .B(new_n464), .C1(new_n465), .C2(new_n291), .ZN(new_n466));
  XNOR2_X1  g0266(.A(new_n466), .B(KEYINPUT88), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n265), .A2(new_n211), .ZN(new_n468));
  OAI21_X1  g0268(.A(KEYINPUT22), .B1(new_n468), .B2(new_n216), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT22), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n265), .A2(new_n470), .A3(new_n211), .A4(G87), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT24), .ZN(new_n473));
  AND3_X1   g0273(.A1(new_n467), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n473), .B1(new_n467), .B2(new_n472), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n298), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n210), .A2(G33), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n303), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n302), .A2(KEYINPUT25), .A3(new_n222), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(KEYINPUT25), .B1(new_n302), .B2(new_n222), .ZN(new_n481));
  OAI22_X1  g0281(.A1(new_n478), .A2(new_n222), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n476), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n265), .A2(G257), .A3(G1698), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G294), .ZN(new_n486));
  OAI211_X1 g0286(.A(G250), .B(new_n266), .C1(new_n259), .C2(new_n260), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n274), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT5), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n210), .B(G45), .C1(new_n490), .C2(G41), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n491), .B1(new_n425), .B2(new_n490), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n493), .A2(G264), .A3(new_n273), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n492), .A2(G274), .A3(new_n273), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n496), .A2(G179), .A3(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT89), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n488), .A2(new_n499), .A3(new_n274), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n500), .A2(new_n497), .A3(new_n494), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n499), .B1(new_n488), .B2(new_n274), .ZN(new_n502));
  OAI21_X1  g0302(.A(G169), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n498), .B1(new_n503), .B2(KEYINPUT90), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT90), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n489), .A2(KEYINPUT89), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n506), .A2(new_n500), .A3(new_n497), .A4(new_n494), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n505), .B1(new_n507), .B2(G169), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n484), .B1(new_n504), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n489), .A2(new_n494), .A3(new_n497), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n258), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n507), .B2(G190), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(new_n476), .A3(new_n483), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT21), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n265), .A2(G257), .A3(new_n266), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n261), .A2(G303), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n516), .B(new_n517), .C1(new_n270), .C2(new_n223), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n274), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n492), .A2(new_n274), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G270), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n519), .A2(new_n497), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G169), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n465), .B1(new_n210), .B2(G33), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n318), .A2(new_n320), .A3(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n301), .A2(G1), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n526), .A2(G20), .A3(new_n465), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(G33), .ZN(new_n529));
  AOI21_X1  g0329(.A(G20), .B1(new_n529), .B2(G97), .ZN(new_n530));
  INV_X1    g0330(.A(G283), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n530), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n465), .A2(G20), .ZN(new_n533));
  AND3_X1   g0333(.A1(new_n298), .A2(KEYINPUT86), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(KEYINPUT86), .B1(new_n298), .B2(new_n533), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n532), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT20), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI211_X1 g0338(.A(KEYINPUT20), .B(new_n532), .C1(new_n534), .C2(new_n535), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n528), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n515), .B1(new_n523), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n538), .A2(new_n539), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n542), .A2(new_n527), .A3(new_n525), .ZN(new_n543));
  INV_X1    g0343(.A(new_n522), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n543), .A2(new_n544), .A3(G179), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n543), .A2(KEYINPUT21), .A3(G169), .A4(new_n522), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n541), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n544), .A2(G190), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n522), .A2(G200), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n548), .A2(new_n540), .A3(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT87), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n548), .A2(new_n549), .A3(KEYINPUT87), .A4(new_n540), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n547), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n265), .A2(G238), .A3(new_n266), .ZN(new_n555));
  NAND2_X1  g0355(.A1(G33), .A2(G116), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n555), .B(new_n556), .C1(new_n270), .C2(new_n221), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n274), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n276), .A2(new_n280), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n217), .B1(new_n210), .B2(G45), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n273), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n562), .A2(new_n258), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n303), .A2(G87), .A3(new_n477), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT85), .ZN(new_n566));
  XNOR2_X1  g0366(.A(new_n565), .B(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT19), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n211), .B1(new_n356), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(G87), .B2(new_n208), .ZN(new_n570));
  INV_X1    g0370(.A(G97), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n568), .B1(new_n291), .B2(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n570), .B(new_n572), .C1(new_n468), .C2(new_n203), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n573), .A2(new_n298), .B1(new_n302), .B2(new_n325), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n558), .A2(new_n561), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n567), .B(new_n574), .C1(new_n575), .C2(new_n336), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(G169), .B1(new_n558), .B2(new_n561), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n578), .B1(new_n342), .B2(new_n562), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n574), .B1(new_n325), .B2(new_n478), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n564), .A2(new_n577), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n520), .A2(G257), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n497), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  OAI22_X1  g0384(.A1(new_n270), .A2(new_n217), .B1(new_n529), .B2(new_n531), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT4), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n265), .A2(G244), .A3(new_n266), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n587), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n589), .A2(KEYINPUT84), .A3(KEYINPUT4), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT84), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(new_n587), .B2(new_n586), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n342), .B(new_n584), .C1(new_n594), .C2(new_n273), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n478), .A2(G97), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(G97), .B2(new_n302), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(KEYINPUT83), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT83), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n596), .B(new_n599), .C1(G97), .C2(new_n302), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT6), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n571), .A2(new_n222), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n602), .B1(new_n603), .B2(new_n207), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n222), .A2(KEYINPUT6), .A3(G97), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n606), .A2(G20), .B1(G77), .B2(new_n293), .ZN(new_n607));
  OAI21_X1  g0407(.A(G107), .B1(new_n410), .B2(new_n411), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n298), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n601), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n273), .B1(new_n588), .B2(new_n593), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n340), .B1(new_n612), .B2(new_n583), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n595), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  OAI211_X1 g0414(.A(G190), .B(new_n584), .C1(new_n594), .C2(new_n273), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n598), .A2(new_n600), .B1(new_n609), .B2(new_n298), .ZN(new_n616));
  OAI21_X1  g0416(.A(G200), .B1(new_n612), .B2(new_n583), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n581), .A2(new_n614), .A3(new_n618), .ZN(new_n619));
  AND4_X1   g0419(.A1(new_n461), .A2(new_n514), .A3(new_n554), .A4(new_n619), .ZN(G372));
  INV_X1    g0420(.A(new_n348), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT92), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n622), .B1(new_n453), .B2(new_n457), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n452), .A2(new_n455), .A3(new_n456), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(KEYINPUT18), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n451), .A2(new_n444), .A3(new_n452), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(new_n626), .A3(KEYINPUT92), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n392), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n390), .A2(KEYINPUT76), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n386), .B(new_n388), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n387), .B1(new_n631), .B2(new_n345), .ZN(new_n632));
  INV_X1    g0432(.A(new_n443), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n628), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n621), .B1(new_n634), .B2(new_n317), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n595), .A2(new_n611), .A3(new_n613), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n636), .A2(KEYINPUT26), .A3(new_n581), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT26), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n575), .A2(new_n340), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n639), .B(new_n580), .C1(G179), .C2(new_n575), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n563), .B2(new_n576), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n638), .B1(new_n614), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n640), .ZN(new_n644));
  INV_X1    g0444(.A(new_n547), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT91), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n646), .B(new_n484), .C1(new_n504), .C2(new_n508), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n503), .A2(KEYINPUT90), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n507), .A2(new_n505), .A3(G169), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(new_n498), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n646), .B1(new_n651), .B2(new_n484), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n645), .B1(new_n648), .B2(new_n652), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n581), .A2(new_n614), .A3(new_n618), .A4(new_n513), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n644), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n635), .B1(new_n460), .B2(new_n656), .ZN(G369));
  NAND2_X1  g0457(.A1(new_n526), .A2(new_n211), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(G213), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(G343), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n540), .A2(new_n664), .ZN(new_n665));
  MUX2_X1   g0465(.A(new_n554), .B(new_n547), .S(new_n665), .Z(new_n666));
  NAND2_X1  g0466(.A1(new_n484), .A2(new_n663), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n514), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n651), .A2(new_n484), .A3(new_n663), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n666), .A2(G330), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  OR3_X1    g0472(.A1(new_n648), .A2(new_n652), .A3(new_n663), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n645), .A2(new_n663), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n514), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n672), .A2(new_n673), .A3(new_n675), .ZN(G399));
  INV_X1    g0476(.A(new_n228), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(new_n425), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR3_X1   g0479(.A1(new_n208), .A2(G87), .A3(G116), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G1), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n232), .B2(new_n679), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT28), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n653), .A2(new_n655), .ZN(new_n684));
  AOI22_X1  g0484(.A1(new_n637), .A2(new_n642), .B1(new_n580), .B2(new_n579), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n663), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT29), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n654), .B1(new_n509), .B2(new_n645), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n664), .B1(new_n644), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT29), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n514), .A2(new_n619), .A3(new_n554), .A4(new_n664), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT31), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n544), .A2(new_n562), .A3(G179), .A4(new_n496), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n612), .A2(new_n583), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(KEYINPUT30), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT30), .ZN(new_n699));
  INV_X1    g0499(.A(new_n697), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n699), .B1(new_n700), .B2(new_n695), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n544), .A2(new_n562), .A3(G179), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n700), .A2(new_n510), .A3(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n698), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n663), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n694), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n704), .A2(KEYINPUT31), .A3(new_n663), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G330), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n692), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT93), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n692), .A2(new_n709), .A3(KEYINPUT93), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n683), .B1(new_n714), .B2(G1), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT94), .ZN(G364));
  AND2_X1   g0516(.A1(new_n666), .A2(G330), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n301), .A2(G20), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n210), .B1(new_n718), .B2(G45), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  OR3_X1    g0520(.A1(new_n678), .A2(KEYINPUT95), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(KEYINPUT95), .B1(new_n678), .B2(new_n720), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n717), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n725), .B1(G330), .B2(new_n666), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n228), .A2(new_n265), .ZN(new_n727));
  INV_X1    g0527(.A(G355), .ZN(new_n728));
  OAI22_X1  g0528(.A1(new_n727), .A2(new_n728), .B1(G116), .B2(new_n228), .ZN(new_n729));
  OR2_X1    g0529(.A1(new_n251), .A2(new_n280), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n677), .A2(new_n265), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n732), .B1(new_n280), .B2(new_n233), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n729), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(G13), .A2(G33), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G20), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n234), .B1(G20), .B2(new_n340), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n724), .B1(new_n734), .B2(new_n741), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n742), .A2(KEYINPUT96), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n211), .A2(new_n342), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(G190), .A3(G200), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT97), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G326), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n211), .A2(new_n336), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n342), .A2(G200), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n211), .A2(G190), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G179), .A2(G200), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI22_X1  g0559(.A1(G322), .A2(new_n755), .B1(new_n759), .B2(G329), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n258), .A2(G179), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n752), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n753), .A2(new_n756), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI22_X1  g0565(.A1(G303), .A2(new_n763), .B1(new_n765), .B2(G311), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n211), .B1(new_n757), .B2(G190), .ZN(new_n767));
  INV_X1    g0567(.A(G294), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n756), .A2(new_n761), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n261), .B1(new_n767), .B2(new_n768), .C1(new_n531), .C2(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n744), .A2(new_n336), .A3(G200), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(KEYINPUT33), .B(G317), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n770), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND4_X1  g0574(.A1(new_n751), .A2(new_n760), .A3(new_n766), .A4(new_n774), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT102), .Z(new_n776));
  OAI22_X1  g0576(.A1(new_n754), .A2(new_n202), .B1(new_n764), .B2(new_n220), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n777), .B1(new_n750), .B2(G50), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT98), .ZN(new_n779));
  XOR2_X1   g0579(.A(KEYINPUT99), .B(G159), .Z(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n758), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT101), .ZN(new_n782));
  XNOR2_X1  g0582(.A(KEYINPUT100), .B(KEYINPUT32), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n763), .A2(G87), .ZN(new_n785));
  INV_X1    g0585(.A(new_n769), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n261), .B1(new_n786), .B2(G107), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n767), .A2(new_n571), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n788), .B1(G68), .B2(new_n772), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n784), .A2(new_n785), .A3(new_n787), .A4(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n776), .B1(new_n779), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n743), .B1(new_n739), .B2(new_n791), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n792), .B1(KEYINPUT96), .B2(new_n742), .C1(new_n666), .C2(new_n738), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n726), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(G396));
  INV_X1    g0595(.A(KEYINPUT104), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n329), .A2(new_n796), .A3(new_n341), .A4(new_n343), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n339), .B(new_n335), .C1(new_n336), .C2(new_n334), .ZN(new_n798));
  OAI21_X1  g0598(.A(KEYINPUT104), .B1(new_n339), .B2(new_n344), .ZN(new_n799));
  AND3_X1   g0599(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n686), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n329), .A2(new_n663), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n797), .A2(new_n799), .A3(new_n798), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n345), .A2(new_n663), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n801), .B1(new_n686), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n724), .B1(new_n806), .B2(new_n709), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n709), .B2(new_n806), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n740), .A2(new_n736), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n724), .B1(G77), .B2(new_n809), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n772), .A2(G283), .B1(new_n765), .B2(G116), .ZN(new_n811));
  INV_X1    g0611(.A(G303), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n749), .B2(new_n812), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT103), .Z(new_n814));
  NOR2_X1   g0614(.A1(new_n769), .A2(new_n216), .ZN(new_n815));
  NOR3_X1   g0615(.A1(new_n815), .A2(new_n788), .A3(new_n265), .ZN(new_n816));
  AOI22_X1  g0616(.A1(G294), .A2(new_n755), .B1(new_n759), .B2(G311), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n816), .B(new_n817), .C1(new_n222), .C2(new_n762), .ZN(new_n818));
  INV_X1    g0618(.A(new_n780), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n765), .A2(new_n819), .B1(new_n755), .B2(G143), .ZN(new_n820));
  INV_X1    g0620(.A(G137), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n820), .B1(new_n292), .B2(new_n771), .C1(new_n749), .C2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(KEYINPUT34), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n265), .B1(new_n762), .B2(new_n201), .ZN(new_n825));
  INV_X1    g0625(.A(G132), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n769), .A2(new_n203), .B1(new_n758), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n767), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n825), .B(new_n827), .C1(G58), .C2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT34), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n829), .B1(new_n822), .B2(new_n830), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n814), .A2(new_n818), .B1(new_n824), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n810), .B1(new_n832), .B2(new_n739), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n805), .B2(new_n736), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n808), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(G384));
  INV_X1    g0636(.A(new_n661), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n452), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT106), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT37), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n452), .A2(KEYINPUT106), .A3(new_n837), .ZN(new_n842));
  AND3_X1   g0642(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  AND3_X1   g0643(.A1(new_n440), .A2(new_n624), .A3(new_n441), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n440), .A2(new_n624), .A3(new_n441), .A4(new_n838), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n843), .A2(new_n844), .B1(KEYINPUT37), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n838), .B1(new_n443), .B2(new_n458), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT38), .ZN(new_n848));
  NOR3_X1   g0648(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n848), .B1(new_n846), .B2(new_n847), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n663), .B1(new_n797), .B2(new_n799), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(new_n686), .B2(new_n800), .ZN(new_n855));
  INV_X1    g0655(.A(new_n386), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n373), .A2(new_n376), .ZN(new_n857));
  INV_X1    g0657(.A(new_n370), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n856), .B(new_n663), .C1(new_n859), .C2(new_n393), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n856), .A2(new_n663), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n631), .B(new_n861), .C1(new_n377), .C2(new_n386), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  NOR3_X1   g0664(.A1(new_n853), .A2(new_n855), .A3(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n628), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n865), .B1(new_n866), .B2(new_n661), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n623), .A2(new_n443), .A3(new_n627), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n840), .A2(new_n842), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n624), .A2(KEYINPUT92), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n452), .A2(new_n455), .A3(new_n622), .A4(new_n456), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n871), .A2(new_n436), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(KEYINPUT37), .B1(new_n873), .B2(new_n869), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n843), .A2(new_n844), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT38), .B1(new_n870), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n849), .B1(new_n877), .B2(KEYINPUT107), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT107), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n869), .A2(new_n868), .B1(new_n874), .B2(new_n875), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n879), .B1(new_n880), .B2(KEYINPUT38), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT39), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n850), .A2(KEYINPUT39), .A3(new_n851), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR3_X1   g0684(.A1(new_n377), .A2(new_n386), .A3(new_n663), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n867), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n635), .B1(new_n692), .B2(new_n460), .ZN(new_n888));
  XOR2_X1   g0688(.A(new_n887), .B(new_n888), .Z(new_n889));
  NAND2_X1  g0689(.A1(new_n870), .A2(new_n876), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n890), .A2(KEYINPUT107), .A3(new_n848), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n881), .A2(new_n891), .A3(new_n850), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(KEYINPUT109), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT109), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n878), .A2(new_n894), .A3(new_n881), .ZN(new_n895));
  INV_X1    g0695(.A(new_n805), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n896), .B1(new_n860), .B2(new_n862), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n693), .A2(KEYINPUT31), .B1(new_n663), .B2(new_n704), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n707), .A2(KEYINPUT108), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT108), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n704), .A2(new_n900), .A3(KEYINPUT31), .A4(new_n663), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n897), .B(KEYINPUT40), .C1(new_n898), .C2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n893), .A2(new_n895), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n706), .A2(new_n899), .A3(new_n901), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n852), .A2(new_n906), .A3(new_n897), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT40), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n461), .A2(new_n906), .ZN(new_n911));
  OAI21_X1  g0711(.A(G330), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n910), .B2(new_n911), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n889), .A2(new_n913), .B1(new_n210), .B2(new_n718), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n889), .B2(new_n913), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n233), .A2(G77), .A3(new_n403), .A4(new_n404), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n201), .A2(G68), .ZN(new_n917));
  AOI211_X1 g0717(.A(new_n210), .B(G13), .C1(new_n916), .C2(new_n917), .ZN(new_n918));
  OR2_X1    g0718(.A1(new_n606), .A2(KEYINPUT35), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n606), .A2(KEYINPUT35), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n919), .A2(G116), .A3(new_n235), .A4(new_n920), .ZN(new_n921));
  XOR2_X1   g0721(.A(KEYINPUT105), .B(KEYINPUT36), .Z(new_n922));
  XNOR2_X1  g0722(.A(new_n921), .B(new_n922), .ZN(new_n923));
  OR3_X1    g0723(.A1(new_n915), .A2(new_n918), .A3(new_n923), .ZN(G367));
  NAND2_X1  g0724(.A1(new_n731), .A2(new_n245), .ZN(new_n925));
  INV_X1    g0725(.A(new_n325), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n741), .B1(new_n677), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n723), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n567), .A2(new_n574), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n663), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n581), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n640), .B2(new_n930), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT46), .B1(new_n763), .B2(G116), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT114), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n934), .B1(G311), .B2(new_n750), .ZN(new_n935));
  INV_X1    g0735(.A(G317), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n758), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n769), .A2(new_n571), .ZN(new_n938));
  AOI211_X1 g0738(.A(new_n937), .B(new_n938), .C1(G303), .C2(new_n755), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n261), .B1(new_n764), .B2(new_n531), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n763), .A2(KEYINPUT46), .A3(G116), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n768), .B2(new_n771), .ZN(new_n942));
  AOI211_X1 g0742(.A(new_n940), .B(new_n942), .C1(G107), .C2(new_n828), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n935), .A2(new_n939), .A3(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n767), .A2(new_n203), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(G150), .B2(new_n755), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT115), .ZN(new_n947));
  OAI22_X1  g0747(.A1(new_n764), .A2(new_n201), .B1(new_n758), .B2(new_n821), .ZN(new_n948));
  OAI221_X1 g0748(.A(new_n265), .B1(new_n762), .B2(new_n202), .C1(new_n780), .C2(new_n771), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n948), .B(new_n949), .C1(G77), .C2(new_n786), .ZN(new_n950));
  INV_X1    g0750(.A(G143), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n950), .B1(new_n951), .B2(new_n749), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n944), .B1(new_n947), .B2(new_n952), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n953), .B(KEYINPUT47), .Z(new_n954));
  OAI221_X1 g0754(.A(new_n928), .B1(new_n738), .B2(new_n932), .C1(new_n954), .C2(new_n740), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n614), .B(new_n618), .C1(new_n616), .C2(new_n664), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n636), .A2(new_n663), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n673), .A2(new_n675), .A3(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT45), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n959), .A2(new_n960), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT113), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n961), .A2(new_n962), .B1(new_n963), .B2(new_n671), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n958), .B1(new_n673), .B2(new_n675), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT44), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n671), .A2(new_n963), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n964), .B(new_n966), .C1(new_n963), .C2(new_n671), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n675), .B1(new_n670), .B2(new_n674), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n717), .B(new_n972), .Z(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(new_n712), .B2(new_n713), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT112), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n971), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AOI211_X1 g0776(.A(KEYINPUT112), .B(new_n973), .C1(new_n712), .C2(new_n713), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n714), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n678), .B(KEYINPUT41), .Z(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n720), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n932), .A2(KEYINPUT43), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT110), .Z(new_n983));
  INV_X1    g0783(.A(KEYINPUT111), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n983), .A2(new_n984), .B1(KEYINPUT43), .B2(new_n932), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n958), .A2(new_n514), .A3(new_n674), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n986), .A2(KEYINPUT42), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(KEYINPUT42), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n614), .B1(new_n956), .B2(new_n509), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n664), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n985), .B1(new_n987), .B2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n958), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n672), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n992), .B(new_n994), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n983), .A2(new_n984), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n995), .B(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n955), .B1(new_n981), .B2(new_n998), .ZN(G387));
  INV_X1    g0799(.A(new_n973), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n668), .A2(new_n669), .A3(new_n737), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n727), .A2(new_n680), .B1(G107), .B2(new_n228), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n242), .A2(new_n280), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n680), .ZN(new_n1004));
  AOI211_X1 g0804(.A(G45), .B(new_n1004), .C1(G68), .C2(G77), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n290), .A2(G50), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT50), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n732), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1002), .B1(new_n1003), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n724), .B1(new_n1009), .B2(new_n741), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n750), .A2(G159), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n762), .A2(new_n220), .B1(new_n764), .B2(new_n203), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n754), .A2(new_n201), .B1(new_n758), .B2(new_n292), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n767), .A2(new_n325), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n290), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n261), .B(new_n938), .C1(new_n1017), .C2(new_n772), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1011), .A2(new_n1014), .A3(new_n1016), .A4(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n265), .B1(new_n759), .B2(G326), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n762), .A2(new_n768), .B1(new_n767), .B2(new_n531), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G317), .A2(new_n755), .B1(new_n765), .B2(G303), .ZN(new_n1022));
  INV_X1    g0822(.A(G311), .ZN(new_n1023));
  INV_X1    g0823(.A(G322), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1022), .B1(new_n1023), .B2(new_n771), .C1(new_n749), .C2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT48), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1021), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n1026), .B2(new_n1025), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT49), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1020), .B1(new_n465), .B2(new_n769), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1019), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1010), .B1(new_n1032), .B2(new_n739), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n1000), .A2(new_n720), .B1(new_n1001), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n714), .A2(new_n1000), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n678), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n714), .A2(new_n1000), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1034), .B1(new_n1036), .B2(new_n1037), .ZN(G393));
  INV_X1    g0838(.A(new_n971), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n679), .B1(new_n1039), .B2(new_n1035), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n977), .B2(new_n976), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n749), .A2(new_n936), .B1(new_n1023), .B2(new_n754), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT52), .Z(new_n1043));
  AOI22_X1  g0843(.A1(G294), .A2(new_n765), .B1(new_n759), .B2(G322), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n531), .B2(new_n762), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n265), .B1(new_n786), .B2(G107), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n465), .B2(new_n767), .C1(new_n812), .C2(new_n771), .ZN(new_n1047));
  NOR3_X1   g0847(.A1(new_n1043), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(G159), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n749), .A2(new_n292), .B1(new_n1049), .B2(new_n754), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT51), .Z(new_n1051));
  AOI22_X1  g0851(.A1(G68), .A2(new_n763), .B1(new_n765), .B2(new_n1017), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n951), .B2(new_n758), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n815), .A2(new_n261), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n828), .A2(G77), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1054), .B(new_n1055), .C1(new_n201), .C2(new_n771), .ZN(new_n1056));
  NOR3_X1   g0856(.A1(new_n1051), .A2(new_n1053), .A3(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n739), .B1(new_n1048), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n256), .A2(new_n731), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n741), .B1(G97), .B2(new_n677), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n723), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT117), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1058), .A2(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT118), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n993), .A2(KEYINPUT116), .A3(new_n737), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(KEYINPUT116), .B1(new_n993), .B2(new_n737), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n971), .B2(new_n720), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1041), .A2(new_n1069), .ZN(G390));
  INV_X1    g0870(.A(new_n885), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n855), .B2(new_n864), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n882), .B2(new_n883), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n664), .B(new_n800), .C1(new_n644), .C2(new_n689), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n854), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n885), .B1(new_n1076), .B2(new_n863), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n893), .A2(new_n895), .A3(new_n1077), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n897), .B(G330), .C1(new_n898), .C2(new_n902), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1079), .A2(KEYINPUT119), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n708), .A2(G330), .A3(new_n805), .A4(new_n863), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n1073), .A2(new_n1078), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT119), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1079), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n1073), .B2(new_n1078), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1087), .A2(new_n719), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n884), .A2(new_n736), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G132), .A2(new_n755), .B1(new_n759), .B2(G125), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1090), .B(new_n265), .C1(new_n201), .C2(new_n769), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n763), .A2(G150), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT53), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1091), .B(new_n1093), .C1(G128), .C2(new_n750), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(KEYINPUT54), .B(G143), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n764), .A2(new_n1095), .B1(new_n767), .B2(new_n1049), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(G137), .B2(new_n772), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT121), .Z(new_n1098));
  NAND2_X1  g0898(.A1(new_n750), .A2(G283), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n785), .A2(new_n261), .A3(new_n1055), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n769), .A2(new_n203), .B1(new_n758), .B2(new_n768), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n754), .A2(new_n465), .B1(new_n764), .B2(new_n571), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n771), .A2(new_n222), .ZN(new_n1103));
  NOR4_X1   g0903(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n1094), .A2(new_n1098), .B1(new_n1099), .B2(new_n1104), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n724), .B1(new_n1017), .B2(new_n809), .C1(new_n1105), .C2(new_n740), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1089), .A2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1088), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n707), .ZN(new_n1109));
  OAI211_X1 g0909(.A(G330), .B(new_n805), .C1(new_n898), .C2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n864), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n1079), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n855), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  OAI211_X1 g0914(.A(G330), .B(new_n805), .C1(new_n898), .C2(new_n902), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n864), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1081), .A2(new_n1116), .A3(new_n1075), .A4(new_n1074), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n461), .A2(new_n906), .A3(G330), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1119), .B(new_n635), .C1(new_n692), .C2(new_n460), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n679), .B1(new_n1087), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1120), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1125));
  AND3_X1   g0925(.A1(new_n1123), .A2(KEYINPUT120), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(KEYINPUT120), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1108), .B1(new_n1126), .B2(new_n1127), .ZN(G378));
  OAI21_X1  g0928(.A(new_n724), .B1(G50), .B2(new_n809), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n317), .A2(new_n348), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n300), .A2(new_n307), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1132), .A2(new_n661), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1130), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1136), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1130), .ZN(new_n1139));
  NOR3_X1   g0939(.A1(new_n1138), .A2(new_n1134), .A3(new_n1139), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT123), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1142), .A2(new_n736), .ZN(new_n1143));
  INV_X1    g0943(.A(G41), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n529), .B(new_n1144), .C1(new_n780), .C2(new_n769), .ZN(new_n1145));
  INV_X1    g0945(.A(G128), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n1146), .A2(new_n754), .B1(new_n762), .B2(new_n1095), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(G137), .B2(new_n765), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n772), .A2(G132), .B1(new_n828), .B2(G150), .ZN(new_n1149));
  INV_X1    g0949(.A(G125), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1148), .B(new_n1149), .C1(new_n1150), .C2(new_n749), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n1151), .A2(KEYINPUT59), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n1145), .B(new_n1152), .C1(G124), .C2(new_n759), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1153), .B1(KEYINPUT59), .B2(new_n1151), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n265), .A2(new_n425), .ZN(new_n1155));
  AOI211_X1 g0955(.A(G50), .B(new_n1155), .C1(new_n529), .C2(new_n1144), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n1156), .B(KEYINPUT122), .Z(new_n1157));
  NAND2_X1  g0957(.A1(new_n750), .A2(G116), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n769), .A2(new_n202), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n754), .A2(new_n222), .B1(new_n764), .B2(new_n325), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1159), .B(new_n1160), .C1(G283), .C2(new_n759), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n772), .A2(G97), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1155), .B1(new_n220), .B2(new_n762), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1163), .A2(new_n945), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1158), .A2(new_n1161), .A3(new_n1162), .A4(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1157), .B1(new_n1166), .B2(KEYINPUT58), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1154), .B(new_n1167), .C1(KEYINPUT58), .C2(new_n1166), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n1129), .B(new_n1143), .C1(new_n739), .C2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n905), .A2(G330), .A3(new_n909), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n1141), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1142), .A2(new_n905), .A3(G330), .A4(new_n909), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n887), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1171), .A2(new_n887), .A3(new_n1172), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1169), .B1(new_n1177), .B2(new_n720), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1125), .A2(new_n1121), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1179), .A2(new_n1175), .A3(KEYINPUT57), .A4(new_n1176), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1180), .A2(KEYINPUT124), .A3(new_n678), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1179), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT57), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1181), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(KEYINPUT124), .B1(new_n1180), .B2(new_n678), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1178), .B1(new_n1185), .B2(new_n1186), .ZN(G375));
  NOR2_X1   g0987(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1188));
  NOR3_X1   g0988(.A1(new_n1188), .A2(new_n1124), .A3(new_n979), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1189), .B(KEYINPUT125), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n864), .A2(new_n735), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n724), .B1(G68), .B2(new_n809), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n265), .B(new_n1015), .C1(G77), .C2(new_n786), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n762), .A2(new_n571), .B1(new_n764), .B2(new_n222), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n754), .A2(new_n531), .B1(new_n758), .B2(new_n812), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1193), .B(new_n1196), .C1(new_n465), .C2(new_n771), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n749), .A2(new_n768), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n749), .A2(new_n826), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n771), .A2(new_n1095), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(new_n1200), .A2(new_n1159), .A3(new_n261), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(G159), .A2(new_n763), .B1(new_n759), .B2(G128), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(G137), .A2(new_n755), .B1(new_n765), .B2(G150), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n828), .A2(G50), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n1197), .A2(new_n1198), .B1(new_n1199), .B2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1192), .B1(new_n1206), .B2(new_n739), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n1118), .A2(new_n720), .B1(new_n1191), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1190), .A2(new_n1208), .ZN(G381));
  NAND2_X1  g1009(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n1108), .ZN(new_n1211));
  INV_X1    g1011(.A(G390), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1212), .A2(new_n1190), .A3(new_n1213), .A4(new_n1208), .ZN(new_n1214));
  OR4_X1    g1014(.A1(G387), .A2(G375), .A3(new_n1211), .A4(new_n1214), .ZN(G407));
  INV_X1    g1015(.A(new_n1211), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n662), .A2(G213), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1219));
  OAI211_X1 g1019(.A(G407), .B(G213), .C1(G375), .C2(new_n1219), .ZN(G409));
  OAI211_X1 g1020(.A(G378), .B(new_n1178), .C1(new_n1185), .C2(new_n1186), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1178), .B1(new_n979), .B2(new_n1182), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n1216), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1221), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n1217), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1122), .A2(KEYINPUT60), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n679), .B1(new_n1226), .B2(new_n1188), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n1188), .B2(new_n1226), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1228), .A2(G384), .A3(new_n1208), .ZN(new_n1229));
  AOI21_X1  g1029(.A(G384), .B1(new_n1228), .B2(new_n1208), .ZN(new_n1230));
  OAI211_X1 g1030(.A(G2897), .B(new_n1218), .C1(new_n1229), .C2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1230), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1228), .A2(G384), .A3(new_n1208), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1218), .A2(G2897), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1232), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1231), .A2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(KEYINPUT61), .B1(new_n1225), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT63), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1238), .B1(new_n1225), .B2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(KEYINPUT126), .B1(G387), .B2(new_n1212), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(G393), .B(new_n794), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1035), .A2(KEYINPUT112), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n974), .A2(new_n975), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1245), .A2(new_n1246), .A3(new_n971), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n979), .B1(new_n1247), .B2(new_n714), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n997), .B1(new_n1248), .B2(new_n720), .ZN(new_n1249));
  AOI21_X1  g1049(.A(G390), .B1(new_n1249), .B2(new_n955), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n955), .B(G390), .C1(new_n981), .C2(new_n998), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n1242), .A2(new_n1244), .B1(new_n1250), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(G387), .A2(new_n1212), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1254), .A2(KEYINPUT126), .A3(new_n1251), .A4(new_n1243), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1253), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1218), .B1(new_n1221), .B2(new_n1223), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1258), .A2(KEYINPUT63), .A3(new_n1239), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1237), .A2(new_n1241), .A3(new_n1257), .A4(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT62), .ZN(new_n1261));
  AND3_X1   g1061(.A1(new_n1258), .A2(new_n1261), .A3(new_n1239), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT61), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1231), .A2(new_n1235), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1263), .B1(new_n1258), .B2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1261), .B1(new_n1258), .B2(new_n1239), .ZN(new_n1266));
  NOR3_X1   g1066(.A1(new_n1262), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1260), .B1(new_n1267), .B2(new_n1257), .ZN(G405));
  INV_X1    g1068(.A(new_n1221), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1180), .A2(new_n678), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT124), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1272), .A2(new_n1184), .A3(new_n1181), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1211), .B1(new_n1273), .B2(new_n1178), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1239), .B1(new_n1269), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(G375), .A2(new_n1216), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(new_n1240), .A3(new_n1221), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1275), .A2(new_n1256), .A3(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1256), .B1(new_n1275), .B2(new_n1277), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT127), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1278), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  AOI211_X1 g1081(.A(KEYINPUT127), .B(new_n1256), .C1(new_n1275), .C2(new_n1277), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(G402));
endmodule


