//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 0 0 1 0 1 1 0 1 1 1 0 0 0 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1277, new_n1278, new_n1279,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1361, new_n1362, new_n1363;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n202), .A2(G50), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT64), .Z(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n217));
  INV_X1    g0017(.A(G77), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  INV_X1    g0019(.A(G107), .ZN(new_n220));
  INV_X1    g0020(.A(G264), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n208), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n211), .B(new_n216), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  AND2_X1   g0044(.A1(KEYINPUT3), .A2(G33), .ZN(new_n245));
  NOR2_X1   g0045(.A1(KEYINPUT3), .A2(G33), .ZN(new_n246));
  NOR2_X1   g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n230), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G238), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G1698), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n247), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  AND2_X1   g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(new_n214), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT3), .B(G33), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n254), .B1(new_n255), .B2(G107), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G274), .ZN(new_n258));
  AND2_X1   g0058(.A1(G1), .A2(G13), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G41), .ZN(new_n262));
  INV_X1    g0062(.A(G45), .ZN(new_n263));
  AOI21_X1  g0063(.A(G1), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n259), .A2(new_n260), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n265), .B1(new_n219), .B2(new_n268), .ZN(new_n269));
  OR2_X1    g0069(.A1(new_n257), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G190), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n257), .A2(new_n269), .ZN(new_n273));
  INV_X1    g0073(.A(G200), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G20), .A2(G77), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT8), .B(G58), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n206), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n206), .A2(G33), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT15), .B(G87), .ZN(new_n281));
  OAI221_X1 g0081(.A(new_n276), .B1(new_n277), .B2(new_n279), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n214), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n282), .A2(new_n284), .B1(new_n218), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT67), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n288), .B1(new_n286), .B2(new_n284), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n205), .A2(G20), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n285), .A2(KEYINPUT67), .A3(new_n214), .A4(new_n283), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n289), .A2(G77), .A3(new_n290), .A4(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  NOR3_X1   g0093(.A1(new_n272), .A2(new_n275), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n255), .A2(G222), .A3(new_n248), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n255), .A2(G223), .A3(G1698), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n295), .B(new_n296), .C1(new_n218), .C2(new_n255), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n254), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n254), .A2(new_n264), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n299), .A2(G226), .B1(new_n264), .B2(new_n261), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G169), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G150), .ZN(new_n304));
  OAI22_X1  g0104(.A1(new_n277), .A2(new_n280), .B1(new_n304), .B2(new_n279), .ZN(new_n305));
  INV_X1    g0105(.A(G50), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n206), .B1(new_n201), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n284), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT65), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI211_X1 g0110(.A(KEYINPUT65), .B(new_n284), .C1(new_n305), .C2(new_n307), .ZN(new_n311));
  OAI21_X1  g0111(.A(G50), .B1(new_n206), .B2(G1), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n312), .B(KEYINPUT66), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n286), .A2(new_n284), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n313), .A2(new_n314), .B1(new_n306), .B2(new_n286), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n310), .A2(new_n311), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G179), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n298), .A2(new_n317), .A3(new_n300), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n303), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n299), .A2(G238), .ZN(new_n321));
  NAND2_X1  g0121(.A1(G33), .A2(G97), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT70), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT70), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n324), .A2(G33), .A3(G97), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(G226), .A2(G1698), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n327), .B1(new_n230), .B2(G1698), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n326), .B1(new_n255), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n321), .B1(new_n329), .B2(new_n266), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT71), .ZN(new_n331));
  OAI21_X1  g0131(.A(G274), .B1(new_n253), .B2(new_n214), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n331), .B1(new_n332), .B2(new_n267), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n261), .A2(KEYINPUT71), .A3(new_n264), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(KEYINPUT13), .B1(new_n330), .B2(new_n335), .ZN(new_n336));
  NOR3_X1   g0136(.A1(new_n254), .A2(new_n264), .A3(new_n250), .ZN(new_n337));
  INV_X1    g0137(.A(G226), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n248), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n230), .A2(G1698), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n339), .B(new_n340), .C1(new_n245), .C2(new_n246), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n341), .A2(new_n323), .A3(new_n325), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n337), .B1(new_n342), .B2(new_n254), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT13), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n333), .A2(new_n334), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n336), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G200), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT72), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(new_n279), .B2(new_n306), .ZN(new_n350));
  NOR2_X1   g0150(.A1(G20), .A2(G33), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n351), .A2(KEYINPUT72), .A3(G50), .ZN(new_n352));
  AND2_X1   g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  OAI22_X1  g0153(.A1(new_n280), .A2(new_n218), .B1(new_n206), .B2(G68), .ZN(new_n354));
  OAI211_X1 g0154(.A(KEYINPUT11), .B(new_n284), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT11), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n354), .B1(new_n350), .B2(new_n352), .ZN(new_n357));
  INV_X1    g0157(.A(new_n284), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n289), .A2(G68), .A3(new_n290), .A4(new_n291), .ZN(new_n360));
  INV_X1    g0160(.A(G68), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n286), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n362), .B(KEYINPUT12), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n355), .A2(new_n359), .A3(new_n360), .A4(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n342), .A2(new_n254), .ZN(new_n365));
  AND4_X1   g0165(.A1(new_n344), .A2(new_n365), .A3(new_n345), .A4(new_n321), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n344), .B1(new_n343), .B2(new_n345), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n364), .B1(new_n368), .B2(G190), .ZN(new_n369));
  AOI211_X1 g0169(.A(new_n294), .B(new_n320), .C1(new_n348), .C2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT16), .ZN(new_n371));
  OR2_X1    g0171(.A1(KEYINPUT3), .A2(G33), .ZN(new_n372));
  NAND2_X1  g0172(.A1(KEYINPUT3), .A2(G33), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n372), .A2(new_n206), .A3(new_n373), .ZN(new_n374));
  XNOR2_X1  g0174(.A(KEYINPUT74), .B(KEYINPUT7), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n372), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n373), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n361), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  AND2_X1   g0178(.A1(G58), .A2(G68), .ZN(new_n379));
  OAI21_X1  g0179(.A(G20), .B1(new_n379), .B2(new_n201), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT75), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n351), .A2(G159), .ZN(new_n383));
  OAI211_X1 g0183(.A(KEYINPUT75), .B(G20), .C1(new_n379), .C2(new_n201), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n371), .B1(new_n378), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n383), .ZN(new_n387));
  XNOR2_X1  g0187(.A(G58), .B(G68), .ZN(new_n388));
  AOI21_X1  g0188(.A(KEYINPUT75), .B1(new_n388), .B2(G20), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n247), .A2(new_n375), .A3(new_n206), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n374), .A2(KEYINPUT7), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n391), .A2(new_n392), .A3(G68), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n390), .A2(new_n393), .A3(KEYINPUT16), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n386), .A2(new_n394), .A3(new_n284), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n299), .A2(G232), .B1(new_n264), .B2(new_n261), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n338), .A2(G1698), .ZN(new_n397));
  OAI221_X1 g0197(.A(new_n397), .B1(G223), .B2(G1698), .C1(new_n245), .C2(new_n246), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G33), .A2(G87), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n396), .B(new_n271), .C1(new_n400), .C2(new_n266), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n266), .B1(new_n398), .B2(new_n399), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n265), .B1(new_n230), .B2(new_n268), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n274), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n277), .B1(new_n205), .B2(G20), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n406), .A2(new_n314), .B1(new_n277), .B2(new_n286), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n395), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT17), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n395), .A2(new_n405), .A3(KEYINPUT17), .A4(new_n407), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n395), .A2(new_n407), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n402), .A2(new_n403), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(G179), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n302), .B2(new_n414), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT18), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n413), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n417), .B1(new_n413), .B2(new_n416), .ZN(new_n420));
  NOR3_X1   g0220(.A1(new_n412), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  XNOR2_X1  g0221(.A(new_n364), .B(KEYINPUT73), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT14), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n423), .B(G169), .C1(new_n366), .C2(new_n367), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n336), .A2(G179), .A3(new_n346), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n423), .B1(new_n347), .B2(G169), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n422), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n270), .A2(new_n302), .B1(new_n287), .B2(new_n292), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n429), .A2(KEYINPUT68), .B1(new_n317), .B2(new_n273), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n293), .B1(G169), .B2(new_n273), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT68), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n370), .A2(new_n421), .A3(new_n428), .A4(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n301), .A2(G200), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n310), .A2(KEYINPUT9), .A3(new_n311), .A4(new_n315), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n298), .A2(G190), .A3(new_n300), .ZN(new_n438));
  AND3_X1   g0238(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT69), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT9), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n316), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n440), .B1(new_n316), .B2(new_n441), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n439), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT10), .ZN(new_n446));
  OR2_X1    g0246(.A1(new_n443), .A2(new_n444), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT10), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n447), .A2(new_n448), .A3(new_n439), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n435), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G116), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n451), .B1(new_n205), .B2(G33), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n289), .A2(new_n291), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT79), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT79), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n289), .A2(new_n455), .A3(new_n291), .A4(new_n452), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n205), .A2(new_n451), .A3(G13), .A4(G20), .ZN(new_n458));
  OR2_X1    g0258(.A1(new_n458), .A2(KEYINPUT80), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(KEYINPUT80), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n283), .A2(new_n214), .B1(G20), .B2(new_n451), .ZN(new_n462));
  NAND2_X1  g0262(.A1(G33), .A2(G283), .ZN(new_n463));
  INV_X1    g0263(.A(G97), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n463), .B(new_n206), .C1(G33), .C2(new_n464), .ZN(new_n465));
  AND3_X1   g0265(.A1(new_n462), .A2(KEYINPUT20), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(KEYINPUT20), .B1(new_n462), .B2(new_n465), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n457), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(G303), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n372), .A2(new_n471), .A3(new_n373), .ZN(new_n472));
  NOR2_X1   g0272(.A1(G257), .A2(G1698), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n473), .B1(new_n221), .B2(G1698), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n254), .B(new_n472), .C1(new_n474), .C2(new_n247), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n263), .A2(G1), .ZN(new_n476));
  XNOR2_X1  g0276(.A(KEYINPUT5), .B(G41), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n261), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  AND2_X1   g0278(.A1(KEYINPUT5), .A2(G41), .ZN(new_n479));
  NOR2_X1   g0279(.A1(KEYINPUT5), .A2(G41), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n476), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n481), .A2(G270), .A3(new_n266), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n475), .A2(new_n478), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G169), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n470), .A2(KEYINPUT21), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT21), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n468), .B1(new_n456), .B2(new_n454), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n487), .B1(new_n488), .B2(new_n484), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n475), .A2(G179), .A3(new_n482), .A4(new_n478), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n470), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n486), .A2(new_n489), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n483), .A2(G200), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n494), .B1(new_n271), .B2(new_n483), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(new_n470), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g0297(.A(G257), .B(G1698), .C1(new_n245), .C2(new_n246), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT83), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT83), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n255), .A2(new_n500), .A3(G257), .A4(G1698), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G33), .A2(G294), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n255), .A2(G250), .A3(new_n248), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n499), .A2(new_n501), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n254), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n254), .B1(new_n476), .B2(new_n477), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G264), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n505), .A2(new_n478), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n302), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT24), .ZN(new_n510));
  INV_X1    g0310(.A(G87), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n511), .A2(KEYINPUT81), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n512), .B(new_n206), .C1(new_n246), .C2(new_n245), .ZN(new_n513));
  XNOR2_X1  g0313(.A(KEYINPUT82), .B(KEYINPUT22), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n255), .A2(new_n514), .A3(new_n206), .A4(new_n512), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n220), .A2(KEYINPUT23), .A3(G20), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT23), .B1(new_n220), .B2(G20), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G33), .A2(G116), .ZN(new_n521));
  OAI22_X1  g0321(.A1(new_n519), .A2(new_n520), .B1(G20), .B2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n510), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  AOI211_X1 g0324(.A(KEYINPUT24), .B(new_n522), .C1(new_n516), .C2(new_n517), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n284), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n314), .B1(G1), .B2(new_n278), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT25), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n285), .B2(G107), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n286), .A2(KEYINPUT25), .A3(new_n220), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n528), .A2(G107), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n505), .A2(new_n478), .A3(new_n507), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n526), .A2(new_n532), .B1(new_n533), .B2(new_n317), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n508), .A2(new_n274), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(G190), .B2(new_n508), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n526), .A2(new_n532), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n509), .A2(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n281), .A2(new_n286), .ZN(new_n539));
  INV_X1    g0339(.A(new_n281), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n314), .B(new_n540), .C1(G1), .C2(new_n278), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n206), .B(G68), .C1(new_n245), .C2(new_n246), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT19), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n280), .B2(new_n464), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n324), .B1(G33), .B2(G97), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n322), .A2(KEYINPUT70), .ZN(new_n547));
  OAI21_X1  g0347(.A(KEYINPUT19), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n206), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n511), .A2(new_n464), .A3(new_n220), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n545), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n539), .B(new_n541), .C1(new_n551), .C2(new_n358), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n261), .A2(new_n476), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n205), .A2(G45), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n266), .A2(G250), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(G244), .B(G1698), .C1(new_n245), .C2(new_n246), .ZN(new_n558));
  OAI211_X1 g0358(.A(G238), .B(new_n248), .C1(new_n245), .C2(new_n246), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n558), .A2(new_n559), .A3(new_n521), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n254), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n302), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n556), .B1(new_n254), .B2(new_n560), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n317), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n552), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n562), .A2(G200), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n543), .B1(new_n323), .B2(new_n325), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n550), .B1(new_n568), .B2(G20), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n542), .A2(new_n544), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n571), .A2(new_n284), .B1(new_n286), .B2(new_n281), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n528), .A2(G87), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n557), .A2(new_n561), .A3(G190), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n567), .A2(new_n572), .A3(new_n573), .A4(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n279), .A2(new_n218), .ZN(new_n576));
  XNOR2_X1  g0376(.A(G97), .B(G107), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT6), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NOR3_X1   g0379(.A1(new_n578), .A2(new_n464), .A3(G107), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n576), .B1(new_n582), .B2(G20), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n376), .A2(new_n377), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(G107), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n358), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n285), .A2(G97), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT76), .ZN(new_n588));
  XNOR2_X1  g0388(.A(new_n587), .B(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(new_n527), .B2(new_n464), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n481), .A2(G257), .A3(new_n266), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n478), .ZN(new_n592));
  OAI211_X1 g0392(.A(G244), .B(new_n248), .C1(new_n245), .C2(new_n246), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT4), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n255), .A2(KEYINPUT4), .A3(G244), .A4(new_n248), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n255), .A2(G250), .A3(G1698), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n595), .A2(new_n596), .A3(new_n463), .A4(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n592), .B1(new_n598), .B2(new_n254), .ZN(new_n599));
  OAI22_X1  g0399(.A1(new_n586), .A2(new_n590), .B1(new_n599), .B2(G169), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n317), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n566), .B(new_n575), .C1(new_n600), .C2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n599), .A2(G190), .ZN(new_n604));
  XNOR2_X1  g0404(.A(new_n604), .B(KEYINPUT78), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n580), .B1(new_n578), .B2(new_n577), .ZN(new_n606));
  OAI22_X1  g0406(.A1(new_n606), .A2(new_n206), .B1(new_n218), .B2(new_n279), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n220), .B1(new_n376), .B2(new_n377), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n284), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n528), .A2(G97), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n609), .A2(new_n610), .A3(new_n589), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n598), .A2(new_n254), .ZN(new_n612));
  INV_X1    g0412(.A(new_n592), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(KEYINPUT77), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT77), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n274), .B1(new_n599), .B2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n611), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n603), .B1(new_n605), .B2(new_n618), .ZN(new_n619));
  AND4_X1   g0419(.A1(new_n450), .A2(new_n497), .A3(new_n538), .A4(new_n619), .ZN(G372));
  NAND2_X1  g0420(.A1(new_n413), .A2(new_n416), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(KEYINPUT18), .ZN(new_n622));
  INV_X1    g0422(.A(new_n428), .ZN(new_n623));
  INV_X1    g0423(.A(new_n434), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n369), .A2(new_n348), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n622), .B(new_n418), .C1(new_n626), .C2(new_n412), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n449), .A2(new_n446), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n320), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n526), .A2(new_n532), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n504), .A2(new_n254), .B1(G264), .B2(new_n506), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n631), .A2(new_n317), .A3(new_n478), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n630), .A2(new_n509), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT84), .B1(new_n633), .B2(new_n493), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n508), .A2(G190), .ZN(new_n635));
  AOI21_X1  g0435(.A(G200), .B1(new_n631), .B2(new_n478), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n526), .B(new_n532), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n486), .A2(new_n492), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n630), .A2(new_n509), .A3(new_n632), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT84), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n638), .A2(new_n639), .A3(new_n640), .A4(new_n489), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n634), .A2(new_n619), .A3(new_n637), .A4(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n566), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n566), .A2(new_n575), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n600), .A2(new_n602), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(KEYINPUT26), .A3(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT26), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n611), .B(new_n601), .C1(G169), .C2(new_n599), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n648), .B1(new_n644), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n643), .B1(new_n647), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n642), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n450), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n629), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g0454(.A(new_n654), .B(KEYINPUT85), .Z(G369));
  NAND3_X1  g0455(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(new_n658), .A3(G213), .ZN(new_n659));
  INV_X1    g0459(.A(G343), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n488), .A2(new_n662), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n493), .A2(new_n496), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT86), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n497), .A2(KEYINPUT86), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n486), .A2(new_n489), .A3(new_n492), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n666), .A2(new_n667), .B1(new_n668), .B2(new_n663), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n637), .B(new_n639), .C1(new_n537), .C2(new_n662), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n633), .A2(new_n661), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n669), .A2(G330), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT87), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n669), .A2(KEYINPUT87), .A3(G330), .A4(new_n672), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n493), .A2(new_n637), .A3(new_n639), .A4(new_n662), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n633), .A2(new_n662), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT88), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n677), .A2(new_n682), .ZN(G399));
  INV_X1    g0483(.A(new_n209), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(G41), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n550), .A2(G116), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(G1), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n212), .B2(new_n686), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT28), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT90), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n633), .B2(new_n493), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n668), .A2(KEYINPUT90), .A3(new_n639), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n692), .A2(new_n619), .A3(new_n693), .A4(new_n637), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(new_n651), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n695), .A2(KEYINPUT29), .A3(new_n662), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n661), .B1(new_n642), .B2(new_n651), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n696), .B1(KEYINPUT29), .B2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(G330), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n631), .A2(new_n599), .A3(new_n491), .A4(new_n564), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT30), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n483), .A2(new_n317), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n508), .A2(new_n614), .A3(new_n562), .A4(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n562), .A2(new_n490), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n705), .A2(KEYINPUT30), .A3(new_n631), .A4(new_n599), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n702), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  AND3_X1   g0507(.A1(new_n707), .A2(KEYINPUT31), .A3(new_n661), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT89), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n702), .A2(new_n704), .A3(KEYINPUT89), .A4(new_n706), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n710), .A2(new_n661), .A3(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT31), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n708), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n619), .A2(new_n497), .A3(new_n538), .A4(new_n662), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n699), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n698), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n690), .B1(new_n719), .B2(G1), .ZN(G364));
  INV_X1    g0520(.A(G13), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(G20), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n205), .B1(new_n722), .B2(G45), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n685), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n725), .B1(new_n669), .B2(G330), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n669), .A2(G330), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(G13), .A2(G33), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(G20), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n669), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n209), .A2(new_n255), .ZN(new_n734));
  INV_X1    g0534(.A(G355), .ZN(new_n735));
  OAI22_X1  g0535(.A1(new_n734), .A2(new_n735), .B1(G116), .B2(new_n209), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n684), .A2(new_n255), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n738), .B1(new_n213), .B2(new_n263), .ZN(new_n739));
  OR2_X1    g0539(.A1(new_n240), .A2(new_n263), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n736), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n214), .B1(G20), .B2(new_n302), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n731), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n725), .B1(new_n741), .B2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n742), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n206), .A2(G179), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G190), .A2(G200), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n750), .A2(KEYINPUT92), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(KEYINPUT92), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G329), .ZN(new_n755));
  INV_X1    g0555(.A(G283), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n747), .A2(new_n271), .A3(G200), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n747), .A2(G190), .A3(G200), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n756), .A2(new_n757), .B1(new_n758), .B2(new_n471), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n206), .A2(new_n317), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G200), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G190), .ZN(new_n762));
  XNOR2_X1  g0562(.A(KEYINPUT33), .B(G317), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n759), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n760), .A2(new_n748), .ZN(new_n765));
  INV_X1    g0565(.A(G311), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n247), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n760), .A2(G190), .A3(new_n274), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n767), .B1(G322), .B2(new_n769), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n271), .A2(G179), .A3(G200), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n206), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n761), .A2(new_n271), .ZN(new_n774));
  AOI22_X1  g0574(.A1(G294), .A2(new_n773), .B1(new_n774), .B2(G326), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n755), .A2(new_n764), .A3(new_n770), .A4(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n774), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n777), .A2(new_n306), .B1(new_n757), .B2(new_n220), .ZN(new_n778));
  INV_X1    g0578(.A(new_n762), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n779), .A2(new_n361), .B1(new_n758), .B2(new_n511), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n772), .B(KEYINPUT91), .Z(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G97), .ZN(new_n783));
  INV_X1    g0583(.A(G159), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n749), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT32), .ZN(new_n786));
  INV_X1    g0586(.A(G58), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n255), .B1(new_n768), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n765), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n788), .B1(G77), .B2(new_n789), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n781), .A2(new_n783), .A3(new_n786), .A4(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n746), .B1(new_n776), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n745), .A2(new_n792), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n726), .A2(new_n728), .B1(new_n733), .B2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(G396));
  AOI21_X1  g0595(.A(new_n662), .B1(new_n287), .B2(new_n292), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n434), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n294), .B1(new_n430), .B2(new_n433), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n797), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n697), .B(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n725), .B1(new_n801), .B2(new_n717), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(new_n717), .B2(new_n801), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n742), .A2(new_n729), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n725), .B1(G77), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n757), .A2(new_n511), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n779), .A2(new_n756), .B1(new_n758), .B2(new_n220), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n807), .B(new_n808), .C1(G303), .C2(new_n774), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n754), .A2(G311), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n247), .B1(new_n765), .B2(new_n451), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(G294), .B2(new_n769), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n809), .A2(new_n783), .A3(new_n810), .A4(new_n812), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n762), .A2(G150), .B1(new_n774), .B2(G137), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT93), .ZN(new_n815));
  INV_X1    g0615(.A(G143), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n768), .A2(new_n816), .B1(new_n765), .B2(new_n784), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(KEYINPUT34), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n754), .A2(G132), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n757), .A2(new_n361), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(new_n247), .ZN(new_n822));
  INV_X1    g0622(.A(new_n758), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n773), .A2(G58), .B1(new_n823), .B2(G50), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n819), .A2(new_n820), .A3(new_n822), .A4(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n818), .A2(KEYINPUT34), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n813), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT94), .ZN(new_n828));
  OR2_X1    g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n746), .B1(new_n827), .B2(new_n828), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n806), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n730), .B2(new_n800), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n803), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(G384));
  NOR2_X1   g0634(.A1(new_n722), .A2(new_n205), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT95), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n428), .A2(new_n836), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n422), .B(KEYINPUT95), .C1(new_n426), .C2(new_n427), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n839), .A2(new_n661), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n394), .A2(new_n284), .ZN(new_n841));
  AOI21_X1  g0641(.A(KEYINPUT16), .B1(new_n390), .B2(new_n393), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n407), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n659), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n843), .A2(new_n416), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n845), .A2(new_n846), .A3(new_n408), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(KEYINPUT37), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n413), .A2(new_n844), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT37), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n621), .A2(new_n849), .A3(new_n850), .A4(new_n408), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n622), .A2(new_n418), .A3(new_n410), .A4(new_n411), .ZN(new_n853));
  INV_X1    g0653(.A(new_n845), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n853), .A2(KEYINPUT97), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT97), .B1(new_n853), .B2(new_n854), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n852), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT38), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n858), .B1(new_n848), .B2(new_n851), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n855), .B2(new_n856), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n859), .A2(KEYINPUT39), .A3(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT98), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n850), .B1(new_n849), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n621), .A2(new_n849), .A3(new_n408), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n864), .B(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n853), .A2(new_n413), .A3(new_n844), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT38), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT99), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n861), .A2(new_n869), .ZN(new_n870));
  OAI211_X1 g0670(.A(KEYINPUT99), .B(new_n860), .C1(new_n855), .C2(new_n856), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n868), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n840), .B(new_n862), .C1(new_n872), .C2(KEYINPUT39), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n434), .A2(new_n661), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(new_n697), .B2(new_n800), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n422), .A2(new_n661), .B1(new_n369), .B2(new_n348), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n837), .A2(new_n838), .A3(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n426), .A2(new_n427), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n625), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(new_n422), .A3(new_n661), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT96), .B1(new_n875), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT96), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n661), .B(new_n799), .C1(new_n642), .C2(new_n651), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n884), .B(new_n881), .C1(new_n885), .C2(new_n874), .ZN(new_n886));
  INV_X1    g0686(.A(new_n852), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT97), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n421), .B2(new_n845), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n853), .A2(KEYINPUT97), .A3(new_n854), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n887), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n861), .B1(new_n891), .B2(KEYINPUT38), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n883), .A2(new_n886), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n659), .B1(new_n419), .B2(new_n420), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n873), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n895), .B(KEYINPUT100), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n696), .B(new_n450), .C1(KEYINPUT29), .C2(new_n697), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n629), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n896), .B(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n868), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n889), .A2(new_n890), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT99), .B1(new_n901), .B2(new_n860), .ZN(new_n902));
  INV_X1    g0702(.A(new_n871), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n900), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n799), .B1(new_n877), .B2(new_n880), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n712), .A2(new_n713), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n710), .A2(KEYINPUT31), .A3(new_n661), .A4(new_n711), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n906), .A2(new_n715), .A3(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT101), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n905), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n910), .A2(KEYINPUT40), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n905), .A2(new_n908), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(KEYINPUT101), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n904), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n912), .B1(new_n859), .B2(new_n861), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n914), .B1(KEYINPUT40), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n450), .A2(new_n908), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(G330), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(new_n916), .B2(new_n917), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n835), .B1(new_n899), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n899), .B2(new_n921), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n582), .A2(KEYINPUT35), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n582), .A2(KEYINPUT35), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n924), .A2(G116), .A3(new_n215), .A4(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT36), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n212), .A2(new_n218), .A3(new_n379), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n361), .A2(G50), .ZN(new_n929));
  OAI211_X1 g0729(.A(G1), .B(new_n721), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n923), .A2(new_n927), .A3(new_n930), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n931), .B(KEYINPUT102), .Z(G367));
  OAI221_X1 g0732(.A(new_n743), .B1(new_n209), .B2(new_n281), .C1(new_n738), .C2(new_n236), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n933), .A2(new_n725), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n662), .B1(new_n572), .B2(new_n573), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n643), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n644), .B2(new_n935), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n768), .A2(new_n304), .B1(new_n765), .B2(new_n306), .ZN(new_n938));
  AOI211_X1 g0738(.A(new_n247), .B(new_n938), .C1(G137), .C2(new_n750), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n782), .A2(G68), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n762), .A2(G159), .B1(new_n774), .B2(G143), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n757), .A2(new_n218), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(G58), .B2(new_n823), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n939), .A2(new_n940), .A3(new_n941), .A4(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n757), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n762), .A2(G294), .B1(new_n945), .B2(G97), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n946), .B1(new_n220), .B2(new_n772), .C1(new_n766), .C2(new_n777), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n769), .A2(G303), .B1(new_n750), .B2(G317), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT46), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n758), .B2(new_n451), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n823), .A2(KEYINPUT46), .A3(G116), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n255), .B1(new_n789), .B2(G283), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n948), .A2(new_n950), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n944), .B1(new_n947), .B2(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT47), .Z(new_n955));
  OAI221_X1 g0755(.A(new_n934), .B1(new_n937), .B2(new_n732), .C1(new_n955), .C2(new_n746), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT103), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n646), .B1(new_n611), .B2(new_n661), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n618), .A2(new_n605), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n649), .A2(new_n662), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n957), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  AOI211_X1 g0763(.A(KEYINPUT103), .B(new_n961), .C1(new_n958), .C2(new_n959), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OR3_X1    g0765(.A1(new_n965), .A2(KEYINPUT104), .A3(new_n678), .ZN(new_n966));
  OAI21_X1  g0766(.A(KEYINPUT104), .B1(new_n965), .B2(new_n678), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(KEYINPUT42), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT42), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n966), .A2(new_n970), .A3(new_n967), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n649), .B1(new_n965), .B2(new_n639), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n662), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n969), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(KEYINPUT105), .B1(new_n677), .B2(new_n965), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT105), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n960), .A2(new_n962), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(KEYINPUT103), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n960), .A2(new_n957), .A3(new_n962), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n675), .A2(new_n980), .A3(new_n676), .A4(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n977), .A2(new_n979), .A3(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n979), .B1(new_n977), .B2(new_n985), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n976), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n977), .A2(new_n985), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n978), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n991), .A2(new_n975), .A3(new_n974), .A4(new_n986), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT44), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n682), .B2(new_n984), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n680), .B(KEYINPUT88), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n996), .A2(KEYINPUT44), .A3(new_n965), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT45), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n996), .B2(new_n965), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n682), .A2(new_n984), .A3(KEYINPUT45), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n998), .A2(new_n1002), .ZN(new_n1003));
  AND2_X1   g0803(.A1(new_n675), .A2(new_n676), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n664), .A2(new_n665), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n663), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1006), .A2(new_n667), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n668), .A2(new_n663), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1008), .A2(G330), .A3(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n668), .A2(new_n661), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n678), .B1(new_n672), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n669), .A2(G330), .A3(new_n1012), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1016), .A2(new_n698), .A3(KEYINPUT106), .A4(new_n717), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1016), .A2(new_n698), .A3(new_n717), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT106), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n677), .A2(new_n998), .A3(new_n1002), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1005), .A2(new_n1017), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(new_n719), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n685), .B(KEYINPUT41), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n724), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n956), .B1(new_n993), .B2(new_n1025), .ZN(G387));
  NAND3_X1  g0826(.A1(new_n670), .A2(new_n671), .A3(new_n731), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n734), .A2(new_n687), .B1(G107), .B2(new_n209), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n277), .A2(G50), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT108), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT107), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1031), .A2(KEYINPUT50), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(KEYINPUT50), .ZN(new_n1033));
  AOI21_X1  g0833(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1032), .A2(new_n687), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n738), .B1(new_n233), .B2(G45), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1028), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n725), .B1(new_n1037), .B2(new_n744), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n768), .A2(new_n306), .B1(new_n749), .B2(new_n304), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n247), .B(new_n1039), .C1(G68), .C2(new_n789), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n782), .A2(new_n540), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n277), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n762), .A2(new_n1042), .B1(new_n945), .B2(G97), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n774), .A2(G159), .B1(new_n823), .B2(G77), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1040), .A2(new_n1041), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n769), .A2(G317), .B1(new_n789), .B2(G303), .ZN(new_n1046));
  INV_X1    g0846(.A(G322), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1046), .B1(new_n779), .B2(new_n766), .C1(new_n1047), .C2(new_n777), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT48), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1051));
  INV_X1    g0851(.A(G294), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n772), .A2(new_n756), .B1(new_n758), .B2(new_n1052), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT109), .Z(new_n1054));
  NAND3_X1  g0854(.A1(new_n1050), .A2(new_n1051), .A3(new_n1054), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT49), .Z(new_n1056));
  AOI21_X1  g0856(.A(new_n255), .B1(new_n750), .B2(G326), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n451), .B2(new_n757), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT110), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1045), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1038), .B1(new_n1060), .B2(new_n742), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n1016), .A2(new_n724), .B1(new_n1027), .B2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n719), .A2(new_n1016), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n685), .B(KEYINPUT111), .Z(new_n1064));
  NAND2_X1  g0864(.A1(new_n1018), .A2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1062), .B1(new_n1063), .B2(new_n1065), .ZN(G393));
  INV_X1    g0866(.A(new_n725), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n737), .A2(new_n243), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n744), .B1(G97), .B2(new_n684), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n772), .A2(new_n451), .B1(new_n765), .B2(new_n1052), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(G317), .A2(new_n774), .B1(new_n769), .B2(G311), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT52), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1071), .B(new_n1073), .C1(G303), .C2(new_n762), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n247), .B1(new_n749), .B2(new_n1047), .C1(new_n220), .C2(new_n757), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(G283), .B2(new_n823), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT112), .Z(new_n1077));
  OAI22_X1  g0877(.A1(new_n361), .A2(new_n758), .B1(new_n757), .B2(new_n511), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n255), .B1(new_n749), .B2(new_n816), .C1(new_n277), .C2(new_n765), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1078), .B(new_n1079), .C1(G50), .C2(new_n762), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n777), .A2(new_n304), .B1(new_n784), .B2(new_n768), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT51), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n782), .A2(G77), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1085));
  AND3_X1   g0885(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1074), .A2(new_n1077), .B1(new_n1080), .B2(new_n1086), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n1070), .B1(new_n746), .B2(new_n1087), .C1(new_n984), .C2(new_n732), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1005), .A2(new_n1021), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1088), .B1(new_n1089), .B2(new_n723), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1021), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n677), .B1(new_n1002), .B2(new_n998), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1018), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1022), .B(new_n1064), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1096), .A2(KEYINPUT113), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT113), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1064), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(new_n1089), .B2(new_n1018), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1098), .B1(new_n1100), .B2(new_n1022), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1091), .B1(new_n1097), .B2(new_n1101), .ZN(G390));
  OAI21_X1  g0902(.A(new_n862), .B1(new_n872), .B2(KEYINPUT39), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n875), .A2(new_n882), .B1(new_n661), .B2(new_n839), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n872), .A2(new_n840), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n661), .B1(new_n694), .B2(new_n651), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n874), .B1(new_n1107), .B2(new_n800), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1108), .A2(new_n882), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1106), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n716), .A2(new_n800), .A3(new_n881), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n1105), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n905), .A2(new_n908), .A3(G330), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(new_n1105), .B2(new_n1111), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT114), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n697), .A2(new_n800), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n874), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n881), .B1(new_n716), .B2(new_n800), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1121), .B1(new_n1122), .B2(new_n1114), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n908), .A2(G330), .A3(new_n800), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n882), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1125), .A2(new_n1108), .A3(new_n1112), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n450), .A2(G330), .A3(new_n908), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n897), .A2(new_n629), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1118), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1131));
  AND3_X1   g0931(.A1(new_n897), .A2(new_n629), .A3(new_n1128), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1131), .A2(new_n1132), .A3(KEYINPUT114), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1099), .B1(new_n1117), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1105), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1103), .A2(new_n1104), .B1(new_n1106), .B2(new_n1110), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1136), .B1(new_n1137), .B2(new_n1115), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n1131), .A2(new_n1132), .A3(KEYINPUT114), .ZN(new_n1139));
  AOI21_X1  g0939(.A(KEYINPUT114), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n1138), .A2(new_n1141), .A3(KEYINPUT115), .ZN(new_n1142));
  AOI21_X1  g0942(.A(KEYINPUT115), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1135), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1117), .A2(new_n724), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n725), .B1(new_n1042), .B2(new_n805), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n220), .A2(new_n779), .B1(new_n777), .B2(new_n756), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n821), .B(new_n1147), .C1(G87), .C2(new_n823), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n754), .A2(G294), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n247), .B1(new_n768), .B2(new_n451), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(G97), .B2(new_n789), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1148), .A2(new_n1084), .A3(new_n1149), .A4(new_n1151), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n758), .A2(new_n304), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT53), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(KEYINPUT54), .B(G143), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n255), .B1(new_n765), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(G132), .B2(new_n769), .ZN(new_n1157));
  INV_X1    g0957(.A(G125), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1154), .B(new_n1157), .C1(new_n1158), .C2(new_n753), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n762), .A2(G137), .B1(new_n945), .B2(G50), .ZN(new_n1160));
  INV_X1    g0960(.A(G128), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n782), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1160), .B1(new_n1161), .B2(new_n777), .C1(new_n1162), .C2(new_n784), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1152), .B1(new_n1159), .B2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1146), .B1(new_n1164), .B2(new_n742), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1103), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1165), .B1(new_n1166), .B2(new_n730), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1145), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1144), .A2(new_n1169), .ZN(G378));
  OAI21_X1  g0970(.A(new_n725), .B1(G50), .B2(new_n805), .ZN(new_n1171));
  XOR2_X1   g0971(.A(new_n1171), .B(KEYINPUT118), .Z(new_n1172));
  NOR2_X1   g0972(.A1(new_n255), .A2(G41), .ZN(new_n1173));
  AOI211_X1 g0973(.A(G50), .B(new_n1173), .C1(new_n278), .C2(new_n262), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n1173), .B1(new_n765), .B2(new_n281), .C1(new_n220), .C2(new_n768), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n754), .B2(G283), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n762), .A2(G97), .B1(new_n823), .B2(G77), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n757), .A2(new_n787), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G116), .B2(new_n774), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1176), .A2(new_n940), .A3(new_n1177), .A4(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT58), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1174), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(G137), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n768), .A2(new_n1161), .B1(new_n765), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(G132), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n779), .A2(new_n1185), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1184), .B(new_n1186), .C1(G125), .C2(new_n774), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n758), .A2(new_n1155), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT116), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1187), .B(new_n1189), .C1(new_n304), .C2(new_n1162), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n945), .A2(G159), .ZN(new_n1192));
  AOI211_X1 g0992(.A(G33), .B(G41), .C1(new_n750), .C2(G124), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1182), .B1(new_n1181), .B2(new_n1180), .C1(new_n1194), .C2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(new_n742), .ZN(new_n1197));
  XOR2_X1   g0997(.A(new_n1197), .B(KEYINPUT117), .Z(new_n1198));
  XOR2_X1   g0998(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n316), .A2(new_n844), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n628), .B2(new_n319), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1201), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n320), .B(new_n1203), .C1(new_n449), .C2(new_n446), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(new_n1202), .A2(new_n1204), .A3(KEYINPUT119), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT119), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n448), .B1(new_n447), .B2(new_n439), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n445), .A2(KEYINPUT10), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n319), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n1203), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n628), .A2(new_n319), .A3(new_n1201), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1206), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1200), .B1(new_n1205), .B2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(KEYINPUT119), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1210), .A2(new_n1211), .A3(new_n1206), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1214), .A2(new_n1215), .A3(new_n1199), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1213), .A2(new_n1216), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1172), .B(new_n1198), .C1(new_n1217), .C2(new_n729), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n873), .A2(new_n893), .A3(new_n894), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n912), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n892), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT40), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n699), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1213), .A2(new_n1216), .ZN(new_n1224));
  AND3_X1   g1024(.A1(new_n1223), .A2(new_n914), .A3(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1224), .B1(new_n1223), .B2(new_n914), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1219), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1223), .A2(new_n914), .A3(new_n1224), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n913), .A2(KEYINPUT40), .A3(new_n910), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1229), .A2(new_n872), .ZN(new_n1230));
  OAI21_X1  g1030(.A(G330), .B1(new_n915), .B2(KEYINPUT40), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1217), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n895), .A2(new_n1228), .A3(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1227), .A2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1218), .B1(new_n1234), .B2(new_n724), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1129), .B(KEYINPUT120), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT57), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(new_n1227), .B2(new_n1233), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n1064), .ZN(new_n1241));
  AOI21_X1  g1041(.A(KEYINPUT57), .B1(new_n1237), .B2(new_n1234), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1235), .B1(new_n1241), .B2(new_n1242), .ZN(G375));
  NOR2_X1   g1043(.A1(new_n881), .A2(new_n730), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n1244), .B(KEYINPUT121), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1067), .B1(new_n361), .B2(new_n804), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n777), .A2(new_n1052), .B1(new_n758), .B2(new_n464), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n942), .B(new_n1247), .C1(G116), .C2(new_n762), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n754), .A2(G303), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n247), .B1(new_n765), .B2(new_n220), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(G283), .B2(new_n769), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1248), .A2(new_n1041), .A3(new_n1249), .A4(new_n1251), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n777), .A2(new_n1185), .B1(new_n758), .B2(new_n784), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n779), .A2(new_n1155), .ZN(new_n1254));
  NOR3_X1   g1054(.A1(new_n1253), .A2(new_n1254), .A3(new_n1178), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n754), .A2(G128), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n782), .A2(G50), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n255), .B1(new_n768), .B2(new_n1183), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(G150), .B2(new_n789), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1255), .A2(new_n1256), .A3(new_n1257), .A4(new_n1259), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1252), .A2(new_n1260), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1245), .B(new_n1246), .C1(new_n746), .C2(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(new_n1127), .B2(new_n723), .ZN(new_n1263));
  XOR2_X1   g1063(.A(new_n1263), .B(KEYINPUT122), .Z(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1141), .A2(new_n1024), .A3(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1265), .A2(new_n1267), .ZN(G381));
  OR3_X1    g1068(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1269));
  NOR4_X1   g1069(.A1(G381), .A2(G390), .A3(G387), .A4(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1143), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1138), .A2(new_n1141), .A3(KEYINPUT115), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1168), .B1(new_n1273), .B2(new_n1135), .ZN(new_n1274));
  INV_X1    g1074(.A(G375), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1270), .A2(new_n1274), .A3(new_n1275), .ZN(G407));
  NAND2_X1  g1076(.A1(new_n660), .A2(G213), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1275), .A2(new_n1274), .A3(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(G407), .A2(G213), .A3(new_n1279), .ZN(G409));
  XNOR2_X1  g1080(.A(G393), .B(new_n794), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n992), .B(new_n989), .C1(new_n1282), .C2(new_n724), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(G390), .A2(new_n1283), .A3(new_n956), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1096), .A2(KEYINPUT113), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1100), .A2(new_n1098), .A3(new_n1022), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1090), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(G387), .A2(new_n1287), .A3(KEYINPUT125), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1284), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT125), .B1(G387), .B2(new_n1287), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1281), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(G387), .A2(new_n1287), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(KEYINPUT126), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1281), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT126), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(G387), .A2(new_n1287), .A3(new_n1295), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1293), .A2(new_n1294), .A3(new_n1284), .A4(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1291), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT62), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1237), .A2(new_n1024), .A3(new_n1234), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1235), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1301), .A2(new_n1144), .A3(new_n1169), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1302), .B1(G375), .B2(new_n1274), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1127), .A2(KEYINPUT60), .A3(new_n1129), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1064), .ZN(new_n1305));
  XOR2_X1   g1105(.A(KEYINPUT123), .B(KEYINPUT60), .Z(new_n1306));
  NAND3_X1  g1106(.A1(new_n1130), .A2(new_n1133), .A3(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(new_n1266), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1305), .B1(new_n1308), .B2(KEYINPUT124), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT124), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1307), .A2(new_n1310), .A3(new_n1266), .ZN(new_n1311));
  AOI211_X1 g1111(.A(new_n833), .B(new_n1264), .C1(new_n1309), .C2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1308), .A2(KEYINPUT124), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1305), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1313), .A2(new_n1311), .A3(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(G384), .B1(new_n1315), .B2(new_n1265), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1312), .A2(new_n1316), .ZN(new_n1317));
  AND4_X1   g1117(.A1(new_n1299), .A2(new_n1303), .A3(new_n1277), .A4(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n840), .B1(new_n1121), .B2(new_n881), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT39), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n904), .A2(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1319), .B1(new_n1321), .B2(new_n862), .ZN(new_n1322));
  NOR3_X1   g1122(.A1(new_n1109), .A2(new_n872), .A3(new_n840), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1114), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1324));
  OAI211_X1 g1124(.A(new_n1324), .B(new_n1136), .C1(new_n1140), .C2(new_n1139), .ZN(new_n1325));
  AOI22_X1  g1125(.A1(new_n1325), .A2(new_n1236), .B1(new_n1233), .B2(new_n1227), .ZN(new_n1326));
  OAI211_X1 g1126(.A(new_n1240), .B(new_n1064), .C1(new_n1326), .C2(KEYINPUT57), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(G378), .A2(new_n1327), .A3(new_n1235), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1278), .B1(new_n1328), .B2(new_n1302), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1299), .B1(new_n1329), .B2(new_n1317), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1318), .A2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1278), .A2(G2897), .ZN(new_n1332));
  AOI22_X1  g1132(.A1(new_n1303), .A2(new_n1277), .B1(new_n1317), .B2(new_n1332), .ZN(new_n1333));
  OAI211_X1 g1133(.A(G2897), .B(new_n1278), .C1(new_n1312), .C2(new_n1316), .ZN(new_n1334));
  AOI21_X1  g1134(.A(KEYINPUT61), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1298), .B1(new_n1331), .B2(new_n1335), .ZN(new_n1336));
  AOI21_X1  g1136(.A(KEYINPUT61), .B1(new_n1291), .B2(new_n1297), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1329), .A2(KEYINPUT63), .A3(new_n1317), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1303), .A2(new_n1277), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1317), .A2(new_n1332), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1340), .A2(new_n1334), .A3(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(KEYINPUT63), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1303), .A2(new_n1277), .A3(new_n1317), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1339), .B1(new_n1343), .B2(new_n1344), .ZN(new_n1345));
  OAI21_X1  g1145(.A(KEYINPUT127), .B1(new_n1336), .B2(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1344), .A2(KEYINPUT62), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT61), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1329), .A2(new_n1299), .A3(new_n1317), .ZN(new_n1349));
  NAND4_X1  g1149(.A1(new_n1342), .A2(new_n1347), .A3(new_n1348), .A4(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1298), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1352));
  AND2_X1   g1152(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT63), .ZN(new_n1354));
  AOI21_X1  g1154(.A(new_n1354), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1355));
  INV_X1    g1155(.A(new_n1344), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1353), .B1(new_n1355), .B2(new_n1356), .ZN(new_n1357));
  INV_X1    g1157(.A(KEYINPUT127), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1352), .A2(new_n1357), .A3(new_n1358), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1346), .A2(new_n1359), .ZN(G405));
  NAND2_X1  g1160(.A1(G375), .A2(new_n1274), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1361), .A2(new_n1328), .ZN(new_n1362));
  XNOR2_X1  g1162(.A(new_n1298), .B(new_n1362), .ZN(new_n1363));
  XOR2_X1   g1163(.A(new_n1363), .B(new_n1317), .Z(G402));
endmodule


