//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 0 0 0 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1 0 0 1 0 0 0 1 0 0 0 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1247, new_n1248, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  INV_X1    g0003(.A(G68), .ZN(new_n204));
  INV_X1    g0004(.A(G238), .ZN(new_n205));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G257), .ZN(new_n207));
  OAI22_X1  g0007(.A1(new_n204), .A2(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT65), .ZN(new_n210));
  AOI211_X1 g0010(.A(new_n208), .B(new_n210), .C1(G77), .C2(G244), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G87), .A2(G250), .ZN(new_n212));
  INV_X1    g0012(.A(G58), .ZN(new_n213));
  INV_X1    g0013(.A(G232), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n211), .B(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AND2_X1   g0015(.A1(G107), .A2(G264), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n203), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT1), .ZN(new_n218));
  NOR2_X1   g0018(.A1(G58), .A2(G68), .ZN(new_n219));
  OR2_X1    g0019(.A1(new_n219), .A2(KEYINPUT64), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(KEYINPUT64), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n220), .A2(G50), .A3(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  NOR3_X1   g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n203), .A2(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT0), .Z(new_n228));
  NOR3_X1   g0028(.A1(new_n218), .A2(new_n225), .A3(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G264), .ZN(new_n235));
  INV_X1    g0035(.A(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n233), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(KEYINPUT3), .ZN(new_n246));
  INV_X1    g0046(.A(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G1698), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G222), .ZN(new_n252));
  INV_X1    g0052(.A(G223), .ZN(new_n253));
  OAI211_X1 g0053(.A(new_n250), .B(new_n252), .C1(new_n253), .C2(new_n251), .ZN(new_n254));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  OAI211_X1 g0055(.A(G1), .B(G13), .C1(new_n247), .C2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  OAI211_X1 g0057(.A(new_n254), .B(new_n257), .C1(G77), .C2(new_n250), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n259), .B1(G41), .B2(G45), .ZN(new_n260));
  INV_X1    g0060(.A(G274), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n256), .A2(new_n260), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G226), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n258), .A2(new_n263), .A3(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G190), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n223), .A2(G33), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n270), .B(KEYINPUT67), .ZN(new_n271));
  NOR2_X1   g0071(.A1(KEYINPUT8), .A2(G58), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT66), .B(G58), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n272), .B1(new_n273), .B2(KEYINPUT8), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G50), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n223), .B1(new_n219), .B2(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G20), .A2(G33), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n277), .B1(G150), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n224), .ZN(new_n282));
  INV_X1    g0082(.A(G13), .ZN(new_n283));
  NOR3_X1   g0083(.A1(new_n283), .A2(new_n223), .A3(G1), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n280), .A2(new_n282), .B1(new_n276), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n282), .B1(new_n259), .B2(G20), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n285), .B1(new_n276), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT71), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n288), .A2(new_n289), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n269), .B1(new_n293), .B2(KEYINPUT9), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT10), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT9), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n291), .A2(new_n296), .A3(new_n292), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n267), .A2(G200), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n294), .A2(new_n295), .A3(new_n297), .A4(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n292), .ZN(new_n300));
  OAI21_X1  g0100(.A(KEYINPUT9), .B1(new_n300), .B2(new_n290), .ZN(new_n301));
  INV_X1    g0101(.A(new_n269), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n301), .A2(new_n297), .A3(new_n298), .A4(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT10), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n299), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n284), .A2(new_n204), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n306), .A2(KEYINPUT12), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(KEYINPUT12), .ZN(new_n308));
  OAI22_X1  g0108(.A1(new_n307), .A2(new_n308), .B1(new_n287), .B2(new_n204), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n271), .A2(G77), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n278), .A2(G50), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n204), .A2(G20), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n282), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT11), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT11), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n313), .A2(new_n316), .A3(new_n282), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n309), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT13), .ZN(new_n319));
  AND2_X1   g0119(.A1(KEYINPUT3), .A2(G33), .ZN(new_n320));
  NOR2_X1   g0120(.A1(KEYINPUT3), .A2(G33), .ZN(new_n321));
  OAI211_X1 g0121(.A(G226), .B(new_n251), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  OAI211_X1 g0122(.A(G232), .B(G1698), .C1(new_n320), .C2(new_n321), .ZN(new_n323));
  NAND2_X1  g0123(.A1(G33), .A2(G97), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n257), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n265), .A2(G238), .ZN(new_n327));
  AND4_X1   g0127(.A1(new_n319), .A2(new_n326), .A3(new_n327), .A4(new_n263), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n262), .B1(new_n325), .B2(new_n257), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n319), .B1(new_n329), .B2(new_n327), .ZN(new_n330));
  OAI21_X1  g0130(.A(G200), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n330), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n329), .A2(new_n319), .A3(new_n327), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n332), .A2(G190), .A3(new_n333), .ZN(new_n334));
  AND3_X1   g0134(.A1(new_n318), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n328), .A2(new_n330), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT14), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n336), .A2(G179), .B1(KEYINPUT72), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(G169), .B1(new_n328), .B2(new_n330), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n337), .A2(KEYINPUT72), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI221_X1 g0141(.A(G169), .B1(KEYINPUT72), .B2(new_n337), .C1(new_n328), .C2(new_n330), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n338), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n318), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n335), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n267), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n288), .B1(G169), .B2(new_n346), .ZN(new_n347));
  XOR2_X1   g0147(.A(new_n347), .B(KEYINPUT68), .Z(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(G179), .B2(new_n267), .ZN(new_n349));
  XNOR2_X1  g0149(.A(KEYINPUT8), .B(G58), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n351), .A2(new_n278), .B1(G20), .B2(G77), .ZN(new_n352));
  XOR2_X1   g0152(.A(KEYINPUT15), .B(G87), .Z(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n352), .B1(new_n270), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G77), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n355), .A2(new_n282), .B1(new_n356), .B2(new_n284), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n286), .A2(G77), .ZN(new_n358));
  AND3_X1   g0158(.A1(new_n357), .A2(KEYINPUT70), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(KEYINPUT70), .B1(new_n357), .B2(new_n358), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n320), .A2(new_n321), .ZN(new_n362));
  OAI21_X1  g0162(.A(KEYINPUT69), .B1(new_n362), .B2(new_n205), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(G1698), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n250), .A2(KEYINPUT69), .A3(G232), .A4(new_n251), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n362), .A2(G107), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT69), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n362), .B2(new_n214), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n364), .A2(new_n365), .A3(new_n366), .A4(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n262), .B1(new_n369), .B2(new_n257), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n265), .A2(G244), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n361), .B1(new_n268), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n372), .ZN(new_n374));
  INV_X1    g0174(.A(G200), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OR2_X1    g0176(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n305), .A2(new_n345), .A3(new_n349), .A4(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT18), .ZN(new_n379));
  INV_X1    g0179(.A(new_n284), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n274), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n381), .B1(new_n286), .B2(new_n274), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n248), .A2(new_n223), .A3(new_n249), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT7), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT73), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n248), .A2(KEYINPUT7), .A3(new_n223), .A4(new_n249), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n388), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT73), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n389), .A2(G68), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n278), .ZN(new_n393));
  INV_X1    g0193(.A(G159), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n213), .A2(KEYINPUT66), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT66), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(G58), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n396), .A2(new_n398), .A3(G68), .ZN(new_n399));
  INV_X1    g0199(.A(new_n219), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n395), .B1(new_n401), .B2(G20), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n392), .A2(KEYINPUT16), .A3(new_n402), .ZN(new_n403));
  AND2_X1   g0203(.A1(new_n403), .A2(new_n282), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT16), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n219), .B1(new_n273), .B2(G68), .ZN(new_n406));
  OAI22_X1  g0206(.A1(new_n406), .A2(new_n223), .B1(new_n394), .B2(new_n393), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n204), .B1(new_n386), .B2(new_n388), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n405), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT74), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(KEYINPUT7), .B1(new_n362), .B2(new_n223), .ZN(new_n412));
  OAI21_X1  g0212(.A(G68), .B1(new_n412), .B2(new_n390), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n402), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n414), .A2(KEYINPUT74), .A3(new_n405), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n383), .B1(new_n404), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n262), .B1(new_n265), .B2(G232), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n253), .A2(new_n251), .ZN(new_n419));
  OAI221_X1 g0219(.A(new_n419), .B1(G226), .B2(new_n251), .C1(new_n320), .C2(new_n321), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G33), .A2(G87), .ZN(new_n421));
  AND2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n418), .B(G179), .C1(new_n256), .C2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n256), .B1(new_n420), .B2(new_n421), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n263), .B1(new_n264), .B2(new_n214), .ZN(new_n425));
  OAI21_X1  g0225(.A(G169), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n379), .B1(new_n417), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n403), .A2(new_n282), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n430), .B1(new_n411), .B2(new_n415), .ZN(new_n431));
  OAI211_X1 g0231(.A(KEYINPUT18), .B(new_n427), .C1(new_n431), .C2(new_n383), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT75), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT17), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n418), .B(G190), .C1(new_n422), .C2(new_n256), .ZN(new_n436));
  OAI21_X1  g0236(.A(G200), .B1(new_n424), .B2(new_n425), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(new_n382), .A3(new_n437), .ZN(new_n438));
  AOI211_X1 g0238(.A(new_n435), .B(new_n438), .C1(new_n404), .C2(new_n416), .ZN(new_n439));
  AOI21_X1  g0239(.A(KEYINPUT74), .B1(new_n414), .B2(new_n405), .ZN(new_n440));
  AOI211_X1 g0240(.A(new_n410), .B(KEYINPUT16), .C1(new_n413), .C2(new_n402), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n282), .B(new_n403), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n438), .ZN(new_n443));
  AOI21_X1  g0243(.A(KEYINPUT17), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n434), .B1(new_n439), .B2(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n440), .A2(new_n441), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n443), .B1(new_n446), .B2(new_n430), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n435), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n442), .A2(KEYINPUT17), .A3(new_n443), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n448), .A2(KEYINPUT75), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n433), .A2(new_n445), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n361), .ZN(new_n452));
  INV_X1    g0252(.A(G169), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n372), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(G179), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n374), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n452), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  OR2_X1    g0258(.A1(new_n451), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n378), .A2(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(G264), .B(G1698), .C1(new_n320), .C2(new_n321), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT80), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT80), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n250), .A2(new_n463), .A3(G264), .A4(G1698), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n362), .A2(G303), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n250), .A2(G257), .A3(new_n251), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n462), .A2(new_n464), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n257), .ZN(new_n468));
  INV_X1    g0268(.A(G45), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(G1), .ZN(new_n470));
  AND2_X1   g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  NOR2_X1   g0271(.A1(KEYINPUT5), .A2(G41), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n256), .ZN(new_n474));
  OAI21_X1  g0274(.A(KEYINPUT79), .B1(new_n474), .B2(new_n236), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT79), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n473), .A2(new_n476), .A3(G270), .A4(new_n256), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  OR2_X1    g0278(.A1(new_n473), .A2(new_n261), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n468), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n247), .A2(G1), .ZN(new_n481));
  NOR3_X1   g0281(.A1(new_n284), .A2(new_n282), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G116), .ZN(new_n483));
  INV_X1    g0283(.A(G116), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n284), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G283), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n486), .B(new_n223), .C1(G33), .C2(new_n206), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n487), .B(new_n282), .C1(new_n223), .C2(G116), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT20), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n488), .A2(new_n489), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n483), .B(new_n485), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n480), .A2(new_n492), .A3(G169), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT81), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(KEYINPUT21), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT21), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n493), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n480), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n499), .A2(G179), .A3(new_n492), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n480), .A2(G200), .ZN(new_n501));
  INV_X1    g0301(.A(new_n492), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n501), .B(new_n502), .C1(new_n268), .C2(new_n480), .ZN(new_n503));
  AND4_X1   g0303(.A1(new_n496), .A2(new_n498), .A3(new_n500), .A4(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n470), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n256), .A2(new_n505), .A3(G250), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n250), .A2(G244), .A3(G1698), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n250), .A2(G238), .A3(new_n251), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G33), .A2(G116), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n507), .B1(new_n511), .B2(new_n257), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n470), .A2(G274), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT76), .ZN(new_n514));
  XNOR2_X1  g0314(.A(new_n513), .B(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n512), .A2(G190), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT78), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT78), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n512), .A2(new_n518), .A3(G190), .A4(new_n515), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(G97), .A2(G107), .ZN(new_n521));
  INV_X1    g0321(.A(G87), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n324), .A2(new_n223), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(KEYINPUT19), .A3(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n223), .B(G68), .C1(new_n320), .C2(new_n321), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n324), .A2(G20), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n525), .B(new_n526), .C1(KEYINPUT19), .C2(new_n527), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n528), .A2(new_n282), .B1(new_n284), .B2(new_n354), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n482), .A2(G87), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n511), .A2(new_n257), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n532), .A2(new_n506), .A3(new_n515), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n531), .B1(G200), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT77), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n482), .A2(new_n353), .ZN(new_n536));
  AND3_X1   g0336(.A1(new_n529), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n535), .B1(new_n529), .B2(new_n536), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n533), .A2(G169), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n512), .A2(G179), .A3(new_n515), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n520), .A2(new_n534), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT6), .ZN(new_n544));
  NOR3_X1   g0344(.A1(new_n544), .A2(new_n206), .A3(G107), .ZN(new_n545));
  XNOR2_X1  g0345(.A(G97), .B(G107), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n545), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  OAI22_X1  g0347(.A1(new_n547), .A2(new_n223), .B1(new_n356), .B2(new_n393), .ZN(new_n548));
  INV_X1    g0348(.A(G107), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n386), .B2(new_n388), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n282), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n482), .A2(G97), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n284), .A2(new_n206), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(G244), .B1(new_n320), .B2(new_n321), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT4), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n555), .A2(new_n556), .B1(G33), .B2(G283), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n250), .A2(KEYINPUT4), .A3(G244), .A4(new_n251), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n556), .B1(new_n250), .B2(G250), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n560), .A2(new_n251), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n257), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n474), .A2(new_n207), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n562), .A2(new_n455), .A3(new_n479), .A4(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n479), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n557), .B(new_n558), .C1(new_n251), .C2(new_n560), .ZN(new_n567));
  AOI211_X1 g0367(.A(new_n563), .B(new_n566), .C1(new_n567), .C2(new_n257), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n554), .B(new_n565), .C1(new_n568), .C2(G169), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n562), .A2(new_n479), .A3(new_n564), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G200), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n563), .B1(new_n567), .B2(new_n257), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n573), .A2(G190), .A3(new_n479), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n571), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n543), .A2(new_n569), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n482), .A2(G107), .ZN(new_n577));
  AOI21_X1  g0377(.A(KEYINPUT25), .B1(new_n284), .B2(new_n549), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n284), .A2(KEYINPUT25), .A3(new_n549), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n577), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n250), .A2(G257), .A3(G1698), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n250), .A2(G250), .A3(new_n251), .ZN(new_n583));
  XNOR2_X1  g0383(.A(KEYINPUT84), .B(G294), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n582), .B(new_n583), .C1(new_n247), .C2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n257), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n473), .A2(G264), .A3(new_n256), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n479), .A3(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n589), .A2(new_n268), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT83), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n510), .A2(G20), .ZN(new_n592));
  AND3_X1   g0392(.A1(new_n549), .A2(KEYINPUT23), .A3(G20), .ZN(new_n593));
  AOI21_X1  g0393(.A(KEYINPUT23), .B1(new_n549), .B2(G20), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n223), .B(G87), .C1(new_n320), .C2(new_n321), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT22), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT22), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n250), .A2(new_n598), .A3(new_n223), .A4(G87), .ZN(new_n599));
  AOI211_X1 g0399(.A(new_n592), .B(new_n595), .C1(new_n597), .C2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT24), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n591), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT82), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n600), .A2(new_n603), .A3(new_n601), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n597), .A2(new_n599), .ZN(new_n605));
  INV_X1    g0405(.A(new_n592), .ZN(new_n606));
  INV_X1    g0406(.A(new_n595), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n605), .A2(new_n601), .A3(new_n606), .A4(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(KEYINPUT82), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n610), .A2(KEYINPUT83), .A3(KEYINPUT24), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n602), .A2(new_n604), .A3(new_n609), .A4(new_n611), .ZN(new_n612));
  AOI211_X1 g0412(.A(new_n581), .B(new_n590), .C1(new_n612), .C2(new_n282), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n589), .A2(G200), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n612), .A2(new_n282), .ZN(new_n615));
  INV_X1    g0415(.A(new_n581), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n589), .A2(new_n453), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n618), .B1(G179), .B2(new_n589), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n613), .A2(new_n614), .B1(new_n617), .B2(new_n620), .ZN(new_n621));
  AND4_X1   g0421(.A1(new_n460), .A2(new_n504), .A3(new_n576), .A4(new_n621), .ZN(G372));
  INV_X1    g0422(.A(KEYINPUT26), .ZN(new_n623));
  INV_X1    g0423(.A(new_n569), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n623), .B1(new_n543), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n529), .A2(new_n536), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n542), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n533), .A2(G200), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n628), .A2(new_n529), .A3(new_n530), .A4(new_n516), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n630), .A2(KEYINPUT26), .A3(new_n569), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n625), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n575), .A2(new_n569), .A3(new_n629), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n590), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n615), .A2(new_n616), .A3(new_n614), .A4(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n496), .A2(new_n498), .A3(new_n500), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n619), .B1(new_n615), .B2(new_n616), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n634), .B(new_n636), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n632), .A2(new_n639), .A3(new_n627), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n460), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n335), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n343), .A2(new_n344), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n642), .B1(new_n458), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n445), .A2(new_n450), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n433), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n305), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n648), .A2(new_n349), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n641), .A2(new_n649), .ZN(G369));
  NAND3_X1  g0450(.A1(new_n259), .A2(new_n223), .A3(G13), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n651), .B(KEYINPUT85), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT27), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(new_n655), .A3(G213), .ZN(new_n656));
  INV_X1    g0456(.A(G343), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n504), .B1(new_n502), .B2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n637), .A2(new_n492), .A3(new_n658), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(G330), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n617), .A2(new_n658), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n638), .B1(new_n664), .B2(new_n636), .ZN(new_n665));
  INV_X1    g0465(.A(new_n282), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n610), .A2(KEYINPUT83), .A3(KEYINPUT24), .ZN(new_n667));
  AOI21_X1  g0467(.A(KEYINPUT83), .B1(new_n610), .B2(KEYINPUT24), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n608), .B(new_n603), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n666), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n620), .B1(new_n671), .B2(new_n581), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(new_n658), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n665), .A2(new_n673), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n493), .A2(new_n494), .A3(new_n497), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n497), .B1(new_n493), .B2(new_n494), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n658), .B1(new_n677), .B2(new_n500), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n663), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n673), .B1(new_n621), .B2(new_n678), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(G399));
  NOR2_X1   g0483(.A1(new_n523), .A2(G116), .ZN(new_n684));
  XOR2_X1   g0484(.A(new_n684), .B(KEYINPUT86), .Z(new_n685));
  INV_X1    g0485(.A(new_n226), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(G41), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n685), .A2(new_n688), .A3(G1), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n222), .B2(new_n688), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT28), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT88), .ZN(new_n692));
  INV_X1    g0492(.A(new_n627), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n672), .A2(new_n677), .A3(new_n500), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n633), .B1(new_n613), .B2(new_n614), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n658), .B1(new_n696), .B2(new_n632), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n692), .B1(new_n697), .B2(KEYINPUT29), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n640), .A2(new_n659), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT29), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(KEYINPUT88), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(KEYINPUT26), .B1(new_n630), .B2(new_n569), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n543), .A2(new_n623), .A3(new_n624), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n639), .A2(new_n627), .A3(new_n702), .A4(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n704), .A2(KEYINPUT29), .A3(new_n659), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n698), .A2(new_n701), .A3(new_n705), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n621), .A2(new_n576), .A3(new_n504), .A4(new_n659), .ZN(new_n707));
  INV_X1    g0507(.A(new_n541), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n499), .A2(new_n708), .A3(new_n573), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT30), .ZN(new_n710));
  OR3_X1    g0510(.A1(new_n709), .A2(new_n710), .A3(new_n589), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n710), .B1(new_n709), .B2(new_n589), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n570), .A2(new_n480), .A3(new_n589), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(new_n455), .A3(new_n533), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n711), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  AOI22_X1  g0515(.A1(new_n707), .A2(KEYINPUT31), .B1(new_n658), .B2(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n712), .A2(new_n714), .A3(KEYINPUT87), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n711), .ZN(new_n718));
  AOI21_X1  g0518(.A(KEYINPUT87), .B1(new_n712), .B2(new_n714), .ZN(new_n719));
  OAI211_X1 g0519(.A(KEYINPUT31), .B(new_n658), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(G330), .B1(new_n716), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n706), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n691), .B1(new_n724), .B2(G1), .ZN(G364));
  AOI21_X1  g0525(.A(new_n224), .B1(G20), .B2(new_n453), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n726), .A2(KEYINPUT91), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(KEYINPUT91), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n223), .A2(new_n268), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n455), .A2(G200), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(G322), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n455), .A2(new_n375), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n730), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  XOR2_X1   g0537(.A(KEYINPUT92), .B(G326), .Z(new_n738));
  NOR2_X1   g0538(.A1(G179), .A2(G200), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G190), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G20), .ZN(new_n741));
  AOI22_X1  g0541(.A1(new_n737), .A2(new_n738), .B1(new_n741), .B2(new_n584), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(KEYINPUT93), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n223), .A2(G190), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n731), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI211_X1 g0546(.A(new_n250), .B(new_n743), .C1(G311), .C2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n375), .A2(G179), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n730), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G303), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n735), .A2(new_n744), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(G317), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(KEYINPUT33), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n754), .A2(KEYINPUT33), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n753), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n748), .A2(new_n744), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n744), .A2(new_n739), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI22_X1  g0561(.A1(G283), .A2(new_n759), .B1(new_n761), .B2(G329), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT94), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n747), .A2(new_n751), .A3(new_n757), .A4(new_n763), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n734), .B(new_n764), .C1(KEYINPUT93), .C2(new_n742), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n737), .A2(G50), .B1(new_n746), .B2(G77), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n766), .B1(new_n549), .B2(new_n758), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n760), .A2(new_n394), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT32), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n741), .A2(G97), .ZN(new_n770));
  INV_X1    g0570(.A(new_n732), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(new_n273), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n362), .B1(new_n750), .B2(G87), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n769), .A2(new_n770), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n767), .B(new_n774), .C1(G68), .C2(new_n753), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n729), .B1(new_n765), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n283), .A2(G20), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n259), .B1(new_n777), .B2(G45), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n687), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G13), .A2(G33), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT90), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G20), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n729), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  OR2_X1    g0586(.A1(new_n222), .A2(G45), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n686), .A2(new_n250), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n787), .B(new_n788), .C1(new_n241), .C2(new_n469), .ZN(new_n789));
  INV_X1    g0589(.A(G355), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n250), .A2(new_n226), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n789), .B1(G116), .B2(new_n226), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT89), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n776), .B(new_n780), .C1(new_n786), .C2(new_n793), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT95), .ZN(new_n795));
  INV_X1    g0595(.A(new_n784), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n795), .B1(new_n662), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(G330), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n798), .B1(new_n660), .B2(new_n661), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(new_n780), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(G330), .B2(new_n662), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(G396));
  AND4_X1   g0603(.A1(new_n452), .A2(new_n454), .A3(new_n456), .A4(new_n659), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n373), .A2(new_n376), .B1(new_n361), .B2(new_n659), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n804), .B1(new_n805), .B2(new_n457), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n640), .A2(new_n659), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(KEYINPUT98), .ZN(new_n808));
  INV_X1    g0608(.A(new_n806), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n699), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n808), .B(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n722), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n812), .A2(KEYINPUT99), .ZN(new_n813));
  INV_X1    g0613(.A(new_n780), .ZN(new_n814));
  OR2_X1    g0614(.A1(new_n811), .A2(new_n722), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n812), .A2(KEYINPUT99), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n813), .A2(new_n814), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(G303), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n770), .B1(new_n549), .B2(new_n749), .C1(new_n818), .C2(new_n736), .ZN(new_n819));
  INV_X1    g0619(.A(G311), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n758), .A2(new_n522), .B1(new_n760), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n362), .B1(new_n745), .B2(new_n484), .ZN(new_n822));
  NOR3_X1   g0622(.A1(new_n819), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(G283), .ZN(new_n824));
  INV_X1    g0624(.A(G294), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n823), .B1(new_n824), .B2(new_n752), .C1(new_n825), .C2(new_n732), .ZN(new_n826));
  XOR2_X1   g0626(.A(KEYINPUT97), .B(G143), .Z(new_n827));
  AOI22_X1  g0627(.A1(new_n771), .A2(new_n827), .B1(new_n746), .B2(G159), .ZN(new_n828));
  INV_X1    g0628(.A(G137), .ZN(new_n829));
  INV_X1    g0629(.A(G150), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n828), .B1(new_n829), .B2(new_n736), .C1(new_n830), .C2(new_n752), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT34), .ZN(new_n832));
  INV_X1    g0632(.A(new_n273), .ZN(new_n833));
  INV_X1    g0633(.A(new_n741), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n832), .B1(new_n204), .B2(new_n758), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(G132), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n250), .B1(new_n760), .B2(new_n836), .C1(new_n276), .C2(new_n749), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n826), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n729), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n729), .A2(new_n781), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n814), .B1(new_n840), .B2(new_n356), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n841), .B(KEYINPUT96), .Z(new_n842));
  OAI211_X1 g0642(.A(new_n839), .B(new_n842), .C1(new_n806), .C2(new_n783), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n817), .A2(new_n843), .ZN(G384));
  INV_X1    g0644(.A(KEYINPUT35), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n223), .B(new_n224), .C1(new_n547), .C2(new_n845), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n846), .B(G116), .C1(new_n845), .C2(new_n547), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT36), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n204), .A2(G50), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n849), .B(KEYINPUT100), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n399), .A2(G77), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n850), .B1(new_n222), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n852), .A2(G1), .A3(new_n283), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT103), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT38), .ZN(new_n855));
  AND3_X1   g0655(.A1(new_n656), .A2(new_n423), .A3(new_n426), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n392), .A2(new_n402), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n405), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n858), .A2(new_n282), .A3(new_n403), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n856), .B1(new_n859), .B2(new_n382), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n438), .B1(new_n404), .B2(new_n416), .ZN(new_n861));
  OAI21_X1  g0661(.A(KEYINPUT37), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT37), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n447), .B(new_n863), .C1(new_n417), .C2(new_n856), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n656), .B1(new_n859), .B2(new_n382), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n855), .B(new_n865), .C1(new_n451), .C2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n451), .A2(new_n866), .ZN(new_n868));
  INV_X1    g0668(.A(new_n865), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT38), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n854), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT102), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n804), .B1(new_n697), .B2(new_n806), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n344), .A2(new_n658), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n345), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT101), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n345), .A2(KEYINPUT101), .A3(new_n874), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n877), .A2(new_n878), .B1(new_n644), .B2(new_n658), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n872), .B1(new_n873), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n868), .A2(new_n869), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n855), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n868), .A2(KEYINPUT38), .A3(new_n869), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n882), .A2(KEYINPUT103), .A3(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n804), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n807), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n644), .A2(new_n658), .ZN(new_n887));
  AND4_X1   g0687(.A1(KEYINPUT101), .A2(new_n643), .A3(new_n642), .A4(new_n874), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT101), .B1(new_n345), .B2(new_n874), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n886), .A2(KEYINPUT102), .A3(new_n890), .ZN(new_n891));
  AND4_X1   g0691(.A1(new_n871), .A2(new_n880), .A3(new_n884), .A4(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT39), .ZN(new_n893));
  OAI21_X1  g0693(.A(KEYINPUT104), .B1(new_n439), .B2(new_n444), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT104), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n448), .A2(new_n895), .A3(new_n449), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n433), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n417), .ZN(new_n898));
  INV_X1    g0698(.A(new_n656), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n447), .B1(new_n417), .B2(new_n856), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT37), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n864), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT38), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n893), .B1(new_n904), .B2(new_n867), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n882), .A2(KEYINPUT39), .A3(new_n883), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n644), .A2(new_n659), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n905), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n433), .A2(new_n899), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(KEYINPUT105), .B1(new_n892), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n912), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT105), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n880), .A2(new_n871), .A3(new_n891), .A4(new_n884), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n460), .A2(new_n705), .A3(new_n698), .A4(new_n701), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n649), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n918), .B(new_n920), .Z(new_n921));
  AND3_X1   g0721(.A1(new_n715), .A2(KEYINPUT31), .A3(new_n658), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n707), .A2(KEYINPUT31), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n715), .A2(new_n658), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n890), .A2(new_n806), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n927), .A2(new_n884), .A3(new_n871), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT40), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n904), .A2(new_n867), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n930), .A2(new_n929), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n928), .A2(new_n929), .B1(new_n931), .B2(new_n927), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n932), .B(new_n460), .C1(new_n716), .C2(new_n922), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n928), .A2(new_n929), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n931), .A2(new_n927), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n934), .A2(G330), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(G330), .B1(new_n716), .B2(new_n922), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n460), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n933), .A2(new_n940), .ZN(new_n941));
  OAI22_X1  g0741(.A1(new_n921), .A2(new_n941), .B1(new_n259), .B2(new_n777), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT106), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n921), .A2(new_n941), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n848), .B(new_n853), .C1(new_n943), .C2(new_n944), .ZN(G367));
  OAI211_X1 g0745(.A(new_n575), .B(new_n569), .C1(new_n572), .C2(new_n659), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n569), .B2(new_n659), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n680), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n678), .A2(new_n621), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n949), .A2(new_n946), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT42), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n569), .B1(new_n672), .B2(new_n946), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n659), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n658), .A2(new_n531), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n693), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n630), .B2(new_n955), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(KEYINPUT108), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT107), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n954), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n958), .A2(KEYINPUT108), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n963), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n954), .A2(new_n965), .A3(new_n959), .A4(new_n961), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n948), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT109), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n964), .A2(new_n948), .A3(new_n966), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n687), .B(KEYINPUT41), .Z(new_n970));
  INV_X1    g0770(.A(KEYINPUT111), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n680), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n679), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n799), .B1(new_n973), .B2(new_n949), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(KEYINPUT111), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT110), .ZN(new_n978));
  NOR3_X1   g0778(.A1(new_n977), .A2(new_n978), .A3(new_n723), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n682), .A2(new_n947), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT44), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n682), .A2(new_n947), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT45), .ZN(new_n984));
  OR3_X1    g0784(.A1(new_n982), .A2(new_n680), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n979), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n970), .B1(new_n986), .B2(new_n724), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n968), .B(new_n969), .C1(new_n987), .C2(new_n779), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n834), .A2(new_n549), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n362), .B1(new_n760), .B2(new_n754), .C1(new_n206), .C2(new_n758), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n991), .A2(KEYINPUT112), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT46), .ZN(new_n993));
  NOR3_X1   g0793(.A1(new_n749), .A2(new_n993), .A3(new_n484), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n585), .A2(new_n752), .B1(new_n736), .B2(new_n820), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n994), .B(new_n995), .C1(G283), .C2(new_n746), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n993), .B1(new_n749), .B2(new_n484), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n991), .A2(KEYINPUT112), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n992), .A2(new_n996), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n989), .B(new_n999), .C1(G303), .C2(new_n771), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n771), .A2(G150), .B1(new_n741), .B2(G68), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(KEYINPUT113), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(G159), .A2(new_n753), .B1(new_n759), .B2(G77), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n1002), .B2(KEYINPUT113), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n737), .A2(new_n827), .B1(new_n746), .B2(G50), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1006), .B(new_n250), .C1(new_n833), .C2(new_n749), .ZN(new_n1007));
  XOR2_X1   g0807(.A(KEYINPUT114), .B(G137), .Z(new_n1008));
  NOR2_X1   g0808(.A1(new_n1008), .A2(new_n760), .ZN(new_n1009));
  NOR3_X1   g0809(.A1(new_n1005), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1000), .B1(new_n1003), .B2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT47), .Z(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n729), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n957), .A2(new_n796), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n788), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n785), .B1(new_n226), .B2(new_n354), .C1(new_n237), .C2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1013), .A2(new_n780), .A3(new_n1014), .A4(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n988), .A2(new_n1017), .ZN(G387));
  INV_X1    g0818(.A(new_n977), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n724), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n688), .B1(new_n977), .B2(new_n723), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n784), .B1(new_n665), .B2(new_n673), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n729), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G322), .A2(new_n737), .B1(new_n753), .B2(G311), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1025), .B1(new_n818), .B2(new_n745), .C1(new_n754), .C2(new_n732), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT48), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(new_n824), .B2(new_n834), .C1(new_n585), .C2(new_n749), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT49), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n761), .A2(new_n738), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n250), .B1(new_n759), .B2(G116), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n274), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n1033), .A2(new_n752), .B1(new_n204), .B2(new_n745), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(G50), .B2(new_n771), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n834), .A2(new_n354), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n736), .A2(new_n394), .B1(new_n760), .B2(new_n830), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n750), .A2(G77), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n362), .B1(new_n759), .B2(G97), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1035), .A2(new_n1038), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1024), .B1(new_n1032), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n788), .B1(new_n233), .B2(new_n469), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n685), .B2(new_n791), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n685), .B(new_n469), .C1(new_n204), .C2(new_n356), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n351), .A2(new_n276), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT50), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1044), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n686), .A2(new_n549), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n786), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NOR3_X1   g0850(.A1(new_n1042), .A2(new_n814), .A3(new_n1050), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n1019), .A2(new_n779), .B1(new_n1023), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1022), .A2(new_n1052), .ZN(G393));
  OAI21_X1  g0853(.A(new_n680), .B1(new_n982), .B2(new_n984), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n985), .A2(new_n1054), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n1020), .A2(new_n1055), .B1(new_n979), .B2(new_n985), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n985), .A2(new_n779), .A3(new_n1054), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n785), .B1(new_n244), .B2(new_n1015), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G97), .B2(new_n686), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n736), .A2(new_n754), .B1(new_n732), .B2(new_n820), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT52), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n834), .A2(new_n484), .B1(new_n825), .B2(new_n745), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n362), .B1(new_n752), .B2(new_n818), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n758), .A2(new_n549), .B1(new_n760), .B2(new_n733), .ZN(new_n1064));
  NOR3_X1   g0864(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1061), .B(new_n1065), .C1(new_n824), .C2(new_n749), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n753), .A2(G50), .B1(new_n746), .B2(new_n351), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT115), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1069), .B(new_n1070), .C1(new_n356), .C2(new_n834), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1071), .B(KEYINPUT116), .Z(new_n1072));
  NAND2_X1  g0872(.A1(new_n761), .A2(new_n827), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G68), .A2(new_n750), .B1(new_n759), .B2(G87), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1072), .A2(new_n250), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n736), .A2(new_n830), .B1(new_n732), .B2(new_n394), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT51), .Z(new_n1077));
  OAI21_X1  g0877(.A(new_n1066), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n814), .B(new_n1059), .C1(new_n1078), .C2(new_n729), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n796), .B2(new_n947), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1057), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT117), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1057), .A2(KEYINPUT117), .A3(new_n1080), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n1056), .A2(new_n687), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(G390));
  NOR2_X1   g0886(.A1(new_n879), .A2(new_n809), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1087), .B(G330), .C1(new_n716), .C2(new_n922), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n886), .A2(new_n890), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n907), .A2(new_n1089), .B1(new_n905), .B2(new_n906), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n904), .A2(new_n867), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n805), .A2(new_n457), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n704), .A2(new_n659), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n885), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n890), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n907), .B(KEYINPUT118), .ZN(new_n1096));
  AND3_X1   g0896(.A1(new_n1091), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1088), .B1(new_n1090), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1089), .A2(new_n907), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n905), .A2(new_n906), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  OAI211_X1 g0901(.A(G330), .B(new_n806), .C1(new_n716), .C2(new_n721), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1102), .A2(new_n879), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1091), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1101), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1098), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n919), .A2(new_n939), .A3(new_n649), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1102), .A2(new_n879), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1088), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n886), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n879), .B1(new_n937), .B2(new_n809), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1094), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1112), .B(new_n1113), .C1(new_n879), .C2(new_n1102), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1108), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT119), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AOI211_X1 g0917(.A(KEYINPUT119), .B(new_n1108), .C1(new_n1111), .C2(new_n1114), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1107), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1106), .A2(new_n1115), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1119), .A2(new_n687), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n778), .B1(new_n1098), .B2(new_n1105), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1100), .A2(new_n782), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n362), .B1(new_n749), .B2(new_n522), .ZN(new_n1124));
  XOR2_X1   g0924(.A(new_n1124), .B(KEYINPUT120), .Z(new_n1125));
  OAI22_X1  g0925(.A1(new_n834), .A2(new_n356), .B1(new_n204), .B2(new_n758), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n752), .A2(new_n549), .B1(new_n745), .B2(new_n206), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n736), .A2(new_n824), .ZN(new_n1128));
  NOR4_X1   g0928(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1129), .B1(new_n484), .B2(new_n732), .C1(new_n825), .C2(new_n760), .ZN(new_n1130));
  OAI21_X1  g0930(.A(KEYINPUT53), .B1(new_n749), .B2(new_n830), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n394), .B2(new_n834), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n250), .B1(new_n758), .B2(new_n276), .C1(new_n752), .C2(new_n1008), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n749), .A2(KEYINPUT53), .A3(new_n830), .ZN(new_n1134));
  NOR3_X1   g0934(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n737), .A2(G128), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n761), .A2(G125), .ZN(new_n1137));
  XOR2_X1   g0937(.A(KEYINPUT54), .B(G143), .Z(new_n1138));
  AOI22_X1  g0938(.A1(G132), .A2(new_n771), .B1(new_n746), .B2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .A4(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1024), .B1(new_n1130), .B2(new_n1140), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n814), .B(new_n1141), .C1(new_n1033), .C2(new_n840), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1123), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  OR3_X1    g0944(.A1(new_n1122), .A2(KEYINPUT121), .A3(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(KEYINPUT121), .B1(new_n1122), .B2(new_n1144), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1121), .A2(new_n1147), .ZN(G378));
  NAND2_X1  g0948(.A1(new_n305), .A2(new_n349), .ZN(new_n1149));
  XOR2_X1   g0949(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1149), .B(new_n1151), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n293), .A2(new_n656), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1149), .B(new_n1150), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1153), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AND2_X1   g0957(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n936), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n932), .A2(new_n1160), .A3(G330), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n918), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1159), .A2(new_n913), .A3(new_n917), .A4(new_n1161), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n840), .A2(new_n276), .ZN(new_n1166));
  AOI21_X1  g0966(.A(G50), .B1(new_n249), .B2(new_n255), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n833), .A2(new_n758), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n732), .A2(new_n549), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT122), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n761), .A2(G283), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1169), .A2(new_n1172), .A3(new_n1039), .A4(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n752), .A2(new_n206), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n255), .B1(new_n834), .B2(new_n204), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n362), .B1(new_n736), .B2(new_n484), .ZN(new_n1177));
  NOR4_X1   g0977(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1178), .B1(new_n1171), .B2(new_n1170), .C1(new_n354), .C2(new_n745), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT58), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(G128), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n732), .A2(new_n1182), .B1(new_n745), .B2(new_n829), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1138), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n834), .A2(new_n830), .B1(new_n1184), .B2(new_n749), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n1183), .B(new_n1185), .C1(G125), .C2(new_n737), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n836), .B2(new_n752), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(KEYINPUT59), .ZN(new_n1188));
  OR2_X1    g0988(.A1(KEYINPUT123), .A2(G124), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(KEYINPUT123), .A2(G124), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n761), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n255), .B(new_n1191), .C1(new_n1187), .C2(KEYINPUT59), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n758), .A2(new_n394), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1192), .A2(G33), .A3(new_n1193), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1167), .B(new_n1181), .C1(new_n1188), .C2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n780), .B1(new_n1195), .B2(new_n1024), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(new_n1160), .B2(new_n782), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1165), .A2(new_n779), .B1(new_n1166), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1108), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1120), .A2(new_n1199), .ZN(new_n1200));
  AND4_X1   g1000(.A1(new_n917), .A2(new_n1159), .A3(new_n913), .A4(new_n1161), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1159), .A2(new_n1161), .B1(new_n913), .B2(new_n917), .ZN(new_n1202));
  OAI211_X1 g1002(.A(KEYINPUT57), .B(new_n1200), .C1(new_n1201), .C2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n687), .ZN(new_n1204));
  AOI21_X1  g1004(.A(KEYINPUT57), .B1(new_n1165), .B2(new_n1200), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1198), .B1(new_n1204), .B2(new_n1205), .ZN(G375));
  OAI221_X1 g1006(.A(new_n362), .B1(new_n745), .B2(new_n549), .C1(new_n206), .C2(new_n749), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n736), .A2(new_n825), .B1(new_n758), .B2(new_n356), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n760), .A2(new_n818), .ZN(new_n1209));
  NOR4_X1   g1009(.A1(new_n1207), .A2(new_n1036), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1210), .B1(new_n484), .B2(new_n752), .C1(new_n824), .C2(new_n732), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n736), .A2(new_n836), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n1184), .A2(new_n752), .B1(new_n732), .B2(new_n1008), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(G150), .C2(new_n746), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n741), .A2(G50), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n749), .A2(new_n394), .B1(new_n760), .B2(new_n1182), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1216), .B(KEYINPUT124), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1214), .A2(new_n250), .A3(new_n1215), .A4(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1211), .B1(new_n1218), .B2(new_n1168), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n814), .B1(new_n1219), .B2(new_n729), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n840), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1220), .B1(G68), .B2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n879), .B2(new_n781), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1223), .B1(new_n1224), .B2(new_n779), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1111), .A2(new_n1108), .A3(new_n1114), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n1118), .B2(new_n1117), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1225), .B1(new_n1227), .B2(new_n970), .ZN(G381));
  OAI21_X1  g1028(.A(new_n779), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1197), .A2(new_n1166), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1108), .B1(new_n1106), .B2(new_n1224), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n688), .B1(new_n1233), .B2(KEYINPUT57), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1200), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT57), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1231), .B1(new_n1234), .B2(new_n1237), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1122), .A2(new_n1144), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1121), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1238), .A2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n988), .A2(new_n1017), .A3(new_n1085), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(new_n1241), .A2(G381), .A3(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(G384), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(G393), .A2(G396), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .ZN(G407));
  NAND2_X1  g1046(.A1(new_n657), .A2(G213), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(KEYINPUT125), .ZN(new_n1248));
  OAI211_X1 g1048(.A(G407), .B(G213), .C1(new_n1241), .C2(new_n1248), .ZN(G409));
  AOI21_X1  g1049(.A(new_n802), .B1(new_n1022), .B2(new_n1052), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1245), .A2(new_n1250), .ZN(new_n1251));
  AND3_X1   g1051(.A1(new_n988), .A2(new_n1017), .A3(new_n1085), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1085), .B1(new_n988), .B2(new_n1017), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1251), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(G387), .A2(G390), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1251), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1255), .A2(new_n1242), .A3(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1254), .A2(new_n1257), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1235), .A2(new_n970), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1240), .B1(new_n1231), .B2(new_n1259), .ZN(new_n1260));
  OAI211_X1 g1060(.A(G378), .B(new_n1198), .C1(new_n1204), .C2(new_n1205), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT60), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n688), .B1(new_n1226), .B2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1115), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1264), .B(new_n1265), .C1(new_n1263), .C2(new_n1226), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n1225), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1244), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1266), .A2(G384), .A3(new_n1225), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1262), .A2(new_n1247), .A3(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT62), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1248), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1274), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1270), .A2(new_n1273), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n1272), .A2(new_n1273), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT61), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n657), .A2(G213), .A3(G2897), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1248), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n1271), .A2(new_n1279), .B1(new_n1280), .B2(G2897), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1278), .B1(new_n1282), .B2(new_n1275), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1258), .B1(new_n1277), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT63), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1270), .A2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1258), .B1(new_n1275), .B2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1262), .A2(new_n1247), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1285), .B1(new_n1288), .B2(new_n1281), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1272), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1287), .B(new_n1278), .C1(new_n1289), .C2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1284), .A2(new_n1291), .ZN(G405));
  AND2_X1   g1092(.A1(new_n1254), .A2(new_n1257), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1240), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1261), .B(new_n1270), .C1(new_n1238), .C2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(G375), .A2(new_n1240), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1270), .B1(new_n1297), .B2(new_n1261), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1293), .B1(new_n1296), .B2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT127), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  OAI211_X1 g1101(.A(new_n1293), .B(KEYINPUT127), .C1(new_n1296), .C2(new_n1298), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1261), .B1(new_n1238), .B2(new_n1294), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1271), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1304), .A2(new_n1258), .A3(new_n1295), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(KEYINPUT126), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT126), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1304), .A2(new_n1307), .A3(new_n1258), .A4(new_n1295), .ZN(new_n1308));
  AOI22_X1  g1108(.A1(new_n1301), .A2(new_n1302), .B1(new_n1306), .B2(new_n1308), .ZN(G402));
endmodule


