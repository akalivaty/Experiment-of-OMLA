//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 0 0 0 1 1 1 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 1 0 0 1 1 0 1 1 0 0 0 0 0 0 0 0 1 0 0 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n841, new_n842,
    new_n843, new_n845, new_n846, new_n847, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961;
  XOR2_X1   g000(.A(KEYINPUT92), .B(KEYINPUT15), .Z(new_n202));
  INV_X1    g001(.A(G43gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G50gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT93), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n203), .A2(G50gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n202), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n204), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT15), .ZN(new_n210));
  NOR3_X1   g009(.A1(new_n209), .A2(new_n207), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(G29gat), .A2(G36gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT14), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n213), .B(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G29gat), .A2(G36gat), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n208), .A2(new_n212), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT91), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n213), .A2(new_n218), .A3(new_n214), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(new_n216), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n211), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n217), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n223), .B(KEYINPUT17), .ZN(new_n224));
  XOR2_X1   g023(.A(G15gat), .B(G22gat), .Z(new_n225));
  INV_X1    g024(.A(G1gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT94), .ZN(new_n228));
  XNOR2_X1  g027(.A(G15gat), .B(G22gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT16), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n229), .B1(new_n230), .B2(G1gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n228), .A2(new_n232), .A3(G8gat), .ZN(new_n233));
  INV_X1    g032(.A(G8gat), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n227), .B(new_n231), .C1(KEYINPUT94), .C2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n224), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT95), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n236), .B(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(new_n223), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(G229gat), .A2(G233gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n242), .A2(KEYINPUT18), .A3(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n240), .B(new_n223), .ZN(new_n245));
  XOR2_X1   g044(.A(new_n243), .B(KEYINPUT13), .Z(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n238), .A2(new_n241), .A3(new_n243), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT18), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n244), .A2(new_n247), .A3(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G113gat), .B(G141gat), .ZN(new_n252));
  INV_X1    g051(.A(G197gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT11), .B(G169gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n256), .B(KEYINPUT12), .Z(new_n257));
  NAND2_X1  g056(.A1(new_n251), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n257), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n244), .A2(new_n247), .A3(new_n250), .A4(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT77), .ZN(new_n263));
  INV_X1    g062(.A(G141gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n264), .A2(G148gat), .ZN(new_n265));
  INV_X1    g064(.A(G148gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n266), .A2(G141gat), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n263), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT2), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n266), .A2(G141gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n264), .A2(G148gat), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n270), .A2(new_n271), .A3(KEYINPUT77), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n268), .A2(new_n269), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(G155gat), .A2(G162gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(G155gat), .A2(G162gat), .ZN(new_n275));
  XOR2_X1   g074(.A(new_n275), .B(KEYINPUT76), .Z(new_n276));
  NAND3_X1  g075(.A1(new_n273), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n269), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(new_n274), .ZN(new_n279));
  XOR2_X1   g078(.A(KEYINPUT78), .B(G141gat), .Z(new_n280));
  NOR2_X1   g079(.A1(new_n280), .A2(new_n266), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT79), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n270), .B(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n279), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n277), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT72), .B(KEYINPUT22), .ZN(new_n286));
  INV_X1    g085(.A(G211gat), .ZN(new_n287));
  INV_X1    g086(.A(G218gat), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(G211gat), .B(G218gat), .Z(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G197gat), .B(G204gat), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n289), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  OR2_X1    g092(.A1(new_n293), .A2(KEYINPUT74), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(KEYINPUT74), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n289), .A2(new_n292), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n291), .B1(new_n297), .B2(KEYINPUT73), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n298), .B1(KEYINPUT73), .B2(new_n297), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT29), .B1(new_n296), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n285), .B1(new_n300), .B2(KEYINPUT3), .ZN(new_n301));
  AND2_X1   g100(.A1(G228gat), .A2(G233gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n296), .A2(new_n299), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT3), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n277), .A2(new_n284), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT29), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n301), .A2(new_n302), .A3(new_n309), .ZN(new_n310));
  AOI22_X1  g109(.A1(new_n294), .A2(new_n295), .B1(new_n290), .B2(new_n297), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n305), .B1(new_n311), .B2(KEYINPUT29), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(new_n285), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n302), .B1(new_n313), .B2(new_n309), .ZN(new_n314));
  OAI21_X1  g113(.A(G22gat), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n301), .A2(new_n302), .A3(new_n309), .ZN(new_n316));
  INV_X1    g115(.A(G22gat), .ZN(new_n317));
  AOI22_X1  g116(.A1(new_n312), .A2(new_n285), .B1(new_n304), .B2(new_n308), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n316), .B(new_n317), .C1(new_n302), .C2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n315), .A2(new_n319), .A3(KEYINPUT84), .ZN(new_n320));
  XNOR2_X1  g119(.A(G78gat), .B(G106gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(KEYINPUT31), .B(G50gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n321), .B(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n310), .A2(new_n314), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT84), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n325), .A2(new_n326), .A3(new_n317), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n320), .A2(new_n324), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n315), .A2(new_n319), .A3(new_n323), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT85), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n315), .A2(new_n319), .A3(KEYINPUT85), .A4(new_n323), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n328), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT83), .ZN(new_n334));
  INV_X1    g133(.A(G127gat), .ZN(new_n335));
  INV_X1    g134(.A(G134gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(G127gat), .A2(G134gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT66), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n337), .A2(KEYINPUT66), .A3(new_n338), .ZN(new_n342));
  XNOR2_X1  g141(.A(G113gat), .B(G120gat), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n341), .B(new_n342), .C1(KEYINPUT1), .C2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT68), .ZN(new_n345));
  INV_X1    g144(.A(G120gat), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n345), .B1(new_n346), .B2(G113gat), .ZN(new_n347));
  INV_X1    g146(.A(G113gat), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT67), .B1(new_n348), .B2(G120gat), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT67), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n350), .A2(new_n346), .A3(G113gat), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n348), .A2(KEYINPUT68), .A3(G120gat), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n347), .A2(new_n349), .A3(new_n351), .A4(new_n352), .ZN(new_n353));
  OR2_X1    g152(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n354));
  NAND2_X1  g153(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n353), .A2(new_n354), .A3(new_n339), .A4(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n344), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT4), .B1(new_n285), .B2(new_n357), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n344), .A2(new_n356), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT4), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n359), .A2(new_n360), .A3(new_n284), .A4(new_n277), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(G225gat), .A2(G233gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n285), .A2(KEYINPUT3), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n364), .A2(new_n357), .A3(new_n306), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n362), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n363), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n285), .A2(new_n357), .ZN(new_n368));
  AOI22_X1  g167(.A1(new_n277), .A2(new_n284), .B1(new_n356), .B2(new_n344), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT5), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  XOR2_X1   g171(.A(G57gat), .B(G85gat), .Z(new_n373));
  XNOR2_X1  g172(.A(G1gat), .B(G29gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n375), .B(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n362), .A2(new_n365), .A3(KEYINPUT5), .A4(new_n363), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n372), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT6), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT81), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n306), .A2(new_n357), .ZN(new_n384));
  AOI22_X1  g183(.A1(new_n384), .A2(new_n364), .B1(new_n358), .B2(new_n361), .ZN(new_n385));
  AOI22_X1  g184(.A1(new_n385), .A2(new_n363), .B1(KEYINPUT5), .B2(new_n370), .ZN(new_n386));
  INV_X1    g185(.A(new_n379), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n377), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n383), .B1(new_n388), .B2(new_n381), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n378), .B1(new_n372), .B2(new_n379), .ZN(new_n390));
  NOR3_X1   g189(.A1(new_n390), .A2(KEYINPUT81), .A3(KEYINPUT6), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  XOR2_X1   g191(.A(new_n380), .B(KEYINPUT82), .Z(new_n393));
  AOI21_X1  g192(.A(new_n382), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(G226gat), .ZN(new_n395));
  INV_X1    g194(.A(G233gat), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(G190gat), .ZN(new_n398));
  AND2_X1   g197(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n399));
  NOR2_X1   g198(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT28), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT27), .B(G183gat), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n404), .A2(KEYINPUT28), .A3(new_n398), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  AND2_X1   g205(.A1(G169gat), .A2(G176gat), .ZN(new_n407));
  NOR2_X1   g206(.A1(G169gat), .A2(G176gat), .ZN(new_n408));
  OR3_X1    g207(.A1(new_n407), .A2(new_n408), .A3(KEYINPUT26), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(KEYINPUT26), .ZN(new_n410));
  NAND2_X1  g209(.A1(G183gat), .A2(G190gat), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n406), .A2(new_n409), .A3(new_n410), .A4(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n407), .B1(KEYINPUT23), .B2(new_n408), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT24), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(G183gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n398), .ZN(new_n417));
  NAND3_X1  g216(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n415), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT64), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n420), .B1(new_n408), .B2(KEYINPUT23), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT23), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n422), .B(KEYINPUT64), .C1(G169gat), .C2(G176gat), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n413), .A2(new_n419), .A3(new_n421), .A4(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT25), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n424), .A2(KEYINPUT65), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT65), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n427), .A2(KEYINPUT25), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(KEYINPUT25), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n428), .B1(new_n424), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n412), .B1(new_n426), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n397), .B1(new_n431), .B2(new_n307), .ZN(new_n432));
  INV_X1    g231(.A(new_n397), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n424), .A2(new_n429), .ZN(new_n434));
  INV_X1    g233(.A(new_n428), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n424), .A2(KEYINPUT65), .A3(new_n425), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n433), .B1(new_n438), .B2(new_n412), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT75), .B1(new_n432), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT75), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT29), .B1(new_n438), .B2(new_n412), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n441), .B1(new_n442), .B2(new_n397), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n440), .A2(new_n304), .A3(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n303), .B1(new_n432), .B2(new_n439), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(G8gat), .B(G36gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(G64gat), .B(G92gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n447), .B(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n444), .A2(new_n445), .A3(new_n449), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(KEYINPUT30), .A3(new_n452), .ZN(new_n453));
  AOI211_X1 g252(.A(KEYINPUT30), .B(new_n449), .C1(new_n444), .C2(new_n445), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n334), .B1(new_n394), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n388), .A2(new_n383), .A3(new_n381), .ZN(new_n459));
  OR2_X1    g258(.A1(new_n380), .A2(KEYINPUT82), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT81), .B1(new_n390), .B2(KEYINPUT6), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n380), .A2(KEYINPUT82), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n459), .A2(new_n460), .A3(new_n461), .A4(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n382), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n465), .A2(KEYINPUT83), .A3(new_n456), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n333), .B1(new_n458), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT36), .ZN(new_n468));
  XNOR2_X1  g267(.A(G71gat), .B(G99gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n469), .B(KEYINPUT70), .ZN(new_n470));
  XOR2_X1   g269(.A(G15gat), .B(G43gat), .Z(new_n471));
  XNOR2_X1  g270(.A(new_n470), .B(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(G227gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n431), .A2(new_n357), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n438), .A2(new_n359), .A3(new_n412), .ZN(new_n475));
  AOI211_X1 g274(.A(new_n473), .B(new_n396), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n472), .B1(new_n476), .B2(KEYINPUT33), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n474), .A2(new_n475), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n473), .A2(new_n396), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT32), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n474), .B(new_n475), .C1(new_n473), .C2(new_n396), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n484), .B(KEYINPUT34), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT33), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n480), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n481), .A2(new_n488), .A3(new_n472), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n483), .A2(new_n486), .A3(KEYINPUT71), .A4(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n489), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n481), .B1(new_n488), .B2(new_n472), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n485), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n483), .A2(new_n486), .A3(new_n489), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n468), .B(new_n490), .C1(new_n495), .C2(KEYINPUT71), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n493), .A2(new_n494), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT36), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT86), .B1(new_n467), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT37), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n450), .B1(new_n446), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT38), .ZN(new_n503));
  OR3_X1    g302(.A1(new_n432), .A2(new_n439), .A3(new_n303), .ZN(new_n504));
  AND2_X1   g303(.A1(new_n440), .A2(new_n443), .ZN(new_n505));
  OAI211_X1 g304(.A(KEYINPUT37), .B(new_n504), .C1(new_n505), .C2(new_n304), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n502), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n390), .A2(KEYINPUT6), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n382), .B1(new_n508), .B2(new_n380), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n507), .A2(new_n509), .A3(new_n451), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n444), .A2(KEYINPUT37), .A3(new_n445), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n503), .B1(new_n502), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n333), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  NOR3_X1   g313(.A1(new_n385), .A2(KEYINPUT39), .A3(new_n363), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n515), .A2(new_n378), .ZN(new_n516));
  OR3_X1    g315(.A1(new_n368), .A2(new_n367), .A3(new_n369), .ZN(new_n517));
  OAI211_X1 g316(.A(KEYINPUT39), .B(new_n517), .C1(new_n385), .C2(new_n363), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT40), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(new_n380), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n516), .A2(KEYINPUT40), .A3(new_n518), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n524), .B(KEYINPUT88), .ZN(new_n525));
  AND3_X1   g324(.A1(new_n453), .A2(new_n455), .A3(KEYINPUT87), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT87), .B1(new_n453), .B2(new_n455), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n523), .B(new_n525), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n528), .A2(KEYINPUT89), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT89), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT87), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n452), .A2(KEYINPUT30), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n449), .B1(new_n444), .B2(new_n445), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n531), .B1(new_n534), .B2(new_n454), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n453), .A2(new_n455), .A3(KEYINPUT87), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n522), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n530), .B1(new_n537), .B2(new_n525), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n514), .B1(new_n529), .B2(new_n538), .ZN(new_n539));
  AND3_X1   g338(.A1(new_n328), .A2(new_n331), .A3(new_n332), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n465), .A2(KEYINPUT83), .A3(new_n456), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT83), .B1(new_n465), .B2(new_n456), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT86), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n496), .A2(new_n498), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n500), .A2(new_n539), .A3(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n490), .B1(new_n495), .B2(KEYINPUT71), .ZN(new_n548));
  AND2_X1   g347(.A1(new_n548), .A2(new_n333), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n526), .A2(new_n527), .ZN(new_n550));
  XOR2_X1   g349(.A(KEYINPUT90), .B(KEYINPUT35), .Z(new_n551));
  NOR2_X1   g350(.A1(new_n509), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n549), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n333), .A2(new_n497), .ZN(new_n554));
  NOR3_X1   g353(.A1(new_n541), .A2(new_n542), .A3(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT35), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n553), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n262), .B1(new_n547), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G127gat), .B(G155gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(G231gat), .A2(G233gat), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n559), .B(new_n560), .Z(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT96), .B(G211gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n236), .B(KEYINPUT95), .ZN(new_n567));
  XNOR2_X1  g366(.A(G57gat), .B(G64gat), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G71gat), .B(G78gat), .ZN(new_n571));
  OR2_X1    g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n571), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT21), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n567), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(G183gat), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n567), .A2(new_n416), .A3(new_n576), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n575), .A2(KEYINPUT21), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n580), .A2(new_n581), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n566), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n584), .ZN(new_n586));
  NOR3_X1   g385(.A1(new_n586), .A2(new_n565), .A3(new_n582), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n562), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G85gat), .A2(G92gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT7), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT8), .ZN(new_n591));
  AND2_X1   g390(.A1(G99gat), .A2(G106gat), .ZN(new_n592));
  OAI221_X1 g391(.A(new_n590), .B1(new_n591), .B2(new_n592), .C1(G85gat), .C2(G92gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(G99gat), .B(G106gat), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n593), .B(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n224), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n593), .B(new_n594), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(new_n223), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n597), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G190gat), .B(G218gat), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n601), .B(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(G134gat), .B(G162gat), .Z(new_n605));
  AOI21_X1  g404(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n604), .B(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n565), .B1(new_n586), .B2(new_n582), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n583), .A2(new_n566), .A3(new_n584), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n609), .A2(new_n610), .A3(new_n561), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n588), .A2(new_n608), .A3(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT97), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n588), .A2(new_n608), .A3(KEYINPUT97), .A4(new_n611), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(G230gat), .A2(G233gat), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n596), .A2(new_n574), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n599), .A2(new_n575), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT10), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n599), .A2(KEYINPUT10), .A3(new_n575), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n618), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n617), .B1(new_n619), .B2(new_n620), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT98), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n625), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G120gat), .B(G148gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(G176gat), .B(G204gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n633), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n625), .A2(new_n628), .A3(new_n635), .A4(new_n629), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT99), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n634), .A2(KEYINPUT99), .A3(new_n636), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n616), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n558), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n465), .B(KEYINPUT100), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(new_n226), .ZN(G1324gat));
  INV_X1    g447(.A(new_n644), .ZN(new_n649));
  INV_X1    g448(.A(new_n550), .ZN(new_n650));
  XOR2_X1   g449(.A(KEYINPUT16), .B(G8gat), .Z(new_n651));
  NAND3_X1  g450(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT42), .ZN(new_n653));
  OR2_X1    g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(G8gat), .B1(new_n644), .B2(new_n550), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n652), .A2(new_n653), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(G1325gat));
  INV_X1    g456(.A(G15gat), .ZN(new_n658));
  NOR3_X1   g457(.A1(new_n644), .A2(new_n658), .A3(new_n545), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n649), .A2(new_n548), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n659), .B1(new_n658), .B2(new_n660), .ZN(G1326gat));
  NOR2_X1   g460(.A1(new_n644), .A2(new_n333), .ZN(new_n662));
  XOR2_X1   g461(.A(KEYINPUT43), .B(G22gat), .Z(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1327gat));
  NAND2_X1  g463(.A1(new_n547), .A2(new_n557), .ZN(new_n665));
  INV_X1    g464(.A(new_n608), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n588), .A2(new_n611), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n667), .A2(new_n641), .A3(new_n261), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n665), .A2(new_n666), .A3(new_n669), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n670), .A2(G29gat), .A3(new_n646), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n671), .B(KEYINPUT45), .Z(new_n672));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n673), .B1(new_n665), .B2(new_n666), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n604), .A2(new_n607), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n601), .A2(new_n602), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n601), .A2(new_n602), .ZN(new_n678));
  AND3_X1   g477(.A1(new_n677), .A2(new_n607), .A3(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n676), .A2(KEYINPUT102), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT102), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(new_n675), .B2(new_n679), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n458), .A2(new_n466), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n499), .B1(new_n685), .B2(new_n540), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n539), .A2(new_n686), .ZN(new_n687));
  AOI211_X1 g486(.A(KEYINPUT44), .B(new_n684), .C1(new_n687), .C2(new_n557), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n674), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n668), .B(KEYINPUT101), .Z(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(G29gat), .B1(new_n691), .B2(new_n646), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n672), .A2(new_n692), .ZN(G1328gat));
  OAI21_X1  g492(.A(G36gat), .B1(new_n691), .B2(new_n550), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n670), .A2(G36gat), .A3(new_n550), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT46), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(G1329gat));
  NAND4_X1  g496(.A1(new_n689), .A2(G43gat), .A3(new_n499), .A4(new_n690), .ZN(new_n698));
  INV_X1    g497(.A(new_n548), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n203), .B1(new_n670), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(KEYINPUT47), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT47), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n698), .A2(new_n703), .A3(new_n700), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(G1330gat));
  NAND4_X1  g504(.A1(new_n689), .A2(G50gat), .A3(new_n540), .A4(new_n690), .ZN(new_n706));
  INV_X1    g505(.A(G50gat), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n707), .B1(new_n670), .B2(new_n333), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(KEYINPUT48), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT48), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n706), .A2(new_n711), .A3(new_n708), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(G1331gat));
  AOI21_X1  g512(.A(new_n261), .B1(new_n687), .B2(new_n557), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n616), .A2(new_n641), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n645), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g518(.A(KEYINPUT49), .B(G64gat), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n717), .A2(new_n650), .A3(new_n720), .ZN(new_n721));
  OAI22_X1  g520(.A1(new_n716), .A2(new_n550), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g522(.A(new_n723), .B(KEYINPUT103), .Z(G1333gat));
  NAND3_X1  g523(.A1(new_n717), .A2(G71gat), .A3(new_n499), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n716), .A2(new_n699), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n725), .B1(G71gat), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g527(.A1(new_n716), .A2(new_n333), .ZN(new_n729));
  XOR2_X1   g528(.A(KEYINPUT104), .B(G78gat), .Z(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(G1335gat));
  NAND2_X1  g530(.A1(new_n667), .A2(new_n262), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n732), .A2(new_n641), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n689), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(G85gat), .B1(new_n734), .B2(new_n646), .ZN(new_n735));
  INV_X1    g534(.A(new_n732), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n543), .A2(new_n545), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n528), .A2(KEYINPUT89), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n537), .A2(new_n530), .A3(new_n525), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n513), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n554), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n742), .A2(new_n458), .A3(new_n466), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n550), .A2(new_n333), .A3(new_n548), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  AOI22_X1  g544(.A1(new_n743), .A2(KEYINPUT35), .B1(new_n745), .B2(new_n552), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n666), .B(new_n736), .C1(new_n741), .C2(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n747), .A2(KEYINPUT105), .A3(KEYINPUT51), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n732), .B1(new_n687), .B2(new_n557), .ZN(new_n749));
  NAND2_X1  g548(.A1(KEYINPUT105), .A2(KEYINPUT51), .ZN(new_n750));
  OR2_X1    g549(.A1(KEYINPUT105), .A2(KEYINPUT51), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n749), .A2(new_n666), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n646), .A2(G85gat), .A3(new_n641), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT106), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n735), .B1(new_n753), .B2(new_n755), .ZN(G1336gat));
  NAND3_X1  g555(.A1(new_n689), .A2(new_n650), .A3(new_n733), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT107), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n550), .A2(new_n641), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n760), .A2(G92gat), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n753), .B1(new_n758), .B2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n761), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT107), .ZN(new_n764));
  AOI22_X1  g563(.A1(G92gat), .A2(new_n757), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n757), .A2(G92gat), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n766), .B1(new_n753), .B2(new_n763), .ZN(new_n768));
  OAI22_X1  g567(.A1(new_n765), .A2(new_n766), .B1(new_n767), .B2(new_n768), .ZN(G1337gat));
  OAI21_X1  g568(.A(G99gat), .B1(new_n734), .B2(new_n545), .ZN(new_n770));
  OR3_X1    g569(.A1(new_n699), .A2(G99gat), .A3(new_n641), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n770), .B1(new_n753), .B2(new_n771), .ZN(G1338gat));
  INV_X1    g571(.A(KEYINPUT110), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT53), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n540), .B(new_n733), .C1(new_n674), .C2(new_n688), .ZN(new_n775));
  XNOR2_X1  g574(.A(KEYINPUT108), .B(G106gat), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n748), .A2(new_n752), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n641), .A2(new_n333), .A3(G106gat), .ZN(new_n779));
  XOR2_X1   g578(.A(new_n779), .B(KEYINPUT109), .Z(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n774), .B1(new_n777), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n748), .A2(new_n752), .A3(new_n779), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n774), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n784), .B1(new_n775), .B2(new_n776), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n773), .B1(new_n782), .B2(new_n785), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n783), .A2(new_n774), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n777), .ZN(new_n788));
  AOI22_X1  g587(.A1(new_n775), .A2(new_n776), .B1(new_n778), .B2(new_n780), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n788), .B(KEYINPUT110), .C1(new_n789), .C2(new_n774), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n786), .A2(new_n790), .ZN(G1339gat));
  INV_X1    g590(.A(new_n667), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n242), .A2(new_n243), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n245), .A2(new_n246), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n256), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n260), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n796), .A2(new_n640), .A3(new_n639), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n635), .B1(new_n624), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n622), .A2(new_n618), .A3(new_n623), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(KEYINPUT54), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n799), .B1(new_n801), .B2(new_n624), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n636), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT111), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n802), .A2(new_n803), .ZN(new_n807));
  OAI211_X1 g606(.A(KEYINPUT111), .B(new_n636), .C1(new_n802), .C2(new_n803), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n797), .B1(new_n809), .B2(new_n262), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n684), .ZN(new_n811));
  INV_X1    g610(.A(new_n809), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n812), .A2(new_n681), .A3(new_n683), .A4(new_n796), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n792), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  AND4_X1   g613(.A1(new_n614), .A2(new_n615), .A3(new_n641), .A4(new_n262), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT112), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT112), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n614), .A2(new_n615), .A3(new_n641), .A4(new_n262), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n681), .A2(new_n683), .A3(new_n796), .ZN(new_n819));
  AOI22_X1  g618(.A1(new_n819), .A2(new_n812), .B1(new_n810), .B2(new_n684), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n817), .B(new_n818), .C1(new_n820), .C2(new_n792), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n816), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n822), .A2(new_n645), .A3(new_n745), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n261), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n825), .A2(KEYINPUT113), .A3(G113gat), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(KEYINPUT113), .B1(new_n825), .B2(G113gat), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n816), .A2(new_n821), .A3(new_n645), .A4(new_n742), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n829), .A2(new_n650), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n261), .A2(new_n348), .ZN(new_n832));
  XOR2_X1   g631(.A(new_n832), .B(KEYINPUT114), .Z(new_n833));
  OAI22_X1  g632(.A1(new_n827), .A2(new_n828), .B1(new_n831), .B2(new_n833), .ZN(G1340gat));
  NAND3_X1  g633(.A1(new_n830), .A2(new_n346), .A3(new_n642), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n824), .A2(new_n642), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n836), .A2(KEYINPUT115), .A3(G120gat), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT115), .B1(new_n836), .B2(G120gat), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n835), .B1(new_n838), .B2(new_n839), .ZN(G1341gat));
  NOR3_X1   g639(.A1(new_n823), .A2(new_n335), .A3(new_n667), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n830), .A2(new_n792), .ZN(new_n842));
  XOR2_X1   g641(.A(new_n842), .B(KEYINPUT116), .Z(new_n843));
  AOI21_X1  g642(.A(new_n841), .B1(new_n843), .B2(new_n335), .ZN(G1342gat));
  NAND3_X1  g643(.A1(new_n830), .A2(new_n336), .A3(new_n666), .ZN(new_n845));
  XNOR2_X1  g644(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n846));
  OR2_X1    g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(G134gat), .B1(new_n823), .B2(new_n608), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n845), .A2(new_n846), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(G1343gat));
  NAND2_X1  g649(.A1(new_n797), .A2(KEYINPUT118), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n802), .A2(new_n803), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n261), .A2(new_n636), .A3(new_n807), .A4(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT118), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n796), .A2(new_n854), .A3(new_n640), .A4(new_n639), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n851), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n608), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n813), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n815), .B1(new_n858), .B2(new_n667), .ZN(new_n859));
  OAI21_X1  g658(.A(KEYINPUT57), .B1(new_n859), .B2(new_n333), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n816), .A2(new_n821), .A3(new_n861), .A4(new_n540), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n645), .A2(new_n550), .A3(new_n545), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n860), .A2(new_n261), .A3(new_n862), .A4(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT120), .B1(new_n865), .B2(new_n280), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(KEYINPUT58), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n822), .A2(new_n540), .A3(new_n864), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n261), .A2(new_n264), .ZN(new_n869));
  XOR2_X1   g668(.A(new_n869), .B(KEYINPUT119), .Z(new_n870));
  NOR2_X1   g669(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n871), .B1(new_n865), .B2(new_n280), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n867), .B(new_n872), .ZN(G1344gat));
  INV_X1    g672(.A(KEYINPUT59), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n816), .A2(new_n540), .A3(new_n821), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(KEYINPUT57), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n809), .A2(new_n608), .ZN(new_n877));
  OR2_X1    g676(.A1(new_n877), .A2(KEYINPUT122), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(KEYINPUT122), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n878), .A2(new_n796), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n792), .B1(new_n880), .B2(new_n857), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n861), .B(new_n540), .C1(new_n881), .C2(new_n815), .ZN(new_n882));
  XOR2_X1   g681(.A(new_n863), .B(KEYINPUT121), .Z(new_n883));
  NAND4_X1  g682(.A1(new_n876), .A2(new_n642), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n884), .A2(KEYINPUT123), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n266), .B1(new_n884), .B2(KEYINPUT123), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n874), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n860), .A2(new_n862), .A3(new_n864), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n874), .B1(new_n888), .B2(new_n641), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n889), .A2(new_n266), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n642), .A2(new_n266), .ZN(new_n891));
  OAI22_X1  g690(.A1(new_n887), .A2(new_n890), .B1(new_n868), .B2(new_n891), .ZN(G1345gat));
  AND2_X1   g691(.A1(new_n860), .A2(new_n864), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n893), .A2(G155gat), .A3(new_n792), .A4(new_n862), .ZN(new_n894));
  INV_X1    g693(.A(G155gat), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n895), .B1(new_n868), .B2(new_n667), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(KEYINPUT124), .ZN(G1346gat));
  OAI21_X1  g697(.A(G162gat), .B1(new_n888), .B2(new_n684), .ZN(new_n899));
  OR2_X1    g698(.A1(new_n868), .A2(G162gat), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(new_n608), .ZN(G1347gat));
  NAND3_X1  g700(.A1(new_n816), .A2(new_n646), .A3(new_n821), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(KEYINPUT125), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT125), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n816), .A2(new_n821), .A3(new_n904), .A4(new_n646), .ZN(new_n905));
  AOI211_X1 g704(.A(new_n554), .B(new_n550), .C1(new_n903), .C2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(G169gat), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n906), .A2(new_n907), .A3(new_n261), .ZN(new_n908));
  AND3_X1   g707(.A1(new_n816), .A2(new_n646), .A3(new_n821), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(new_n549), .A3(new_n650), .ZN(new_n910));
  OAI21_X1  g709(.A(G169gat), .B1(new_n910), .B2(new_n262), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n908), .A2(new_n911), .ZN(G1348gat));
  INV_X1    g711(.A(KEYINPUT126), .ZN(new_n913));
  AOI21_X1  g712(.A(G176gat), .B1(new_n906), .B2(new_n642), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n909), .A2(G176gat), .A3(new_n549), .A4(new_n759), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n913), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n554), .B1(new_n903), .B2(new_n905), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n918), .A2(new_n642), .A3(new_n650), .ZN(new_n919));
  INV_X1    g718(.A(G176gat), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n921), .A2(KEYINPUT126), .A3(new_n915), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n917), .A2(new_n922), .ZN(G1349gat));
  NAND4_X1  g722(.A1(new_n918), .A2(new_n792), .A3(new_n404), .A4(new_n650), .ZN(new_n924));
  OAI21_X1  g723(.A(G183gat), .B1(new_n910), .B2(new_n667), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(KEYINPUT60), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT60), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n924), .A2(new_n928), .A3(new_n925), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(G1350gat));
  INV_X1    g729(.A(new_n684), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n906), .A2(new_n398), .A3(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(new_n910), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n398), .B1(new_n933), .B2(new_n666), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT61), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n934), .A2(new_n935), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n932), .B1(new_n936), .B2(new_n937), .ZN(G1351gat));
  AND2_X1   g737(.A1(new_n876), .A2(new_n882), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n499), .A2(new_n550), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n941), .A2(new_n645), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g742(.A(G197gat), .B1(new_n943), .B2(new_n262), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n941), .B1(new_n903), .B2(new_n905), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n945), .A2(new_n253), .A3(new_n540), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n944), .B1(new_n262), .B2(new_n946), .ZN(G1352gat));
  INV_X1    g746(.A(G204gat), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n945), .A2(new_n948), .A3(new_n642), .A4(new_n540), .ZN(new_n949));
  XNOR2_X1  g748(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n950));
  OR2_X1    g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n950), .ZN(new_n952));
  AND3_X1   g751(.A1(new_n939), .A2(new_n642), .A3(new_n942), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n951), .B(new_n952), .C1(new_n948), .C2(new_n953), .ZN(G1353gat));
  NAND4_X1  g753(.A1(new_n945), .A2(new_n287), .A3(new_n792), .A4(new_n540), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n939), .A2(new_n792), .A3(new_n942), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n956), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT63), .B1(new_n956), .B2(G211gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(G1354gat));
  NOR3_X1   g758(.A1(new_n943), .A2(new_n288), .A3(new_n608), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n945), .A2(new_n540), .A3(new_n931), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n960), .B1(new_n961), .B2(new_n288), .ZN(G1355gat));
endmodule


