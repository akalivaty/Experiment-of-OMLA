

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590;

  XNOR2_X1 U325 ( .A(n451), .B(KEYINPUT113), .ZN(n549) );
  XNOR2_X1 U326 ( .A(KEYINPUT96), .B(KEYINPUT26), .ZN(n471) );
  XOR2_X1 U327 ( .A(n390), .B(n389), .Z(n517) );
  XNOR2_X1 U328 ( .A(KEYINPUT37), .B(KEYINPUT103), .ZN(n488) );
  XOR2_X1 U329 ( .A(KEYINPUT110), .B(n393), .Z(n293) );
  XNOR2_X1 U330 ( .A(n472), .B(n471), .ZN(n553) );
  INV_X1 U331 ( .A(KEYINPUT83), .ZN(n341) );
  XNOR2_X1 U332 ( .A(n382), .B(KEYINPUT68), .ZN(n383) );
  XNOR2_X1 U333 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U334 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U335 ( .A(n384), .B(n383), .ZN(n388) );
  XNOR2_X1 U336 ( .A(n344), .B(n343), .ZN(n440) );
  XNOR2_X1 U337 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U338 ( .A(n489), .B(n488), .ZN(n531) );
  NOR2_X1 U339 ( .A1(n483), .A2(n482), .ZN(n498) );
  AND2_X1 U340 ( .A1(n450), .A2(n540), .ZN(n451) );
  INV_X1 U341 ( .A(G190GAT), .ZN(n468) );
  INV_X1 U342 ( .A(G127GAT), .ZN(n452) );
  XNOR2_X1 U343 ( .A(n468), .B(KEYINPUT58), .ZN(n469) );
  XNOR2_X1 U344 ( .A(n452), .B(KEYINPUT50), .ZN(n453) );
  XNOR2_X1 U345 ( .A(n492), .B(G43GAT), .ZN(n493) );
  XNOR2_X1 U346 ( .A(n470), .B(n469), .ZN(G1351GAT) );
  XNOR2_X1 U347 ( .A(n494), .B(n493), .ZN(G1330GAT) );
  XOR2_X1 U348 ( .A(KEYINPUT79), .B(KEYINPUT12), .Z(n295) );
  XNOR2_X1 U349 ( .A(KEYINPUT78), .B(KEYINPUT14), .ZN(n294) );
  XNOR2_X1 U350 ( .A(n295), .B(n294), .ZN(n313) );
  XOR2_X1 U351 ( .A(KEYINPUT80), .B(KEYINPUT81), .Z(n297) );
  XNOR2_X1 U352 ( .A(G22GAT), .B(G64GAT), .ZN(n296) );
  XNOR2_X1 U353 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U354 ( .A(G211GAT), .B(G78GAT), .Z(n299) );
  XNOR2_X1 U355 ( .A(G71GAT), .B(G155GAT), .ZN(n298) );
  XNOR2_X1 U356 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U357 ( .A(n301), .B(n300), .ZN(n311) );
  XNOR2_X1 U358 ( .A(G8GAT), .B(G183GAT), .ZN(n302) );
  XNOR2_X1 U359 ( .A(n302), .B(KEYINPUT77), .ZN(n327) );
  XOR2_X1 U360 ( .A(KEYINPUT15), .B(n327), .Z(n304) );
  NAND2_X1 U361 ( .A1(G231GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U362 ( .A(n304), .B(n303), .ZN(n307) );
  XOR2_X1 U363 ( .A(KEYINPUT13), .B(KEYINPUT69), .Z(n306) );
  XNOR2_X1 U364 ( .A(G57GAT), .B(KEYINPUT70), .ZN(n305) );
  XNOR2_X1 U365 ( .A(n306), .B(n305), .ZN(n362) );
  XOR2_X1 U366 ( .A(n307), .B(n362), .Z(n309) );
  XOR2_X1 U367 ( .A(G1GAT), .B(KEYINPUT67), .Z(n377) );
  XOR2_X1 U368 ( .A(G15GAT), .B(G127GAT), .Z(n435) );
  XNOR2_X1 U369 ( .A(n377), .B(n435), .ZN(n308) );
  XNOR2_X1 U370 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U371 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U372 ( .A(n313), .B(n312), .Z(n582) );
  XOR2_X1 U373 ( .A(KEYINPUT19), .B(KEYINPUT86), .Z(n315) );
  XNOR2_X1 U374 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n314) );
  XNOR2_X1 U375 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U376 ( .A(G169GAT), .B(n316), .Z(n447) );
  XOR2_X1 U377 ( .A(G64GAT), .B(KEYINPUT73), .Z(n318) );
  XNOR2_X1 U378 ( .A(G176GAT), .B(G204GAT), .ZN(n317) );
  XNOR2_X1 U379 ( .A(n318), .B(n317), .ZN(n363) );
  XOR2_X1 U380 ( .A(G36GAT), .B(G190GAT), .Z(n396) );
  XOR2_X1 U381 ( .A(n363), .B(n396), .Z(n320) );
  NAND2_X1 U382 ( .A1(G226GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U383 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U384 ( .A(KEYINPUT91), .B(KEYINPUT93), .Z(n322) );
  XNOR2_X1 U385 ( .A(G92GAT), .B(KEYINPUT92), .ZN(n321) );
  XNOR2_X1 U386 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U387 ( .A(n324), .B(n323), .Z(n329) );
  XOR2_X1 U388 ( .A(G211GAT), .B(KEYINPUT21), .Z(n326) );
  XNOR2_X1 U389 ( .A(G197GAT), .B(G218GAT), .ZN(n325) );
  XNOR2_X1 U390 ( .A(n326), .B(n325), .ZN(n420) );
  XNOR2_X1 U391 ( .A(n420), .B(n327), .ZN(n328) );
  XNOR2_X1 U392 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U393 ( .A(n447), .B(n330), .Z(n523) );
  XOR2_X1 U394 ( .A(KEYINPUT27), .B(KEYINPUT94), .Z(n331) );
  XOR2_X1 U395 ( .A(n523), .B(n331), .Z(n473) );
  XOR2_X1 U396 ( .A(G155GAT), .B(KEYINPUT3), .Z(n333) );
  XNOR2_X1 U397 ( .A(KEYINPUT2), .B(KEYINPUT88), .ZN(n332) );
  XNOR2_X1 U398 ( .A(n333), .B(n332), .ZN(n432) );
  XOR2_X1 U399 ( .A(G85GAT), .B(n432), .Z(n335) );
  NAND2_X1 U400 ( .A1(G225GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U401 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U402 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n337) );
  XNOR2_X1 U403 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n336) );
  XNOR2_X1 U404 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U405 ( .A(n339), .B(n338), .Z(n346) );
  XNOR2_X1 U406 ( .A(KEYINPUT0), .B(KEYINPUT82), .ZN(n340) );
  XNOR2_X1 U407 ( .A(n340), .B(KEYINPUT84), .ZN(n344) );
  XNOR2_X1 U408 ( .A(G113GAT), .B(G134GAT), .ZN(n342) );
  XNOR2_X1 U409 ( .A(G29GAT), .B(n440), .ZN(n345) );
  XNOR2_X1 U410 ( .A(n346), .B(n345), .ZN(n354) );
  XOR2_X1 U411 ( .A(KEYINPUT6), .B(KEYINPUT90), .Z(n348) );
  XNOR2_X1 U412 ( .A(G141GAT), .B(G57GAT), .ZN(n347) );
  XNOR2_X1 U413 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U414 ( .A(G162GAT), .B(G148GAT), .Z(n350) );
  XNOR2_X1 U415 ( .A(G120GAT), .B(G127GAT), .ZN(n349) );
  XNOR2_X1 U416 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U417 ( .A(n352), .B(n351), .Z(n353) );
  XOR2_X1 U418 ( .A(n354), .B(n353), .Z(n534) );
  INV_X1 U419 ( .A(n534), .ZN(n519) );
  NOR2_X1 U420 ( .A1(n473), .A2(n519), .ZN(n355) );
  XOR2_X1 U421 ( .A(KEYINPUT95), .B(n355), .Z(n480) );
  XNOR2_X1 U422 ( .A(G106GAT), .B(G78GAT), .ZN(n356) );
  XNOR2_X1 U423 ( .A(n356), .B(G148GAT), .ZN(n431) );
  XOR2_X1 U424 ( .A(KEYINPUT71), .B(G92GAT), .Z(n358) );
  XNOR2_X1 U425 ( .A(G99GAT), .B(G85GAT), .ZN(n357) );
  XNOR2_X1 U426 ( .A(n358), .B(n357), .ZN(n397) );
  XOR2_X1 U427 ( .A(n431), .B(n397), .Z(n371) );
  XOR2_X1 U428 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n360) );
  NAND2_X1 U429 ( .A1(G230GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U430 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U431 ( .A(n361), .B(KEYINPUT33), .Z(n365) );
  XNOR2_X1 U432 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U433 ( .A(n365), .B(n364), .ZN(n369) );
  XOR2_X1 U434 ( .A(G120GAT), .B(G71GAT), .Z(n436) );
  XNOR2_X1 U435 ( .A(n436), .B(KEYINPUT72), .ZN(n367) );
  INV_X1 U436 ( .A(KEYINPUT74), .ZN(n366) );
  XNOR2_X1 U437 ( .A(n371), .B(n370), .ZN(n578) );
  XOR2_X1 U438 ( .A(n578), .B(KEYINPUT64), .Z(n372) );
  XNOR2_X1 U439 ( .A(n372), .B(KEYINPUT41), .ZN(n566) );
  XOR2_X1 U440 ( .A(G197GAT), .B(G113GAT), .Z(n374) );
  XNOR2_X1 U441 ( .A(G169GAT), .B(G15GAT), .ZN(n373) );
  XNOR2_X1 U442 ( .A(n374), .B(n373), .ZN(n390) );
  XOR2_X1 U443 ( .A(KEYINPUT66), .B(KEYINPUT65), .Z(n376) );
  XNOR2_X1 U444 ( .A(G8GAT), .B(KEYINPUT30), .ZN(n375) );
  XNOR2_X1 U445 ( .A(n376), .B(n375), .ZN(n381) );
  XOR2_X1 U446 ( .A(G50GAT), .B(G36GAT), .Z(n378) );
  XNOR2_X1 U447 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U448 ( .A(G141GAT), .B(G22GAT), .Z(n424) );
  XNOR2_X1 U449 ( .A(n379), .B(n424), .ZN(n380) );
  XOR2_X1 U450 ( .A(n381), .B(n380), .Z(n384) );
  NAND2_X1 U451 ( .A1(G229GAT), .A2(G233GAT), .ZN(n382) );
  XOR2_X1 U452 ( .A(G29GAT), .B(G43GAT), .Z(n386) );
  XNOR2_X1 U453 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n385) );
  XNOR2_X1 U454 ( .A(n386), .B(n385), .ZN(n401) );
  XOR2_X1 U455 ( .A(n401), .B(KEYINPUT29), .Z(n387) );
  XNOR2_X1 U456 ( .A(n388), .B(n387), .ZN(n389) );
  INV_X1 U457 ( .A(n517), .ZN(n573) );
  NOR2_X1 U458 ( .A1(n566), .A2(n573), .ZN(n391) );
  XNOR2_X1 U459 ( .A(n391), .B(KEYINPUT46), .ZN(n392) );
  INV_X1 U460 ( .A(n582), .ZN(n484) );
  NOR2_X1 U461 ( .A1(n392), .A2(n484), .ZN(n393) );
  XOR2_X1 U462 ( .A(KEYINPUT75), .B(KEYINPUT10), .Z(n395) );
  XNOR2_X1 U463 ( .A(G106GAT), .B(KEYINPUT11), .ZN(n394) );
  XNOR2_X1 U464 ( .A(n395), .B(n394), .ZN(n408) );
  XOR2_X1 U465 ( .A(n397), .B(n396), .Z(n399) );
  NAND2_X1 U466 ( .A1(G232GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U467 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U468 ( .A(n400), .B(KEYINPUT76), .Z(n403) );
  XNOR2_X1 U469 ( .A(n401), .B(KEYINPUT9), .ZN(n402) );
  XNOR2_X1 U470 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U471 ( .A(n404), .B(G218GAT), .Z(n406) );
  XOR2_X1 U472 ( .A(G50GAT), .B(G162GAT), .Z(n419) );
  XNOR2_X1 U473 ( .A(G134GAT), .B(n419), .ZN(n405) );
  XNOR2_X1 U474 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U475 ( .A(n408), .B(n407), .ZN(n495) );
  NOR2_X1 U476 ( .A1(n293), .A2(n495), .ZN(n409) );
  XNOR2_X1 U477 ( .A(n409), .B(KEYINPUT47), .ZN(n416) );
  XNOR2_X1 U478 ( .A(KEYINPUT36), .B(KEYINPUT101), .ZN(n410) );
  XNOR2_X1 U479 ( .A(n495), .B(n410), .ZN(n587) );
  NOR2_X1 U480 ( .A1(n582), .A2(n587), .ZN(n411) );
  XNOR2_X1 U481 ( .A(n411), .B(KEYINPUT45), .ZN(n412) );
  NAND2_X1 U482 ( .A1(n412), .A2(n578), .ZN(n413) );
  XNOR2_X1 U483 ( .A(n413), .B(KEYINPUT111), .ZN(n414) );
  NAND2_X1 U484 ( .A1(n414), .A2(n573), .ZN(n415) );
  NAND2_X1 U485 ( .A1(n416), .A2(n415), .ZN(n417) );
  XNOR2_X1 U486 ( .A(n417), .B(KEYINPUT48), .ZN(n455) );
  NAND2_X1 U487 ( .A1(n480), .A2(n455), .ZN(n418) );
  XNOR2_X1 U488 ( .A(n418), .B(KEYINPUT112), .ZN(n554) );
  XOR2_X1 U489 ( .A(n420), .B(n419), .Z(n422) );
  NAND2_X1 U490 ( .A1(G228GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U491 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U492 ( .A(n423), .B(G204GAT), .Z(n426) );
  XNOR2_X1 U493 ( .A(n424), .B(KEYINPUT24), .ZN(n425) );
  XNOR2_X1 U494 ( .A(n426), .B(n425), .ZN(n430) );
  XOR2_X1 U495 ( .A(KEYINPUT89), .B(KEYINPUT87), .Z(n428) );
  XNOR2_X1 U496 ( .A(KEYINPUT22), .B(KEYINPUT23), .ZN(n427) );
  XNOR2_X1 U497 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U498 ( .A(n430), .B(n429), .Z(n434) );
  XNOR2_X1 U499 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U500 ( .A(n434), .B(n433), .ZN(n475) );
  XOR2_X1 U501 ( .A(n475), .B(KEYINPUT28), .Z(n528) );
  INV_X1 U502 ( .A(n528), .ZN(n543) );
  NOR2_X1 U503 ( .A1(n554), .A2(n543), .ZN(n450) );
  XOR2_X1 U504 ( .A(G183GAT), .B(G190GAT), .Z(n438) );
  XNOR2_X1 U505 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U506 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U507 ( .A(n439), .B(G99GAT), .Z(n442) );
  XNOR2_X1 U508 ( .A(G43GAT), .B(n440), .ZN(n441) );
  XNOR2_X1 U509 ( .A(n442), .B(n441), .ZN(n446) );
  XOR2_X1 U510 ( .A(KEYINPUT20), .B(KEYINPUT85), .Z(n444) );
  NAND2_X1 U511 ( .A1(G227GAT), .A2(G233GAT), .ZN(n443) );
  XOR2_X1 U512 ( .A(n444), .B(n443), .Z(n445) );
  XNOR2_X1 U513 ( .A(n446), .B(n445), .ZN(n449) );
  XNOR2_X1 U514 ( .A(n447), .B(G176GAT), .ZN(n448) );
  XOR2_X1 U515 ( .A(n449), .B(n448), .Z(n525) );
  INV_X1 U516 ( .A(n525), .ZN(n540) );
  NOR2_X1 U517 ( .A1(n582), .A2(n549), .ZN(n454) );
  XNOR2_X1 U518 ( .A(n454), .B(n453), .ZN(G1342GAT) );
  INV_X1 U519 ( .A(n523), .ZN(n537) );
  NAND2_X1 U520 ( .A1(n455), .A2(n537), .ZN(n457) );
  XOR2_X1 U521 ( .A(KEYINPUT118), .B(KEYINPUT54), .Z(n456) );
  XNOR2_X1 U522 ( .A(n457), .B(n456), .ZN(n458) );
  NAND2_X1 U523 ( .A1(n458), .A2(n519), .ZN(n572) );
  NOR2_X1 U524 ( .A1(n475), .A2(n572), .ZN(n460) );
  XNOR2_X1 U525 ( .A(KEYINPUT119), .B(KEYINPUT55), .ZN(n459) );
  XNOR2_X1 U526 ( .A(n460), .B(n459), .ZN(n461) );
  NAND2_X1 U527 ( .A1(n461), .A2(n540), .ZN(n567) );
  NOR2_X1 U528 ( .A1(n573), .A2(n567), .ZN(n464) );
  INV_X1 U529 ( .A(G169GAT), .ZN(n462) );
  XNOR2_X1 U530 ( .A(n462), .B(KEYINPUT120), .ZN(n463) );
  XNOR2_X1 U531 ( .A(n464), .B(n463), .ZN(G1348GAT) );
  NOR2_X1 U532 ( .A1(n582), .A2(n567), .ZN(n467) );
  INV_X1 U533 ( .A(G183GAT), .ZN(n465) );
  XNOR2_X1 U534 ( .A(n465), .B(KEYINPUT122), .ZN(n466) );
  XNOR2_X1 U535 ( .A(n467), .B(n466), .ZN(G1350GAT) );
  INV_X1 U536 ( .A(n495), .ZN(n564) );
  NOR2_X1 U537 ( .A1(n564), .A2(n567), .ZN(n470) );
  AND2_X1 U538 ( .A1(n578), .A2(n517), .ZN(n499) );
  INV_X1 U539 ( .A(KEYINPUT102), .ZN(n486) );
  NAND2_X1 U540 ( .A1(n525), .A2(n475), .ZN(n472) );
  NOR2_X1 U541 ( .A1(n553), .A2(n473), .ZN(n478) );
  NOR2_X1 U542 ( .A1(n523), .A2(n525), .ZN(n474) );
  NOR2_X1 U543 ( .A1(n475), .A2(n474), .ZN(n476) );
  XOR2_X1 U544 ( .A(KEYINPUT25), .B(n476), .Z(n477) );
  NOR2_X1 U545 ( .A1(n478), .A2(n477), .ZN(n479) );
  NOR2_X1 U546 ( .A1(n479), .A2(n534), .ZN(n483) );
  NAND2_X1 U547 ( .A1(n480), .A2(n525), .ZN(n481) );
  NOR2_X1 U548 ( .A1(n481), .A2(n543), .ZN(n482) );
  NOR2_X1 U549 ( .A1(n498), .A2(n484), .ZN(n485) );
  XNOR2_X1 U550 ( .A(n486), .B(n485), .ZN(n487) );
  NOR2_X1 U551 ( .A1(n587), .A2(n487), .ZN(n489) );
  NAND2_X1 U552 ( .A1(n499), .A2(n531), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n490), .B(KEYINPUT38), .ZN(n491) );
  XNOR2_X1 U554 ( .A(KEYINPUT104), .B(n491), .ZN(n514) );
  NOR2_X1 U555 ( .A1(n525), .A2(n514), .ZN(n494) );
  INV_X1 U556 ( .A(KEYINPUT40), .ZN(n492) );
  NOR2_X1 U557 ( .A1(n582), .A2(n495), .ZN(n496) );
  XOR2_X1 U558 ( .A(KEYINPUT16), .B(n496), .Z(n497) );
  NOR2_X1 U559 ( .A1(n498), .A2(n497), .ZN(n518) );
  NAND2_X1 U560 ( .A1(n499), .A2(n518), .ZN(n500) );
  XNOR2_X1 U561 ( .A(KEYINPUT97), .B(n500), .ZN(n508) );
  NAND2_X1 U562 ( .A1(n508), .A2(n534), .ZN(n504) );
  XOR2_X1 U563 ( .A(KEYINPUT99), .B(KEYINPUT34), .Z(n502) );
  XNOR2_X1 U564 ( .A(G1GAT), .B(KEYINPUT98), .ZN(n501) );
  XNOR2_X1 U565 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U566 ( .A(n504), .B(n503), .ZN(G1324GAT) );
  NAND2_X1 U567 ( .A1(n537), .A2(n508), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n505), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U569 ( .A(G15GAT), .B(KEYINPUT35), .Z(n507) );
  NAND2_X1 U570 ( .A1(n508), .A2(n540), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(G1326GAT) );
  NAND2_X1 U572 ( .A1(n543), .A2(n508), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n509), .B(KEYINPUT100), .ZN(n510) );
  XNOR2_X1 U574 ( .A(G22GAT), .B(n510), .ZN(G1327GAT) );
  NOR2_X1 U575 ( .A1(n519), .A2(n514), .ZN(n512) );
  XNOR2_X1 U576 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n512), .B(n511), .ZN(G1328GAT) );
  NOR2_X1 U578 ( .A1(n523), .A2(n514), .ZN(n513) );
  XOR2_X1 U579 ( .A(G36GAT), .B(n513), .Z(G1329GAT) );
  NOR2_X1 U580 ( .A1(n528), .A2(n514), .ZN(n516) );
  XNOR2_X1 U581 ( .A(G50GAT), .B(KEYINPUT105), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n516), .B(n515), .ZN(G1331GAT) );
  NOR2_X1 U583 ( .A1(n517), .A2(n566), .ZN(n532) );
  NAND2_X1 U584 ( .A1(n532), .A2(n518), .ZN(n527) );
  NOR2_X1 U585 ( .A1(n519), .A2(n527), .ZN(n521) );
  XNOR2_X1 U586 ( .A(KEYINPUT106), .B(KEYINPUT42), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U588 ( .A(G57GAT), .B(n522), .Z(G1332GAT) );
  NOR2_X1 U589 ( .A1(n523), .A2(n527), .ZN(n524) );
  XOR2_X1 U590 ( .A(G64GAT), .B(n524), .Z(G1333GAT) );
  NOR2_X1 U591 ( .A1(n525), .A2(n527), .ZN(n526) );
  XOR2_X1 U592 ( .A(G71GAT), .B(n526), .Z(G1334GAT) );
  NOR2_X1 U593 ( .A1(n528), .A2(n527), .ZN(n530) );
  XNOR2_X1 U594 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n529) );
  XNOR2_X1 U595 ( .A(n530), .B(n529), .ZN(G1335GAT) );
  NAND2_X1 U596 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U597 ( .A(n533), .B(KEYINPUT107), .ZN(n542) );
  NAND2_X1 U598 ( .A1(n542), .A2(n534), .ZN(n535) );
  XNOR2_X1 U599 ( .A(n535), .B(KEYINPUT108), .ZN(n536) );
  XNOR2_X1 U600 ( .A(G85GAT), .B(n536), .ZN(G1336GAT) );
  XOR2_X1 U601 ( .A(G92GAT), .B(KEYINPUT109), .Z(n539) );
  NAND2_X1 U602 ( .A1(n542), .A2(n537), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(G1337GAT) );
  NAND2_X1 U604 ( .A1(n542), .A2(n540), .ZN(n541) );
  XNOR2_X1 U605 ( .A(n541), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U606 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U607 ( .A(n544), .B(KEYINPUT44), .ZN(n545) );
  XNOR2_X1 U608 ( .A(G106GAT), .B(n545), .ZN(G1339GAT) );
  NOR2_X1 U609 ( .A1(n573), .A2(n549), .ZN(n546) );
  XOR2_X1 U610 ( .A(G113GAT), .B(n546), .Z(G1340GAT) );
  NOR2_X1 U611 ( .A1(n566), .A2(n549), .ZN(n548) );
  XNOR2_X1 U612 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(G1341GAT) );
  NOR2_X1 U614 ( .A1(n564), .A2(n549), .ZN(n551) );
  XNOR2_X1 U615 ( .A(KEYINPUT114), .B(KEYINPUT51), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U617 ( .A(G134GAT), .B(n552), .ZN(G1343GAT) );
  NOR2_X1 U618 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U619 ( .A(KEYINPUT115), .B(n555), .ZN(n563) );
  NOR2_X1 U620 ( .A1(n573), .A2(n563), .ZN(n556) );
  XOR2_X1 U621 ( .A(G141GAT), .B(n556), .Z(n557) );
  XNOR2_X1 U622 ( .A(KEYINPUT116), .B(n557), .ZN(G1344GAT) );
  NOR2_X1 U623 ( .A1(n563), .A2(n566), .ZN(n561) );
  XOR2_X1 U624 ( .A(KEYINPUT117), .B(KEYINPUT52), .Z(n559) );
  XNOR2_X1 U625 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(G1345GAT) );
  NOR2_X1 U628 ( .A1(n582), .A2(n563), .ZN(n562) );
  XOR2_X1 U629 ( .A(G155GAT), .B(n562), .Z(G1346GAT) );
  NOR2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U631 ( .A(G162GAT), .B(n565), .Z(G1347GAT) );
  NOR2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n571) );
  XOR2_X1 U633 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n569) );
  XNOR2_X1 U634 ( .A(G176GAT), .B(KEYINPUT121), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1349GAT) );
  OR2_X1 U637 ( .A1(n572), .A2(n553), .ZN(n586) );
  NOR2_X1 U638 ( .A1(n586), .A2(n573), .ZN(n577) );
  XOR2_X1 U639 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n575) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  NOR2_X1 U643 ( .A1(n578), .A2(n586), .ZN(n580) );
  XNOR2_X1 U644 ( .A(KEYINPUT124), .B(KEYINPUT61), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(n581), .ZN(G1353GAT) );
  NOR2_X1 U647 ( .A1(n582), .A2(n586), .ZN(n584) );
  XNOR2_X1 U648 ( .A(KEYINPUT125), .B(KEYINPUT126), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(G211GAT), .B(n585), .ZN(G1354GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n589) );
  XNOR2_X1 U652 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

