//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 0 0 1 0 0 1 0 0 0 1 1 1 1 0 1 0 0 0 1 0 0 1 1 0 1 0 0 0 1 1 1 0 0 0 1 0 1 1 0 0 1 0 1 0 0 1 1 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n811, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n960, new_n961, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1018, new_n1019, new_n1020,
    new_n1021;
  XOR2_X1   g000(.A(G78gat), .B(G106gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT81), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT31), .B(G50gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(KEYINPUT82), .ZN(new_n206));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT2), .ZN(new_n208));
  INV_X1    g007(.A(G148gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n209), .A2(G141gat), .ZN(new_n210));
  INV_X1    g009(.A(G141gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n211), .A2(G148gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n208), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  AND2_X1   g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215));
  NOR3_X1   g014(.A1(new_n214), .A2(new_n215), .A3(KEYINPUT77), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT77), .ZN(new_n217));
  INV_X1    g016(.A(G155gat), .ZN(new_n218));
  INV_X1    g017(.A(G162gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n217), .B1(new_n220), .B2(new_n207), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n213), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT78), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(new_n209), .B2(G141gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n209), .A2(G141gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n211), .A2(KEYINPUT78), .A3(G148gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n207), .B1(new_n220), .B2(KEYINPUT2), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n222), .A2(new_n223), .A3(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT79), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT77), .B1(new_n214), .B2(new_n215), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n220), .A2(new_n217), .A3(new_n207), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  AOI22_X1  g035(.A1(new_n236), .A2(new_n213), .B1(new_n228), .B2(new_n229), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n237), .A2(KEYINPUT79), .A3(new_n223), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT29), .B1(new_n233), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT22), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT73), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT73), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT22), .ZN(new_n243));
  NAND2_X1  g042(.A1(G211gat), .A2(G218gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n241), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT74), .ZN(new_n246));
  XOR2_X1   g045(.A(G197gat), .B(G204gat), .Z(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT74), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n241), .A2(new_n243), .A3(new_n249), .A4(new_n244), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n246), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  XOR2_X1   g050(.A(G211gat), .B(G218gat), .Z(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n247), .B1(new_n245), .B2(KEYINPUT74), .ZN(new_n254));
  INV_X1    g053(.A(new_n252), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n254), .A2(new_n255), .A3(new_n250), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n206), .B1(new_n239), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT29), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT79), .B1(new_n237), .B2(new_n223), .ZN(new_n260));
  AND4_X1   g059(.A1(KEYINPUT79), .A2(new_n222), .A3(new_n223), .A4(new_n230), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n257), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n262), .A2(KEYINPUT82), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n222), .A2(new_n230), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT29), .B1(new_n253), .B2(new_n256), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n265), .B1(new_n266), .B2(KEYINPUT3), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n258), .A2(new_n264), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G228gat), .A2(G233gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G22gat), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT83), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n262), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n239), .A2(KEYINPUT83), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n273), .A2(new_n274), .A3(new_n263), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n251), .A2(new_n252), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n255), .B1(new_n254), .B2(new_n250), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n259), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n237), .B1(new_n278), .B2(new_n223), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n279), .A2(new_n269), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n275), .A2(new_n280), .ZN(new_n281));
  AND3_X1   g080(.A1(new_n270), .A2(new_n271), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n271), .B1(new_n270), .B2(new_n281), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n205), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT84), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI211_X1 g085(.A(KEYINPUT84), .B(new_n205), .C1(new_n282), .C2(new_n283), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n283), .A2(KEYINPUT85), .ZN(new_n288));
  AOI22_X1  g087(.A1(new_n268), .A2(new_n269), .B1(new_n275), .B2(new_n280), .ZN(new_n289));
  NAND2_X1  g088(.A1(KEYINPUT85), .A2(G22gat), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n205), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n286), .A2(new_n287), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n294));
  INV_X1    g093(.A(G227gat), .ZN(new_n295));
  INV_X1    g094(.A(G233gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G113gat), .ZN(new_n298));
  INV_X1    g097(.A(G120gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G113gat), .A2(G120gat), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT68), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G127gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G134gat), .ZN(new_n304));
  INV_X1    g103(.A(G134gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G127gat), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT1), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n304), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n302), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n300), .A2(KEYINPUT68), .A3(new_n301), .ZN(new_n310));
  AND2_X1   g109(.A1(G113gat), .A2(G120gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(G113gat), .A2(G120gat), .ZN(new_n312));
  NOR3_X1   g111(.A1(new_n311), .A2(new_n312), .A3(KEYINPUT1), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n305), .A2(KEYINPUT67), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT67), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(G134gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n315), .A2(new_n317), .A3(G127gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(new_n304), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n309), .A2(new_n310), .B1(new_n314), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT23), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n321), .B1(G169gat), .B2(G176gat), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n322), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(G183gat), .A2(G190gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n322), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(G169gat), .ZN(new_n328));
  INV_X1    g127(.A(G176gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(new_n329), .A3(KEYINPUT23), .ZN(new_n330));
  NAND2_X1  g129(.A1(G169gat), .A2(G176gat), .ZN(new_n331));
  AND2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT25), .B1(new_n327), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n328), .A2(new_n329), .A3(KEYINPUT64), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT64), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n335), .B1(G169gat), .B2(G176gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(new_n336), .A3(KEYINPUT23), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(new_n331), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT65), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n337), .A2(KEYINPUT65), .A3(new_n331), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT25), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n343), .B1(new_n323), .B2(new_n326), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n333), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(G183gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT27), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT27), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(G183gat), .ZN(new_n349));
  INV_X1    g148(.A(G190gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n347), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT28), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n352), .A2(KEYINPUT66), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n351), .A2(new_n353), .B1(G183gat), .B2(G190gat), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT26), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n334), .A2(new_n336), .A3(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n356), .A2(new_n331), .A3(new_n357), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n347), .A2(new_n349), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n359), .A2(new_n360), .A3(new_n350), .ZN(new_n361));
  AND3_X1   g160(.A1(new_n354), .A2(new_n358), .A3(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n320), .B1(new_n345), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n333), .ZN(new_n364));
  AND3_X1   g163(.A1(new_n337), .A2(KEYINPUT65), .A3(new_n331), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT65), .B1(new_n337), .B2(new_n331), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n344), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n307), .B1(new_n305), .B2(G127gat), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n303), .A2(G134gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT68), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n372), .B1(new_n311), .B2(new_n312), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n371), .A2(new_n310), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n304), .ZN(new_n375));
  XNOR2_X1  g174(.A(KEYINPUT67), .B(G134gat), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n375), .B1(new_n376), .B2(G127gat), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n374), .B1(new_n377), .B2(new_n313), .ZN(new_n378));
  INV_X1    g177(.A(new_n362), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n368), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n297), .B1(new_n363), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT34), .ZN(new_n382));
  AND2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n381), .A2(new_n382), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n363), .A2(new_n297), .A3(new_n380), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT33), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(KEYINPUT32), .ZN(new_n389));
  XNOR2_X1  g188(.A(G15gat), .B(G43gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n390), .B(KEYINPUT69), .ZN(new_n391));
  XNOR2_X1  g190(.A(G71gat), .B(G99gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n391), .B(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n388), .A2(new_n389), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT70), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT70), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n388), .A2(new_n389), .A3(new_n396), .A4(new_n393), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n393), .A2(KEYINPUT33), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n386), .A2(KEYINPUT32), .A3(new_n398), .ZN(new_n399));
  AND4_X1   g198(.A1(new_n385), .A2(new_n395), .A3(new_n397), .A4(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n399), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n401), .B1(new_n394), .B2(KEYINPUT70), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n385), .B1(new_n402), .B2(new_n397), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n294), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n395), .A2(new_n385), .A3(new_n397), .A4(new_n399), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT72), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT5), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n265), .A2(new_n378), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n314), .A2(new_n319), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n409), .A2(new_n222), .A3(new_n230), .A4(new_n374), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(G225gat), .A2(G233gat), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n407), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT4), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n410), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n320), .A2(KEYINPUT4), .A3(new_n237), .ZN(new_n418));
  AND2_X1   g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n265), .A2(KEYINPUT3), .B1(new_n409), .B2(new_n374), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n420), .B1(new_n260), .B2(new_n261), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n415), .B1(new_n422), .B2(new_n413), .ZN(new_n423));
  XNOR2_X1  g222(.A(G1gat), .B(G29gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n424), .B(KEYINPUT0), .ZN(new_n425));
  XNOR2_X1  g224(.A(G57gat), .B(G85gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n419), .A2(new_n421), .A3(KEYINPUT5), .A4(new_n412), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n423), .A2(KEYINPUT6), .A3(new_n427), .A4(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n378), .B1(new_n237), .B2(new_n223), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n430), .B1(new_n233), .B2(new_n238), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n417), .A2(new_n418), .ZN(new_n432));
  NOR3_X1   g231(.A1(new_n431), .A2(new_n432), .A3(new_n413), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n427), .B(new_n428), .C1(new_n433), .C2(new_n414), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT6), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n427), .B1(new_n423), .B2(new_n428), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n429), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT35), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT75), .ZN(new_n441));
  NAND2_X1  g240(.A1(G226gat), .A2(G233gat), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n362), .B1(new_n364), .B2(new_n367), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n442), .B1(new_n443), .B2(KEYINPUT29), .ZN(new_n444));
  OAI211_X1 g243(.A(G226gat), .B(G233gat), .C1(new_n345), .C2(new_n362), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n444), .A2(new_n257), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n257), .B1(new_n444), .B2(new_n445), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n441), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n444), .A2(new_n445), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n263), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n444), .A2(new_n257), .A3(new_n445), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n450), .A2(KEYINPUT75), .A3(new_n451), .ZN(new_n452));
  XOR2_X1   g251(.A(G8gat), .B(G36gat), .Z(new_n453));
  XNOR2_X1  g252(.A(G64gat), .B(G92gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n453), .B(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n455), .B(KEYINPUT76), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n448), .A2(new_n452), .A3(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n450), .A2(new_n451), .A3(new_n455), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT30), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n446), .A2(new_n447), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n461), .A2(KEYINPUT30), .A3(new_n455), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n457), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n440), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n293), .A2(new_n404), .A3(new_n406), .A4(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n429), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n436), .A2(new_n437), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT80), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT80), .B1(new_n436), .B2(new_n437), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n463), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n400), .A2(new_n403), .ZN(new_n472));
  INV_X1    g271(.A(new_n205), .ZN(new_n473));
  INV_X1    g272(.A(new_n269), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n262), .A2(new_n263), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n279), .B1(new_n475), .B2(new_n206), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n474), .B1(new_n476), .B2(new_n264), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n275), .A2(new_n280), .ZN(new_n478));
  OAI21_X1  g277(.A(G22gat), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n289), .A2(new_n271), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n473), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n292), .B1(new_n481), .B2(KEYINPUT84), .ZN(new_n482));
  INV_X1    g281(.A(new_n287), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n471), .B(new_n472), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n465), .A2(KEYINPUT88), .B1(new_n484), .B2(KEYINPUT35), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n462), .A2(new_n460), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n486), .A2(new_n439), .A3(new_n438), .A4(new_n457), .ZN(new_n487));
  AOI22_X1  g286(.A1(new_n284), .A2(new_n285), .B1(new_n288), .B2(new_n291), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n487), .B1(new_n488), .B2(new_n287), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n405), .A2(KEYINPUT72), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n395), .A2(new_n397), .A3(new_n399), .ZN(new_n491));
  INV_X1    g290(.A(new_n385), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(new_n405), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n490), .B1(new_n494), .B2(new_n294), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT88), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n489), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT37), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n461), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT38), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT37), .B1(new_n446), .B2(new_n447), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n499), .A2(new_n500), .A3(new_n501), .A4(new_n456), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n429), .B(new_n458), .C1(new_n436), .C2(new_n437), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n448), .A2(new_n452), .A3(KEYINPUT37), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n455), .B1(new_n461), .B2(new_n498), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n502), .B(new_n504), .C1(new_n507), .C2(new_n500), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT40), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n413), .B1(new_n431), .B2(new_n432), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT86), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT86), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n422), .A2(new_n512), .A3(new_n413), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n408), .A2(new_n412), .A3(new_n410), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n511), .A2(new_n513), .A3(KEYINPUT39), .A4(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n427), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(KEYINPUT87), .B(KEYINPUT39), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n518), .B1(new_n511), .B2(new_n513), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n509), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n519), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n521), .A2(KEYINPUT40), .A3(new_n516), .A4(new_n515), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n463), .A2(new_n520), .A3(new_n434), .A4(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(new_n293), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n482), .A2(new_n483), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(new_n471), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT71), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n493), .A2(new_n529), .A3(KEYINPUT36), .A4(new_n405), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n493), .A2(KEYINPUT36), .A3(new_n405), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT71), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n530), .B(new_n532), .C1(new_n495), .C2(KEYINPUT36), .ZN(new_n533));
  AOI22_X1  g332(.A1(new_n485), .A2(new_n497), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(G43gat), .B(G50gat), .ZN(new_n535));
  INV_X1    g334(.A(G29gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT14), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(G36gat), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n536), .A2(KEYINPUT14), .ZN(new_n539));
  OAI211_X1 g338(.A(KEYINPUT15), .B(new_n535), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(G43gat), .B(G50gat), .Z(new_n541));
  INV_X1    g340(.A(KEYINPUT15), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n539), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n535), .A2(KEYINPUT15), .ZN(new_n544));
  INV_X1    g343(.A(G36gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n537), .B(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n540), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT17), .ZN(new_n549));
  XNOR2_X1  g348(.A(G15gat), .B(G22gat), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT90), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(G1gat), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT16), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n552), .A2(new_n553), .B1(new_n554), .B2(new_n550), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n550), .A2(new_n551), .A3(G1gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(G8gat), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT91), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n559), .B1(new_n550), .B2(G1gat), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n557), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n558), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n555), .A2(new_n562), .A3(new_n556), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(KEYINPUT92), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT92), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n561), .A2(new_n566), .A3(new_n563), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n549), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G229gat), .A2(G233gat), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n561), .A2(new_n563), .A3(new_n548), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT93), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT18), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n548), .B1(new_n561), .B2(new_n563), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n575), .A2(KEYINPUT94), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(KEYINPUT94), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n577), .A2(new_n570), .A3(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n569), .B(KEYINPUT13), .Z(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n572), .A2(new_n573), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n568), .A2(new_n569), .A3(new_n570), .A4(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n574), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G113gat), .B(G141gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(G197gat), .ZN(new_n586));
  XOR2_X1   g385(.A(KEYINPUT11), .B(G169gat), .Z(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT89), .B(KEYINPUT12), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n588), .B(new_n589), .Z(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n584), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n574), .A2(new_n581), .A3(new_n590), .A4(new_n583), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n534), .A2(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(G99gat), .B(G106gat), .Z(new_n597));
  INV_X1    g396(.A(KEYINPUT7), .ZN(new_n598));
  NAND2_X1  g397(.A1(G85gat), .A2(G92gat), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT101), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT102), .ZN(new_n602));
  NAND3_X1  g401(.A1(KEYINPUT101), .A2(G85gat), .A3(G92gat), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(G99gat), .ZN(new_n605));
  INV_X1    g404(.A(G106gat), .ZN(new_n606));
  OAI21_X1  g405(.A(KEYINPUT8), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OR2_X1    g406(.A1(KEYINPUT103), .A2(G92gat), .ZN(new_n608));
  INV_X1    g407(.A(G85gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(KEYINPUT103), .A2(G92gat), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n604), .A2(new_n607), .A3(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(KEYINPUT102), .B1(new_n599), .B2(KEYINPUT7), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n613), .B1(new_n603), .B2(new_n601), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n597), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(KEYINPUT104), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT104), .ZN(new_n617));
  OAI211_X1 g416(.A(new_n617), .B(new_n597), .C1(new_n612), .C2(new_n614), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n611), .A2(new_n607), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n601), .A2(new_n603), .ZN(new_n620));
  INV_X1    g419(.A(new_n613), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n597), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n619), .A2(new_n622), .A3(new_n623), .A4(new_n604), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n616), .A2(new_n618), .A3(new_n624), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n549), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G190gat), .B(G218gat), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n627), .A2(KEYINPUT105), .ZN(new_n628));
  AND2_X1   g427(.A1(G232gat), .A2(G233gat), .ZN(new_n629));
  AOI22_X1  g428(.A1(new_n627), .A2(KEYINPUT105), .B1(KEYINPUT41), .B2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n548), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n630), .B1(new_n625), .B2(new_n631), .ZN(new_n632));
  OR3_X1    g431(.A1(new_n626), .A2(new_n628), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n628), .B1(new_n626), .B2(new_n632), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n629), .A2(KEYINPUT41), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT100), .ZN(new_n637));
  XNOR2_X1  g436(.A(G134gat), .B(G162gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n635), .B(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G71gat), .B(G78gat), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(KEYINPUT95), .ZN(new_n645));
  XOR2_X1   g444(.A(G57gat), .B(G64gat), .Z(new_n646));
  INV_X1    g445(.A(KEYINPUT9), .ZN(new_n647));
  INV_X1    g446(.A(G71gat), .ZN(new_n648));
  INV_X1    g447(.A(G78gat), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT95), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n643), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n645), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n644), .A2(new_n646), .A3(KEYINPUT95), .A4(new_n650), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI22_X1  g455(.A1(new_n561), .A2(new_n563), .B1(KEYINPUT21), .B2(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n657), .B(KEYINPUT99), .Z(new_n658));
  XNOR2_X1  g457(.A(G127gat), .B(G155gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT20), .ZN(new_n660));
  NAND2_X1  g459(.A1(G231gat), .A2(G233gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT97), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n660), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n658), .B(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n656), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT96), .B(KEYINPUT21), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g466(.A(KEYINPUT98), .B(KEYINPUT19), .Z(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(G183gat), .B(G211gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n664), .B(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n642), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(G120gat), .B(G148gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(G176gat), .B(G204gat), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n674), .B(new_n675), .Z(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(G230gat), .A2(G233gat), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n656), .A2(new_n615), .A3(new_n624), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n680), .B1(new_n625), .B2(new_n665), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT10), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n625), .A2(new_n682), .A3(new_n665), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n679), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n681), .A2(new_n678), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n677), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  AOI211_X1 g487(.A(KEYINPUT10), .B(new_n680), .C1(new_n665), .C2(new_n625), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n678), .B1(new_n689), .B2(new_n684), .ZN(new_n690));
  INV_X1    g489(.A(new_n687), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n690), .A2(new_n691), .A3(new_n676), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT106), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n688), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  OAI211_X1 g493(.A(KEYINPUT106), .B(new_n677), .C1(new_n686), .C2(new_n687), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n673), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n596), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n469), .A2(new_n470), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(new_n553), .ZN(G1324gat));
  INV_X1    g501(.A(new_n699), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(new_n463), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT42), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n554), .A2(new_n558), .ZN(new_n706));
  NOR2_X1   g505(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OR3_X1    g507(.A1(new_n704), .A2(new_n705), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n705), .B1(new_n704), .B2(new_n708), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n704), .A2(G8gat), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(G1325gat));
  NAND2_X1  g511(.A1(new_n532), .A2(new_n530), .ZN(new_n713));
  AOI21_X1  g512(.A(KEYINPUT36), .B1(new_n404), .B2(new_n406), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n533), .A2(KEYINPUT107), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(G15gat), .B1(new_n699), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n404), .A2(new_n406), .ZN(new_n721));
  OR2_X1    g520(.A1(new_n721), .A2(G15gat), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n720), .B1(new_n699), .B2(new_n722), .ZN(G1326gat));
  NAND3_X1  g522(.A1(new_n703), .A2(KEYINPUT108), .A3(new_n526), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT108), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n725), .B1(new_n699), .B2(new_n293), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(KEYINPUT43), .B(G22gat), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1327gat));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n642), .A2(new_n672), .A3(new_n697), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n596), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT109), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n700), .A2(G29gat), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n733), .B1(new_n732), .B2(new_n734), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n730), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n737), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n739), .A2(KEYINPUT45), .A3(new_n735), .ZN(new_n740));
  INV_X1    g539(.A(new_n672), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n741), .A2(new_n594), .A3(new_n696), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n464), .B1(new_n482), .B2(new_n483), .ZN(new_n743));
  OAI21_X1  g542(.A(KEYINPUT88), .B1(new_n743), .B2(new_n721), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n484), .A2(KEYINPUT35), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n744), .A2(new_n745), .A3(new_n497), .ZN(new_n746));
  AOI22_X1  g545(.A1(new_n508), .A2(new_n523), .B1(new_n488), .B2(new_n287), .ZN(new_n747));
  AND3_X1   g546(.A1(new_n471), .A2(new_n488), .A3(new_n287), .ZN(new_n748));
  OAI22_X1  g547(.A1(new_n747), .A2(new_n748), .B1(new_n713), .B2(new_n714), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT110), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n746), .A2(KEYINPUT110), .A3(new_n749), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n642), .A2(KEYINPUT44), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n750), .A2(new_n641), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT44), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n742), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n700), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n738), .B(new_n740), .C1(new_n536), .C2(new_n760), .ZN(G1328gat));
  AOI21_X1  g560(.A(G36gat), .B1(KEYINPUT111), .B2(KEYINPUT46), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n732), .A2(new_n463), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n763), .B(new_n764), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n758), .A2(new_n463), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n765), .B1(new_n545), .B2(new_n766), .ZN(G1329gat));
  NOR2_X1   g566(.A1(new_n721), .A2(G43gat), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n732), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n769), .A2(KEYINPUT112), .ZN(new_n770));
  INV_X1    g569(.A(G43gat), .ZN(new_n771));
  INV_X1    g570(.A(new_n719), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n771), .B1(new_n758), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(KEYINPUT47), .A2(G43gat), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n775), .B1(new_n758), .B2(new_n715), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n769), .B1(KEYINPUT112), .B2(KEYINPUT47), .ZN(new_n777));
  OAI22_X1  g576(.A1(new_n774), .A2(KEYINPUT47), .B1(new_n776), .B2(new_n777), .ZN(G1330gat));
  NAND3_X1  g577(.A1(new_n758), .A2(G50gat), .A3(new_n526), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(G50gat), .B1(new_n732), .B2(new_n526), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT48), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT48), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n732), .A2(new_n526), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n779), .B(new_n783), .C1(G50gat), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n782), .A2(new_n785), .ZN(G1331gat));
  AND2_X1   g585(.A1(new_n752), .A2(new_n753), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n673), .A2(new_n594), .A3(new_n696), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n759), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g591(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n793), .B1(new_n790), .B2(new_n463), .ZN(new_n794));
  INV_X1    g593(.A(new_n463), .ZN(new_n795));
  XOR2_X1   g594(.A(KEYINPUT49), .B(G64gat), .Z(new_n796));
  NOR3_X1   g595(.A1(new_n789), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT113), .B1(new_n794), .B2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT113), .ZN(new_n799));
  OAI22_X1  g598(.A1(new_n789), .A2(new_n795), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n790), .A2(new_n463), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n799), .B(new_n800), .C1(new_n801), .C2(new_n796), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n798), .A2(new_n802), .ZN(G1333gat));
  OAI21_X1  g602(.A(G71gat), .B1(new_n789), .B2(new_n719), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n787), .A2(new_n648), .A3(new_n495), .A4(new_n788), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT50), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n804), .A2(KEYINPUT50), .A3(new_n805), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(G1334gat));
  NOR2_X1   g609(.A1(new_n789), .A2(new_n293), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(new_n649), .ZN(G1335gat));
  INV_X1    g611(.A(KEYINPUT51), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n672), .A2(new_n594), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n642), .B1(new_n746), .B2(new_n749), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AOI211_X1 g616(.A(KEYINPUT115), .B(new_n642), .C1(new_n746), .C2(new_n749), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n813), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(KEYINPUT115), .B1(new_n534), .B2(new_n642), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n750), .A2(new_n816), .A3(new_n641), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n820), .A2(KEYINPUT51), .A3(new_n814), .A4(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n696), .B1(new_n819), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n823), .A2(new_n609), .A3(new_n759), .ZN(new_n824));
  INV_X1    g623(.A(new_n814), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n825), .A2(new_n696), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n827), .B1(new_n755), .B2(new_n757), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n759), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT114), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(G85gat), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n829), .A2(KEYINPUT114), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n824), .B1(new_n831), .B2(new_n832), .ZN(G1336gat));
  AND2_X1   g632(.A1(new_n608), .A2(new_n610), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n834), .B1(new_n828), .B2(new_n463), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n696), .A2(new_n795), .ZN(new_n837));
  INV_X1    g636(.A(G92gat), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n839), .B1(new_n819), .B2(new_n822), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  XNOR2_X1  g640(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n836), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n842), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n844), .B1(new_n835), .B2(new_n840), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(G1337gat));
  NAND3_X1  g645(.A1(new_n823), .A2(new_n605), .A3(new_n495), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n828), .A2(new_n772), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n847), .B1(new_n605), .B2(new_n848), .ZN(G1338gat));
  NOR2_X1   g648(.A1(new_n293), .A2(G106gat), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  AOI211_X1 g650(.A(new_n696), .B(new_n851), .C1(new_n819), .C2(new_n822), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n606), .B1(new_n828), .B2(new_n526), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT53), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n819), .A2(new_n822), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n697), .A3(new_n850), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n828), .A2(new_n526), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(G106gat), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n856), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n854), .A2(new_n860), .ZN(G1339gat));
  NOR3_X1   g660(.A1(new_n673), .A2(new_n594), .A3(new_n697), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n569), .B1(new_n568), .B2(new_n570), .ZN(new_n863));
  OAI22_X1  g662(.A1(new_n863), .A2(KEYINPUT118), .B1(new_n579), .B2(new_n580), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT118), .ZN(new_n865));
  AOI211_X1 g664(.A(new_n865), .B(new_n569), .C1(new_n568), .C2(new_n570), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n588), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n867), .A2(new_n593), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n697), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n683), .A2(new_n685), .A3(new_n679), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n690), .A2(KEYINPUT54), .A3(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT54), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n872), .B(new_n678), .C1(new_n689), .C2(new_n684), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT117), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n873), .A2(new_n874), .A3(new_n677), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n874), .B1(new_n873), .B2(new_n677), .ZN(new_n876));
  OAI211_X1 g675(.A(KEYINPUT55), .B(new_n871), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n877), .A2(new_n594), .A3(new_n692), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n871), .B1(new_n875), .B2(new_n876), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT55), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n869), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n642), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n879), .A2(new_n880), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n884), .A2(new_n641), .A3(new_n868), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n877), .A2(new_n692), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n862), .B1(new_n888), .B2(new_n741), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n889), .A2(new_n700), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n526), .A2(new_n494), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n890), .A2(new_n795), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(new_n298), .A3(new_n594), .ZN(new_n893));
  INV_X1    g692(.A(new_n862), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n885), .A2(new_n886), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n895), .B1(new_n642), .B2(new_n882), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n894), .B1(new_n896), .B2(new_n672), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n721), .A2(new_n526), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n700), .A2(new_n463), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n298), .B1(new_n901), .B2(new_n594), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT119), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n902), .A2(new_n903), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n893), .B1(new_n904), .B2(new_n905), .ZN(G1340gat));
  AOI21_X1  g705(.A(G120gat), .B1(new_n892), .B2(new_n697), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n696), .A2(new_n299), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n901), .B2(new_n908), .ZN(G1341gat));
  INV_X1    g708(.A(new_n901), .ZN(new_n910));
  OAI21_X1  g709(.A(G127gat), .B1(new_n910), .B2(new_n741), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n892), .A2(new_n303), .A3(new_n672), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1342gat));
  NAND3_X1  g712(.A1(new_n892), .A2(new_n376), .A3(new_n641), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n914), .A2(KEYINPUT56), .ZN(new_n915));
  OAI21_X1  g714(.A(G134gat), .B1(new_n910), .B2(new_n642), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(KEYINPUT56), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(G1343gat));
  AOI21_X1  g717(.A(new_n293), .B1(new_n717), .B2(new_n718), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n890), .A2(new_n795), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n211), .B1(new_n920), .B2(new_n595), .ZN(new_n921));
  AND4_X1   g720(.A1(new_n593), .A2(new_n867), .A3(new_n694), .A4(new_n695), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n879), .A2(KEYINPUT120), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT120), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n924), .B(new_n871), .C1(new_n875), .C2(new_n876), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n923), .A2(new_n880), .A3(new_n925), .ZN(new_n926));
  AND3_X1   g725(.A1(new_n877), .A2(new_n594), .A3(new_n692), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n922), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n887), .B1(new_n928), .B2(new_n641), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n862), .B1(new_n929), .B2(new_n741), .ZN(new_n930));
  OAI21_X1  g729(.A(KEYINPUT57), .B1(new_n930), .B2(new_n293), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT57), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n897), .A2(new_n932), .A3(new_n526), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n533), .A2(new_n900), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n931), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n594), .A2(G141gat), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n921), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT58), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n921), .B(KEYINPUT58), .C1(new_n935), .C2(new_n936), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(G1344gat));
  INV_X1    g740(.A(new_n920), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n942), .A2(new_n209), .A3(new_n697), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT59), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT121), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n672), .B1(new_n929), .B2(new_n945), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n887), .B(KEYINPUT121), .C1(new_n928), .C2(new_n641), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n862), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n526), .A2(new_n932), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g749(.A(KEYINPUT57), .B1(new_n889), .B2(new_n293), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n950), .A2(new_n697), .A3(new_n934), .A4(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n944), .B1(new_n952), .B2(G148gat), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n935), .A2(new_n696), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n954), .A2(KEYINPUT59), .A3(new_n209), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n943), .B1(new_n953), .B2(new_n955), .ZN(G1345gat));
  NAND3_X1  g755(.A1(new_n942), .A2(new_n218), .A3(new_n672), .ZN(new_n957));
  OAI21_X1  g756(.A(G155gat), .B1(new_n935), .B2(new_n741), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1346gat));
  AOI21_X1  g758(.A(G162gat), .B1(new_n942), .B2(new_n641), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n935), .A2(new_n219), .A3(new_n642), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n960), .A2(new_n961), .ZN(G1347gat));
  NOR2_X1   g761(.A1(new_n759), .A2(new_n795), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n899), .A2(new_n963), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n964), .A2(new_n328), .A3(new_n595), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n889), .A2(new_n759), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n966), .A2(new_n891), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n967), .A2(new_n594), .A3(new_n463), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n965), .B1(new_n968), .B2(new_n328), .ZN(G1348gat));
  NAND3_X1  g768(.A1(new_n967), .A2(new_n329), .A3(new_n837), .ZN(new_n970));
  OAI21_X1  g769(.A(G176gat), .B1(new_n964), .B2(new_n696), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT122), .ZN(G1349gat));
  NAND4_X1  g772(.A1(new_n897), .A2(new_n672), .A3(new_n898), .A4(new_n963), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n346), .B1(new_n974), .B2(KEYINPUT123), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n975), .B1(KEYINPUT123), .B2(new_n974), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n967), .A2(new_n463), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n672), .A2(new_n359), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(KEYINPUT60), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT60), .ZN(new_n981));
  OAI211_X1 g780(.A(new_n976), .B(new_n981), .C1(new_n977), .C2(new_n978), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n980), .A2(new_n982), .ZN(G1350gat));
  NAND3_X1  g782(.A1(new_n899), .A2(new_n641), .A3(new_n963), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT61), .ZN(new_n985));
  AND3_X1   g784(.A1(new_n984), .A2(new_n985), .A3(G190gat), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n985), .B1(new_n984), .B2(G190gat), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n641), .A2(new_n350), .ZN(new_n988));
  OAI22_X1  g787(.A1(new_n986), .A2(new_n987), .B1(new_n977), .B2(new_n988), .ZN(G1351gat));
  NAND2_X1  g788(.A1(new_n719), .A2(new_n963), .ZN(new_n990));
  INV_X1    g789(.A(new_n990), .ZN(new_n991));
  OAI211_X1 g790(.A(new_n951), .B(new_n991), .C1(new_n948), .C2(new_n949), .ZN(new_n992));
  INV_X1    g791(.A(G197gat), .ZN(new_n993));
  NOR3_X1   g792(.A1(new_n992), .A2(new_n993), .A3(new_n595), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n966), .A2(new_n463), .A3(new_n919), .ZN(new_n995));
  XNOR2_X1  g794(.A(new_n995), .B(KEYINPUT124), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n996), .A2(new_n594), .ZN(new_n997));
  AOI21_X1  g796(.A(new_n994), .B1(new_n997), .B2(new_n993), .ZN(G1352gat));
  XOR2_X1   g797(.A(KEYINPUT125), .B(G204gat), .Z(new_n999));
  OAI211_X1 g798(.A(new_n697), .B(new_n951), .C1(new_n948), .C2(new_n949), .ZN(new_n1000));
  OAI21_X1  g799(.A(new_n999), .B1(new_n1000), .B2(new_n990), .ZN(new_n1001));
  NOR3_X1   g800(.A1(new_n696), .A2(new_n795), .A3(new_n999), .ZN(new_n1002));
  NAND4_X1  g801(.A1(new_n919), .A2(new_n897), .A3(new_n700), .A4(new_n1002), .ZN(new_n1003));
  INV_X1    g802(.A(KEYINPUT62), .ZN(new_n1004));
  XNOR2_X1  g803(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1001), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g805(.A(KEYINPUT126), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n1001), .A2(KEYINPUT126), .A3(new_n1005), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1008), .A2(new_n1009), .ZN(G1353gat));
  INV_X1    g809(.A(G211gat), .ZN(new_n1011));
  NAND3_X1  g810(.A1(new_n996), .A2(new_n1011), .A3(new_n672), .ZN(new_n1012));
  NAND4_X1  g811(.A1(new_n950), .A2(new_n672), .A3(new_n951), .A4(new_n991), .ZN(new_n1013));
  AOI21_X1  g812(.A(KEYINPUT63), .B1(new_n1013), .B2(G211gat), .ZN(new_n1014));
  OAI211_X1 g813(.A(KEYINPUT63), .B(G211gat), .C1(new_n992), .C2(new_n741), .ZN(new_n1015));
  INV_X1    g814(.A(new_n1015), .ZN(new_n1016));
  OAI21_X1  g815(.A(new_n1012), .B1(new_n1014), .B2(new_n1016), .ZN(G1354gat));
  AOI21_X1  g816(.A(G218gat), .B1(new_n996), .B2(new_n641), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n641), .A2(G218gat), .ZN(new_n1019));
  XOR2_X1   g818(.A(new_n1019), .B(KEYINPUT127), .Z(new_n1020));
  NOR2_X1   g819(.A1(new_n992), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g820(.A1(new_n1018), .A2(new_n1021), .ZN(G1355gat));
endmodule


