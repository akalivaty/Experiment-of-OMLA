//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 1 1 1 1 0 0 0 1 1 0 0 0 1 0 0 1 1 1 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1230, new_n1231,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  AND3_X1   g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G107), .A2(G264), .ZN(new_n208));
  INV_X1    g0008(.A(G68), .ZN(new_n209));
  INV_X1    g0009(.A(G238), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n207), .B(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  AOI21_X1  g0011(.A(new_n211), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G50), .ZN(new_n213));
  INV_X1    g0013(.A(G226), .ZN(new_n214));
  INV_X1    g0014(.A(G244), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n202), .C2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G58), .ZN(new_n217));
  INV_X1    g0017(.A(G232), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n206), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT66), .Z(new_n222));
  NOR2_X1   g0022(.A1(new_n206), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT0), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n222), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OR2_X1    g0030(.A1(new_n203), .A2(KEYINPUT65), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n203), .A2(KEYINPUT65), .ZN(new_n232));
  NAND3_X1  g0032(.A1(new_n231), .A2(G50), .A3(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n227), .B1(new_n230), .B2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G264), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n237), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G226), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n238), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(new_n213), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n217), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  OAI21_X1  g0052(.A(KEYINPUT70), .B1(new_n206), .B2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT70), .ZN(new_n254));
  NAND4_X1  g0054(.A1(new_n254), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n253), .A2(new_n228), .A3(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT71), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G58), .ZN(new_n258));
  XOR2_X1   g0058(.A(new_n258), .B(KEYINPUT8), .Z(new_n259));
  NOR2_X1   g0059(.A1(new_n252), .A2(G20), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G150), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G20), .A2(G33), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  OAI22_X1  g0064(.A1(new_n259), .A2(new_n261), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n229), .B1(new_n201), .B2(new_n203), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n256), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n256), .ZN(new_n268));
  INV_X1    g0068(.A(G1), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT68), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT68), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G1), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G20), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n268), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G50), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT72), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT68), .B(G1), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n278), .A2(new_n229), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G13), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n213), .ZN(new_n281));
  AND3_X1   g0081(.A1(new_n276), .A2(new_n277), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n277), .B1(new_n276), .B2(new_n281), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n267), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT9), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT10), .ZN(new_n287));
  OR2_X1    g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(KEYINPUT3), .A2(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G223), .ZN(new_n291));
  INV_X1    g0091(.A(G1698), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT69), .B(G1698), .ZN(new_n293));
  INV_X1    g0093(.A(G222), .ZN(new_n294));
  OAI221_X1 g0094(.A(new_n290), .B1(new_n291), .B2(new_n292), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G41), .ZN(new_n296));
  OAI211_X1 g0096(.A(G1), .B(G13), .C1(new_n252), .C2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n295), .B(new_n298), .C1(G77), .C2(new_n290), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n269), .B(G274), .C1(G41), .C2(G45), .ZN(new_n300));
  NOR2_X1   g0100(.A1(G41), .A2(G45), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n297), .B1(new_n278), .B2(new_n301), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n299), .B(new_n300), .C1(new_n214), .C2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G190), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI211_X1 g0105(.A(KEYINPUT9), .B(new_n267), .C1(new_n282), .C2(new_n283), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n286), .A2(new_n287), .A3(new_n305), .A4(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT74), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n303), .A2(G200), .ZN(new_n309));
  OR3_X1    g0109(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n308), .B1(new_n307), .B2(new_n309), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n286), .A2(new_n305), .A3(new_n306), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT75), .ZN(new_n314));
  OR2_X1    g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n309), .B1(new_n313), .B2(new_n314), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n287), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n303), .A2(G179), .ZN(new_n320));
  INV_X1    g0120(.A(G169), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n303), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n320), .A2(new_n284), .A3(new_n322), .ZN(new_n323));
  XNOR2_X1  g0123(.A(KEYINPUT8), .B(G58), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n325), .A2(new_n263), .B1(G20), .B2(G77), .ZN(new_n326));
  XOR2_X1   g0126(.A(KEYINPUT15), .B(G87), .Z(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n260), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n268), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n329), .B(KEYINPUT73), .ZN(new_n330));
  INV_X1    g0130(.A(G13), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n274), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n330), .B1(new_n202), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n275), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G77), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  OAI221_X1 g0136(.A(new_n290), .B1(new_n210), .B2(new_n292), .C1(new_n293), .C2(new_n218), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n337), .B(new_n298), .C1(G107), .C2(new_n290), .ZN(new_n338));
  OR2_X1    g0138(.A1(new_n302), .A2(new_n215), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n338), .A2(new_n300), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n321), .ZN(new_n341));
  INV_X1    g0141(.A(new_n340), .ZN(new_n342));
  INV_X1    g0142(.A(G179), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n336), .A2(new_n341), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n319), .A2(new_n323), .A3(new_n345), .ZN(new_n346));
  OAI22_X1  g0146(.A1(new_n293), .A2(new_n214), .B1(new_n218), .B2(new_n292), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n347), .A2(new_n290), .B1(G33), .B2(G97), .ZN(new_n348));
  OAI221_X1 g0148(.A(new_n300), .B1(new_n210), .B2(new_n302), .C1(new_n348), .C2(new_n297), .ZN(new_n349));
  OR2_X1    g0149(.A1(new_n349), .A2(KEYINPUT13), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(KEYINPUT13), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT14), .B1(new_n353), .B2(new_n321), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(G179), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT14), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n352), .A2(new_n356), .A3(G169), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n354), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n332), .A2(new_n209), .ZN(new_n359));
  XNOR2_X1  g0159(.A(new_n359), .B(KEYINPUT12), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n260), .A2(G77), .B1(G20), .B2(new_n209), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(new_n213), .B2(new_n264), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n362), .A2(KEYINPUT11), .A3(new_n256), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT11), .B1(new_n362), .B2(new_n256), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n364), .B1(G68), .B2(new_n334), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n360), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n358), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G200), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n353), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n366), .B1(new_n352), .B2(new_n304), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n259), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n275), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n280), .A2(new_n259), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n288), .A2(new_n229), .A3(new_n289), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT7), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n288), .A2(KEYINPUT7), .A3(new_n229), .A4(new_n289), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G68), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n217), .A2(new_n209), .ZN(new_n385));
  OAI21_X1  g0185(.A(G20), .B1(new_n385), .B2(new_n203), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n263), .A2(G159), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n384), .A2(KEYINPUT16), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n256), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT76), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n381), .A2(new_n392), .A3(new_n382), .ZN(new_n393));
  OR2_X1    g0193(.A1(new_n382), .A2(new_n392), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n393), .A2(G68), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT16), .B1(new_n395), .B2(new_n389), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n378), .B1(new_n391), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n292), .A2(KEYINPUT69), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT69), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G1698), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n291), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n214), .A2(new_n292), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n290), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G33), .A2(G87), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n298), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT78), .ZN(new_n407));
  OAI211_X1 g0207(.A(G232), .B(new_n297), .C1(new_n278), .C2(new_n301), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n407), .B1(new_n408), .B2(new_n300), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n408), .A2(new_n407), .A3(new_n300), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n406), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n321), .ZN(new_n413));
  AND3_X1   g0213(.A1(new_n408), .A2(new_n407), .A3(new_n300), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n414), .A2(new_n409), .ZN(new_n415));
  AOI21_X1  g0215(.A(KEYINPUT77), .B1(new_n405), .B2(new_n298), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT77), .ZN(new_n417));
  AOI211_X1 g0217(.A(new_n417), .B(new_n297), .C1(new_n403), .C2(new_n404), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n415), .B(new_n343), .C1(new_n416), .C2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n397), .A2(new_n413), .A3(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT18), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n397), .A2(KEYINPUT18), .A3(new_n413), .A4(new_n419), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT17), .ZN(new_n425));
  XNOR2_X1  g0225(.A(KEYINPUT79), .B(G190), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n415), .B(new_n427), .C1(new_n416), .C2(new_n418), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n412), .A2(new_n369), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n395), .A2(new_n389), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT16), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n388), .B1(new_n383), .B2(G68), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n268), .B1(new_n434), .B2(KEYINPUT16), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n433), .A2(new_n435), .B1(new_n376), .B2(new_n377), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n430), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n425), .B1(new_n437), .B2(KEYINPUT80), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT80), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n430), .A2(new_n436), .A3(new_n439), .A4(KEYINPUT17), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n424), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n342), .A2(new_n369), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n340), .A2(new_n304), .ZN(new_n443));
  NOR3_X1   g0243(.A1(new_n336), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  OR3_X1    g0244(.A1(new_n374), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n346), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT94), .ZN(new_n448));
  XNOR2_X1  g0248(.A(KEYINPUT88), .B(KEYINPUT22), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n290), .A2(new_n449), .A3(new_n229), .A4(G87), .ZN(new_n450));
  AND2_X1   g0250(.A1(KEYINPUT3), .A2(G33), .ZN(new_n451));
  NOR2_X1   g0251(.A1(KEYINPUT3), .A2(G33), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n229), .B(G87), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT88), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(KEYINPUT22), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n229), .A2(G33), .A3(G116), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT23), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n458), .B1(new_n229), .B2(G107), .ZN(new_n459));
  INV_X1    g0259(.A(G107), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n460), .A2(KEYINPUT23), .A3(G20), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n450), .A2(new_n456), .A3(new_n457), .A4(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT89), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n453), .A2(new_n455), .B1(new_n459), .B2(new_n461), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT89), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n465), .A2(new_n466), .A3(new_n450), .A4(new_n457), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n464), .A2(KEYINPUT24), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(KEYINPUT24), .B1(new_n464), .B2(new_n467), .ZN(new_n469));
  NOR3_X1   g0269(.A1(new_n468), .A2(new_n469), .A3(new_n268), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT91), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n279), .A2(G13), .A3(new_n460), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT25), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n472), .A2(new_n471), .A3(new_n473), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT90), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n477), .B1(new_n472), .B2(new_n473), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n332), .A2(KEYINPUT90), .A3(KEYINPUT25), .A4(new_n460), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n475), .A2(new_n476), .A3(new_n478), .A4(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n273), .A2(G33), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n280), .A2(new_n268), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n480), .B1(new_n460), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(KEYINPUT92), .B1(new_n470), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n464), .A2(new_n467), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT24), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n464), .A2(KEYINPUT24), .A3(new_n467), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n487), .A2(new_n256), .A3(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n476), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n490), .A2(new_n474), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n478), .A2(new_n479), .ZN(new_n492));
  INV_X1    g0292(.A(new_n482), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n491), .A2(new_n492), .B1(G107), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT92), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n489), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  OR2_X1    g0296(.A1(new_n296), .A2(KEYINPUT5), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n273), .A2(G45), .A3(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT83), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n296), .A2(KEYINPUT5), .ZN(new_n501));
  INV_X1    g0301(.A(G45), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n502), .B1(new_n270), .B2(new_n272), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n503), .A2(KEYINPUT83), .A3(new_n497), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n500), .A2(new_n501), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(G264), .A3(new_n297), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(KEYINPUT93), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT93), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n505), .A2(new_n508), .A3(G264), .A4(new_n297), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n451), .A2(new_n452), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n398), .A2(new_n400), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G250), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G257), .A2(G1698), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(G294), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n252), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n298), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n500), .A2(G274), .A3(new_n501), .A4(new_n504), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n518), .B1(new_n519), .B2(new_n298), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n510), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G169), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n510), .A2(G179), .A3(new_n521), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n484), .A2(new_n496), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n520), .B1(new_n507), .B2(new_n509), .ZN(new_n526));
  AND2_X1   g0326(.A1(new_n526), .A2(G190), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n489), .A2(new_n494), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n369), .B1(new_n510), .B2(new_n521), .ZN(new_n529));
  NOR3_X1   g0329(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n448), .B1(new_n525), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n524), .B1(new_n321), .B2(new_n526), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n489), .A2(new_n495), .A3(new_n494), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n495), .B1(new_n489), .B2(new_n494), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n529), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n526), .A2(G190), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n536), .A2(new_n489), .A3(new_n494), .A4(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n535), .A2(KEYINPUT94), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n531), .A2(new_n539), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n500), .A2(new_n504), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n541), .A2(G274), .A3(new_n297), .A4(new_n501), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G264), .A2(G1698), .ZN(new_n543));
  INV_X1    g0343(.A(G257), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n290), .B(new_n543), .C1(new_n293), .C2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(G303), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n297), .B1(new_n511), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(KEYINPUT86), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT86), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n545), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n505), .A2(G270), .A3(new_n297), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n542), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT20), .ZN(new_n555));
  NAND2_X1  g0355(.A1(G33), .A2(G283), .ZN(new_n556));
  OR2_X1    g0356(.A1(KEYINPUT81), .A2(G97), .ZN(new_n557));
  NAND2_X1  g0357(.A1(KEYINPUT81), .A2(G97), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n229), .B(new_n556), .C1(new_n559), .C2(G33), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(G116), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(G20), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n256), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n555), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n560), .A2(KEYINPUT20), .A3(new_n256), .A4(new_n563), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n280), .A2(G116), .A3(new_n268), .A4(new_n481), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n332), .A2(new_n562), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n554), .A2(G169), .A3(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT21), .ZN(new_n572));
  INV_X1    g0372(.A(new_n554), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n565), .A2(new_n566), .B1(new_n562), .B2(new_n332), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n343), .B1(new_n574), .B2(new_n568), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n571), .A2(new_n572), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT87), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(new_n571), .B2(new_n572), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n321), .B1(new_n574), .B2(new_n568), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n579), .A2(KEYINPUT87), .A3(KEYINPUT21), .A4(new_n554), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n576), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n554), .A2(G200), .ZN(new_n582));
  INV_X1    g0382(.A(new_n570), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n582), .B(new_n583), .C1(new_n427), .C2(new_n554), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n505), .A2(G257), .A3(new_n297), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n290), .A2(new_n512), .A3(G244), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT4), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n290), .A2(new_n512), .A3(KEYINPUT4), .A4(G244), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n290), .A2(G250), .A3(G1698), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n589), .A2(new_n556), .A3(new_n590), .A4(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n298), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n542), .A2(new_n586), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G169), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n343), .B2(new_n594), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n557), .A2(KEYINPUT6), .A3(new_n460), .A4(new_n558), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT82), .ZN(new_n598));
  OR2_X1    g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT6), .ZN(new_n600));
  INV_X1    g0400(.A(G97), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n601), .A2(new_n460), .ZN(new_n602));
  NOR2_X1   g0402(.A1(G97), .A2(G107), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n600), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n597), .A2(new_n598), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n599), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G20), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n393), .A2(G107), .A3(new_n394), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n263), .A2(G77), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n610), .A2(new_n256), .B1(new_n601), .B2(new_n332), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT84), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n493), .A2(G97), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n612), .B1(new_n611), .B2(new_n613), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n596), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n493), .A2(new_n327), .ZN(new_n617));
  NAND3_X1  g0417(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n229), .ZN(new_n619));
  INV_X1    g0419(.A(new_n558), .ZN(new_n620));
  NOR2_X1   g0420(.A1(KEYINPUT81), .A2(G97), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(G87), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n460), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n619), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n290), .A2(new_n229), .A3(G68), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n559), .A2(new_n261), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n625), .B(new_n626), .C1(new_n627), .C2(KEYINPUT19), .ZN(new_n628));
  INV_X1    g0428(.A(new_n327), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n628), .A2(new_n256), .B1(new_n332), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT85), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n617), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n631), .B1(new_n617), .B2(new_n630), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(G274), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n503), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(G250), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n637), .B1(new_n278), .B2(new_n502), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n636), .A2(new_n638), .A3(new_n297), .ZN(new_n639));
  OAI22_X1  g0439(.A1(new_n293), .A2(new_n210), .B1(new_n215), .B2(new_n292), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n640), .A2(new_n290), .B1(G33), .B2(G116), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n639), .B1(new_n641), .B2(new_n297), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(G169), .ZN(new_n643));
  OAI211_X1 g0443(.A(G179), .B(new_n639), .C1(new_n641), .C2(new_n297), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n642), .A2(G200), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n493), .A2(G87), .ZN(new_n647));
  OAI211_X1 g0447(.A(G190), .B(new_n639), .C1(new_n641), .C2(new_n297), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n647), .A2(new_n630), .A3(new_n648), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n634), .A2(new_n645), .B1(new_n646), .B2(new_n649), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n594), .A2(new_n304), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n594), .A2(G200), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n651), .A2(new_n613), .A3(new_n611), .A4(new_n652), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n616), .A2(new_n650), .A3(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n540), .A2(new_n585), .A3(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n447), .A2(new_n655), .ZN(G372));
  NAND2_X1  g0456(.A1(new_n617), .A2(new_n630), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n645), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n650), .B(new_n596), .C1(new_n615), .C2(new_n614), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(KEYINPUT26), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n649), .A2(new_n646), .B1(new_n645), .B2(new_n657), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n611), .A2(new_n613), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT26), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n596), .A2(new_n662), .A3(new_n663), .A4(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT95), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n526), .A2(new_n321), .ZN(new_n667));
  AOI211_X1 g0467(.A(new_n343), .B(new_n520), .C1(new_n507), .C2(new_n509), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n666), .B(new_n528), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n666), .B1(new_n532), .B2(new_n528), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n576), .A2(new_n578), .A3(new_n580), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n616), .A2(new_n538), .A3(new_n653), .A4(new_n662), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n661), .B(new_n665), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n446), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n323), .ZN(new_n677));
  INV_X1    g0477(.A(new_n345), .ZN(new_n678));
  AOI22_X1  g0478(.A1(new_n373), .A2(new_n678), .B1(new_n358), .B2(new_n367), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n438), .A2(new_n440), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n424), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n677), .B1(new_n681), .B2(new_n319), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n676), .A2(new_n682), .ZN(G369));
  INV_X1    g0483(.A(G330), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n331), .A2(G20), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  OR3_X1    g0486(.A1(new_n278), .A2(new_n686), .A3(KEYINPUT27), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT27), .B1(new_n278), .B2(new_n686), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(new_n688), .A3(G213), .ZN(new_n689));
  INV_X1    g0489(.A(G343), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  OAI211_X1 g0492(.A(new_n581), .B(new_n584), .C1(new_n583), .C2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n672), .A2(new_n570), .A3(new_n691), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n684), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n691), .B1(new_n533), .B2(new_n534), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n540), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n525), .A2(new_n691), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n695), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n581), .B1(new_n531), .B2(new_n539), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n670), .A2(new_n671), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n692), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n700), .A2(new_n704), .ZN(G399));
  INV_X1    g0505(.A(new_n223), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G41), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G1), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n559), .A2(new_n623), .A3(new_n460), .A4(new_n562), .ZN(new_n710));
  OAI22_X1  g0510(.A1(new_n709), .A2(new_n710), .B1(new_n233), .B2(new_n708), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n596), .A2(new_n662), .A3(new_n663), .A4(KEYINPUT26), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT96), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n660), .A2(new_n664), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n659), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n616), .A2(new_n653), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT97), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n581), .A2(new_n720), .A3(new_n535), .ZN(new_n721));
  OAI21_X1  g0521(.A(KEYINPUT97), .B1(new_n525), .B2(new_n672), .ZN(new_n722));
  INV_X1    g0522(.A(new_n662), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n530), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n719), .A2(new_n721), .A3(new_n722), .A4(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n691), .B1(new_n717), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(KEYINPUT29), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n675), .A2(new_n692), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n727), .B1(new_n729), .B2(KEYINPUT29), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n593), .A2(new_n586), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(new_n642), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n668), .A2(new_n573), .A3(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT30), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n573), .A2(new_n526), .A3(G179), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(new_n642), .A3(new_n594), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n735), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n739), .A2(KEYINPUT31), .A3(new_n691), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n691), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT31), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n740), .B(new_n743), .C1(new_n655), .C2(new_n691), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G330), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n730), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n712), .B1(new_n747), .B2(G1), .ZN(G364));
  NAND2_X1  g0548(.A1(new_n693), .A2(new_n694), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G330), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n709), .B1(G45), .B2(new_n685), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n693), .A2(new_n684), .A3(new_n694), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n750), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  XOR2_X1   g0554(.A(new_n754), .B(KEYINPUT98), .Z(new_n755));
  AOI21_X1  g0555(.A(new_n228), .B1(G20), .B2(new_n321), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n229), .A2(G179), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n758), .A2(new_n304), .A3(G200), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n460), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n343), .A2(new_n369), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n426), .A2(G20), .A3(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n229), .A2(G190), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n763), .A2(G50), .B1(G68), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n343), .A2(G200), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n764), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n767), .B1(new_n202), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n426), .A2(G20), .A3(new_n768), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n217), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G179), .A2(G200), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n764), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  XOR2_X1   g0575(.A(KEYINPUT101), .B(G159), .Z(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT32), .ZN(new_n778));
  OR4_X1    g0578(.A1(new_n760), .A2(new_n770), .A3(new_n772), .A4(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n229), .B1(new_n773), .B2(G190), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n601), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n758), .A2(G190), .A3(G200), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n623), .ZN(new_n783));
  NOR4_X1   g0583(.A1(new_n779), .A2(new_n511), .A3(new_n781), .A4(new_n783), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n784), .B(KEYINPUT102), .Z(new_n785));
  INV_X1    g0585(.A(new_n759), .ZN(new_n786));
  INV_X1    g0586(.A(new_n780), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n786), .A2(G283), .B1(new_n787), .B2(G294), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n775), .A2(G329), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n788), .A2(new_n511), .A3(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G311), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n769), .A2(new_n791), .ZN(new_n792));
  OR2_X1    g0592(.A1(KEYINPUT33), .A2(G317), .ZN(new_n793));
  NAND2_X1  g0593(.A1(KEYINPUT33), .A2(G317), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n765), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n782), .A2(new_n546), .ZN(new_n796));
  NOR4_X1   g0596(.A1(new_n790), .A2(new_n792), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n763), .A2(G326), .ZN(new_n798));
  INV_X1    g0598(.A(G322), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n797), .B(new_n798), .C1(new_n799), .C2(new_n771), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT103), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n757), .B1(new_n785), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(G13), .A2(G33), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(G20), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n756), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  XOR2_X1   g0607(.A(G355), .B(KEYINPUT99), .Z(new_n808));
  NAND3_X1  g0608(.A1(new_n808), .A2(new_n223), .A3(new_n290), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(G116), .B2(new_n223), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT100), .Z(new_n811));
  NAND2_X1  g0611(.A1(new_n247), .A2(G45), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n706), .A2(new_n290), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n812), .B(new_n813), .C1(G45), .C2(new_n233), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n807), .B1(new_n811), .B2(new_n814), .ZN(new_n815));
  NOR3_X1   g0615(.A1(new_n802), .A2(new_n815), .A3(new_n752), .ZN(new_n816));
  INV_X1    g0616(.A(new_n805), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n816), .B1(new_n749), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n755), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT104), .ZN(G396));
  NOR2_X1   g0620(.A1(new_n345), .A2(new_n691), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n692), .B1(new_n333), .B2(new_n335), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n345), .B1(new_n444), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n803), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n756), .A2(new_n803), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n202), .ZN(new_n828));
  INV_X1    g0628(.A(new_n771), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n829), .A2(G143), .B1(G150), .B2(new_n766), .ZN(new_n830));
  INV_X1    g0630(.A(G137), .ZN(new_n831));
  INV_X1    g0631(.A(new_n776), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n830), .B1(new_n831), .B2(new_n762), .C1(new_n832), .C2(new_n769), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT34), .Z(new_n834));
  INV_X1    g0634(.A(G132), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n290), .B1(new_n780), .B2(new_n217), .C1(new_n835), .C2(new_n774), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n782), .A2(new_n213), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n759), .A2(new_n209), .ZN(new_n838));
  NOR4_X1   g0638(.A1(new_n834), .A2(new_n836), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n769), .ZN(new_n840));
  AOI22_X1  g0640(.A1(G283), .A2(new_n766), .B1(new_n840), .B2(G116), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n546), .B2(new_n762), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(G294), .B2(new_n829), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n786), .A2(G87), .ZN(new_n844));
  INV_X1    g0644(.A(new_n782), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n781), .B1(G107), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n843), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n290), .B(new_n847), .C1(G311), .C2(new_n775), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n756), .B1(new_n839), .B2(new_n848), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n826), .A2(new_n751), .A3(new_n828), .A4(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n825), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n728), .B(new_n851), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(new_n745), .Z(new_n853));
  OAI21_X1  g0653(.A(new_n850), .B1(new_n853), .B2(new_n751), .ZN(G384));
  NOR3_X1   g0654(.A1(new_n233), .A2(new_n202), .A3(new_n385), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(G68), .B2(new_n201), .ZN(new_n856));
  NOR3_X1   g0656(.A1(new_n856), .A2(G13), .A3(new_n273), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT105), .Z(new_n858));
  AOI21_X1  g0658(.A(new_n562), .B1(new_n606), .B2(KEYINPUT35), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n859), .B(new_n230), .C1(KEYINPUT35), .C2(new_n606), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(KEYINPUT36), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT108), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n741), .A2(new_n862), .A3(new_n742), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n739), .B(new_n691), .C1(KEYINPUT108), .C2(KEYINPUT31), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n863), .B(new_n864), .C1(new_n655), .C2(new_n691), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n366), .A2(new_n692), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n368), .A2(new_n373), .A3(new_n867), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n367), .B(new_n691), .C1(new_n358), .C2(new_n372), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n825), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n434), .A2(KEYINPUT16), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n378), .B1(new_n391), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n873), .A2(new_n413), .A3(new_n419), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n437), .A2(KEYINPUT106), .A3(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n689), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT106), .B1(new_n437), .B2(new_n874), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT37), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT37), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n397), .A2(new_n876), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n437), .A2(new_n420), .A3(new_n881), .A4(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n877), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n441), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n884), .A2(KEYINPUT107), .A3(KEYINPUT38), .A4(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT38), .ZN(new_n888));
  AOI221_X4 g0688(.A(new_n888), .B1(new_n441), .B2(new_n885), .C1(new_n880), .C2(new_n883), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT107), .ZN(new_n890));
  INV_X1    g0690(.A(new_n882), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n437), .A2(new_n420), .A3(new_n882), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(KEYINPUT37), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n441), .A2(new_n891), .B1(new_n893), .B2(new_n883), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n890), .B1(new_n894), .B2(KEYINPUT38), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n887), .B1(new_n889), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT40), .B1(new_n871), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n884), .A2(new_n886), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n888), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n884), .A2(KEYINPUT38), .A3(new_n886), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT40), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n865), .A2(new_n901), .A3(new_n902), .A4(new_n870), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n897), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n446), .A2(new_n865), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n904), .B(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(G330), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n424), .A2(new_n876), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n868), .A2(new_n869), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n675), .A2(new_n692), .A3(new_n851), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n910), .B1(new_n911), .B2(new_n822), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n908), .B1(new_n912), .B2(new_n901), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT39), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n914), .B(new_n887), .C1(new_n889), .C2(new_n895), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n899), .A2(KEYINPUT39), .A3(new_n900), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n358), .A2(new_n367), .A3(new_n692), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n915), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n913), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n682), .B1(new_n730), .B2(new_n447), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n920), .B(new_n921), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n907), .A2(new_n922), .B1(new_n273), .B2(new_n685), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT109), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n907), .A2(new_n922), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n858), .B(new_n861), .C1(new_n924), .C2(new_n925), .ZN(G367));
  AOI21_X1  g0726(.A(new_n269), .B1(new_n685), .B2(G45), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT45), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT111), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n663), .A2(new_n691), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n719), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n596), .A2(new_n663), .A3(new_n691), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AND3_X1   g0734(.A1(new_n704), .A2(new_n930), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n930), .B1(new_n704), .B2(new_n934), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n929), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT44), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n704), .B2(new_n719), .ZN(new_n939));
  NOR3_X1   g0739(.A1(new_n525), .A2(new_n530), .A3(new_n448), .ZN(new_n940));
  AOI21_X1  g0740(.A(KEYINPUT94), .B1(new_n535), .B2(new_n538), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n672), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n691), .B1(new_n942), .B2(new_n702), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n943), .A2(KEYINPUT44), .A3(new_n718), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n939), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n934), .ZN(new_n946));
  OAI21_X1  g0746(.A(KEYINPUT111), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n704), .A2(new_n930), .A3(new_n934), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n947), .A2(KEYINPUT45), .A3(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n937), .A2(new_n945), .A3(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n700), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n581), .A2(new_n691), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n540), .A2(new_n696), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n750), .A2(new_n955), .A3(new_n698), .ZN(new_n956));
  AND3_X1   g0756(.A1(new_n700), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n954), .B1(new_n700), .B2(new_n956), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n959), .A2(new_n746), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n937), .A2(new_n949), .A3(new_n700), .A4(new_n945), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n952), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n747), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n707), .B(KEYINPUT41), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n928), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n697), .A2(new_n719), .A3(new_n931), .A4(new_n953), .ZN(new_n966));
  XOR2_X1   g0766(.A(KEYINPUT110), .B(KEYINPUT42), .Z(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n616), .B1(new_n946), .B2(new_n535), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n692), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n966), .A2(new_n968), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n969), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n692), .B1(new_n647), .B2(new_n630), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n659), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n723), .B2(new_n974), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(KEYINPUT43), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n973), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n951), .A2(new_n934), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n973), .A2(new_n979), .A3(new_n977), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n976), .A2(KEYINPUT43), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n981), .A2(new_n984), .A3(new_n982), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n976), .A2(new_n817), .ZN(new_n989));
  INV_X1    g0789(.A(new_n813), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n806), .B1(new_n223), .B2(new_n629), .C1(new_n238), .C2(new_n990), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n782), .A2(new_n217), .B1(new_n774), .B2(new_n831), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT112), .Z(new_n993));
  NAND2_X1  g0793(.A1(new_n763), .A2(G143), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n786), .A2(G77), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n787), .A2(G68), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n766), .A2(new_n776), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n994), .A2(new_n995), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n201), .A2(new_n769), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n290), .B1(new_n771), .B2(new_n262), .ZN(new_n1000));
  NOR4_X1   g0800(.A1(new_n993), .A2(new_n998), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n511), .B1(new_n765), .B2(new_n516), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n845), .A2(G116), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT46), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n829), .A2(G303), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n840), .A2(G283), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n763), .A2(G311), .B1(G107), .B2(new_n787), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1002), .B(new_n1008), .C1(G317), .C2(new_n775), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n786), .A2(new_n622), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1001), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT47), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n751), .B(new_n991), .C1(new_n1012), .C2(new_n757), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n965), .A2(new_n988), .B1(new_n989), .B2(new_n1013), .ZN(G387));
  NOR2_X1   g0814(.A1(new_n959), .A2(new_n927), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT113), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n960), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n959), .A2(new_n746), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1017), .A2(new_n707), .A3(new_n1018), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n375), .A2(new_n766), .B1(G97), .B2(new_n786), .ZN(new_n1020));
  INV_X1    g0820(.A(G159), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1020), .B1(new_n213), .B2(new_n771), .C1(new_n1021), .C2(new_n762), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(new_n327), .B2(new_n787), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n840), .A2(G68), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n845), .A2(G77), .B1(new_n775), .B2(G150), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1023), .A2(new_n290), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n787), .A2(G283), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n829), .A2(G317), .B1(G311), .B2(new_n766), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n546), .B2(new_n769), .C1(new_n799), .C2(new_n762), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT48), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1027), .B1(new_n516), .B2(new_n782), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT115), .Z(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(new_n1030), .B2(new_n1029), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(KEYINPUT49), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n786), .A2(G116), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n775), .A2(G326), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1034), .A2(new_n511), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1033), .A2(KEYINPUT49), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1026), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n752), .B1(new_n1039), .B2(new_n756), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n955), .A2(new_n698), .A3(new_n805), .ZN(new_n1041));
  NOR3_X1   g0841(.A1(new_n324), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1042), .A2(new_n710), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(G68), .A2(G77), .ZN(new_n1044));
  OAI21_X1  g0844(.A(KEYINPUT50), .B1(new_n324), .B2(G50), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1043), .A2(new_n502), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n813), .B(new_n1046), .C1(new_n243), .C2(new_n502), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n710), .A2(new_n223), .A3(new_n290), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1047), .B(new_n1048), .C1(G107), .C2(new_n223), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT114), .Z(new_n1050));
  OAI211_X1 g0850(.A(new_n1040), .B(new_n1041), .C1(new_n807), .C2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1016), .A2(new_n1019), .A3(new_n1051), .ZN(G393));
  NAND2_X1  g0852(.A1(new_n952), .A2(new_n961), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n1017), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1054), .A2(new_n707), .A3(new_n962), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT119), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1053), .A2(new_n927), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n946), .A2(new_n805), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n806), .B1(new_n223), .B2(new_n559), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n250), .B2(new_n813), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n201), .A2(new_n765), .B1(new_n780), .B2(new_n202), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n325), .B2(new_n840), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT117), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n511), .B1(new_n845), .B2(G68), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n775), .A2(G143), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1065), .A2(new_n844), .A3(new_n1066), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT116), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n262), .A2(new_n762), .B1(new_n771), .B2(new_n1021), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT51), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1064), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT118), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n765), .A2(new_n546), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G311), .A2(new_n829), .B1(new_n763), .B2(G317), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT52), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1075), .A2(new_n290), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n769), .A2(new_n516), .B1(new_n774), .B2(new_n799), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n760), .B(new_n1077), .C1(G283), .C2(new_n845), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1076), .B(new_n1078), .C1(new_n562), .C2(new_n780), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1072), .B1(new_n1073), .B2(new_n1079), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n752), .B(new_n1061), .C1(new_n1080), .C2(new_n756), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1058), .B1(new_n1059), .B2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1054), .A2(KEYINPUT119), .A3(new_n707), .A4(new_n962), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1057), .A2(new_n1082), .A3(new_n1083), .ZN(G390));
  NAND3_X1  g0884(.A1(new_n446), .A2(G330), .A3(new_n865), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1085), .B(new_n682), .C1(new_n730), .C2(new_n447), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n821), .B1(new_n726), .B2(new_n824), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n825), .A2(new_n684), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n744), .A2(new_n909), .A3(new_n1089), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n865), .A2(new_n1089), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1088), .B(new_n1090), .C1(new_n1091), .C2(new_n909), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n911), .A2(new_n822), .ZN(new_n1093));
  AND3_X1   g0893(.A1(new_n865), .A2(G330), .A3(new_n870), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n909), .B1(new_n744), .B2(new_n1089), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1093), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1092), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1087), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(KEYINPUT121), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n915), .A2(new_n916), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n912), .B2(new_n918), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT120), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n917), .A2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n358), .A2(KEYINPUT120), .A3(new_n367), .A4(new_n692), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n887), .B(new_n1105), .C1(new_n889), .C2(new_n895), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n1088), .B2(new_n910), .ZN(new_n1108));
  AND3_X1   g0908(.A1(new_n1101), .A2(new_n1108), .A3(new_n1090), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n865), .A2(G330), .A3(new_n870), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n1101), .B2(new_n1108), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1099), .A2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1098), .B(KEYINPUT121), .C1(new_n1109), .C2(new_n1111), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1113), .A2(new_n1114), .A3(new_n707), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n259), .A2(new_n827), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n201), .A2(new_n759), .ZN(new_n1117));
  INV_X1    g0917(.A(G125), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n290), .B1(new_n774), .B2(new_n1118), .C1(new_n831), .C2(new_n765), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n1117), .B(new_n1119), .C1(G159), .C2(new_n787), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n829), .A2(G132), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n782), .A2(new_n262), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT53), .ZN(new_n1123));
  XOR2_X1   g0923(.A(KEYINPUT54), .B(G143), .Z(new_n1124));
  AOI22_X1  g0924(.A1(new_n763), .A2(G128), .B1(new_n840), .B2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1120), .A2(new_n1121), .A3(new_n1123), .A4(new_n1125), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n771), .A2(new_n562), .B1(new_n559), .B2(new_n769), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n783), .B(new_n1127), .C1(G77), .C2(new_n787), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n766), .A2(G107), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n290), .B1(new_n763), .B2(G283), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n759), .A2(new_n209), .B1(new_n774), .B2(new_n516), .ZN(new_n1131));
  XOR2_X1   g0931(.A(new_n1131), .B(KEYINPUT122), .Z(new_n1132));
  NAND4_X1  g0932(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .A4(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n757), .B1(new_n1126), .B2(new_n1133), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n752), .B(new_n1134), .C1(new_n1100), .C2(new_n803), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1112), .A2(new_n928), .B1(new_n1116), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1115), .A2(new_n1136), .ZN(G378));
  INV_X1    g0937(.A(KEYINPUT57), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1086), .B1(new_n1112), .B2(new_n1097), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n904), .A2(G330), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n323), .B1(new_n312), .B2(new_n317), .ZN(new_n1141));
  XOR2_X1   g0941(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1142), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n323), .B(new_n1144), .C1(new_n312), .C2(new_n317), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n284), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1146), .B1(new_n1147), .B2(new_n689), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1143), .A2(new_n284), .A3(new_n876), .A4(new_n1145), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  AND3_X1   g0950(.A1(new_n913), .A2(new_n919), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1150), .B1(new_n913), .B2(new_n919), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1140), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1150), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n920), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n684), .B1(new_n897), .B2(new_n903), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n913), .A2(new_n919), .A3(new_n1150), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1153), .A2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1138), .B1(new_n1139), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1101), .A2(new_n1108), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n1094), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1101), .A2(new_n1108), .A3(new_n1090), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(new_n1097), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n1087), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1165), .A2(KEYINPUT57), .A3(new_n1158), .A4(new_n1153), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1160), .A2(new_n707), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1150), .A2(new_n803), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n827), .A2(new_n201), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(G124), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n252), .B1(new_n774), .B2(new_n1171), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n762), .A2(new_n1118), .B1(new_n835), .B2(new_n765), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1124), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n1174), .A2(new_n782), .B1(new_n262), .B2(new_n780), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1173), .B(new_n1175), .C1(G137), .C2(new_n840), .ZN(new_n1176));
  INV_X1    g0976(.A(G128), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1176), .B1(new_n1177), .B2(new_n771), .ZN(new_n1178));
  AOI211_X1 g0978(.A(G41), .B(new_n1172), .C1(new_n1178), .C2(KEYINPUT59), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1179), .B1(KEYINPUT59), .B2(new_n1178), .C1(new_n759), .C2(new_n832), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n213), .B1(new_n451), .B2(G41), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n996), .B1(new_n771), .B2(new_n460), .C1(new_n562), .C2(new_n762), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(G77), .A2(new_n845), .B1(new_n840), .B2(new_n327), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n601), .B2(new_n765), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1182), .B(new_n1184), .C1(G283), .C2(new_n775), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n786), .A2(G58), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1185), .A2(new_n296), .A3(new_n511), .A4(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT58), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1180), .A2(new_n1181), .A3(new_n1188), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n752), .B(new_n1170), .C1(new_n756), .C2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1159), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1190), .B1(new_n1191), .B2(new_n928), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1167), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT123), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1167), .A2(KEYINPUT123), .A3(new_n1192), .ZN(new_n1196));
  AND2_X1   g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(G375));
  NAND3_X1  g0998(.A1(new_n1086), .A2(new_n1096), .A3(new_n1092), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1098), .A2(new_n964), .A3(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n511), .B1(new_n845), .B2(G159), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1201), .B(new_n1186), .C1(new_n765), .C2(new_n1174), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(G150), .A2(new_n840), .B1(new_n775), .B2(G128), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n835), .B2(new_n762), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n780), .A2(new_n213), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n771), .A2(new_n831), .ZN(new_n1206));
  NOR4_X1   g1006(.A1(new_n1202), .A2(new_n1204), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n829), .A2(G283), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(G116), .A2(new_n766), .B1(new_n775), .B2(G303), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1208), .B(new_n1209), .C1(new_n629), .C2(new_n780), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n995), .B(new_n511), .C1(new_n601), .C2(new_n782), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n769), .A2(new_n460), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n762), .A2(new_n516), .ZN(new_n1213));
  NOR4_X1   g1013(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n756), .B1(new_n1207), .B2(new_n1214), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n751), .B(new_n1215), .C1(new_n909), .C2(new_n804), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n209), .B2(new_n827), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n1097), .B2(new_n928), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1200), .A2(new_n1218), .ZN(G381));
  AND2_X1   g1019(.A1(new_n1115), .A2(new_n1136), .ZN(new_n1220));
  AND3_X1   g1020(.A1(new_n1057), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1221));
  NOR4_X1   g1021(.A1(G393), .A2(G381), .A3(G396), .A4(G384), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1013), .A2(new_n989), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n963), .A2(new_n964), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n927), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n986), .A2(new_n987), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1223), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n1221), .A2(new_n1222), .A3(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1197), .A2(new_n1220), .A3(new_n1228), .ZN(G407));
  NOR2_X1   g1029(.A1(new_n1228), .A2(new_n690), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1195), .A2(new_n1220), .A3(new_n1196), .ZN(new_n1231));
  OAI21_X1  g1031(.A(G213), .B1(new_n1230), .B2(new_n1231), .ZN(G409));
  XNOR2_X1  g1032(.A(G393), .B(G396), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1227), .A2(G390), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1227), .A2(G390), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1233), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(KEYINPUT125), .B1(new_n1227), .B2(G390), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1239), .A2(new_n1236), .ZN(new_n1240));
  XOR2_X1   g1040(.A(G393), .B(G396), .Z(new_n1241));
  INV_X1    g1041(.A(KEYINPUT125), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1241), .B1(new_n1234), .B2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT126), .B1(new_n1240), .B2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1221), .A2(new_n1242), .A3(G387), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1245), .A2(new_n1239), .A3(new_n1233), .A4(new_n1236), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT126), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1238), .B1(new_n1244), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n690), .A2(G213), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1193), .A2(G378), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1191), .A2(new_n964), .A3(new_n1165), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1220), .A2(new_n1192), .A3(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT60), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1098), .B(new_n707), .C1(new_n1254), .C2(new_n1199), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1199), .A2(new_n1254), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1218), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1257), .B(G384), .ZN(new_n1258));
  AND4_X1   g1058(.A1(new_n1250), .A2(new_n1251), .A3(new_n1253), .A4(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT61), .B1(new_n1259), .B2(KEYINPUT63), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT63), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1251), .A2(new_n1253), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(KEYINPUT124), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT124), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1251), .A2(new_n1264), .A3(new_n1253), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1263), .A2(new_n1250), .A3(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n690), .A2(G213), .A3(G2897), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1258), .B(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1261), .B1(new_n1266), .B2(new_n1269), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1263), .A2(new_n1250), .A3(new_n1258), .A4(new_n1265), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1249), .B(new_n1260), .C1(new_n1270), .C2(new_n1272), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n1271), .A2(new_n1274), .B1(KEYINPUT62), .B2(new_n1259), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT61), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1262), .B1(G213), .B2(new_n690), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1276), .B1(new_n1277), .B2(new_n1268), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1275), .A2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1273), .B1(new_n1279), .B2(new_n1249), .ZN(G405));
  INV_X1    g1080(.A(new_n1258), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1243), .A2(KEYINPUT126), .A3(new_n1236), .A4(new_n1239), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1283));
  AOI221_X4 g1083(.A(new_n1237), .B1(new_n1231), .B2(new_n1251), .C1(new_n1282), .C2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1231), .A2(new_n1251), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1285), .B1(new_n1286), .B2(new_n1238), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1281), .B1(new_n1284), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1285), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1249), .A2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1286), .A2(new_n1238), .A3(new_n1285), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1290), .A2(new_n1258), .A3(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1288), .A2(new_n1292), .ZN(G402));
endmodule


