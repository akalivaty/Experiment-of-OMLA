//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 0 1 0 0 1 0 1 0 1 1 1 1 0 1 1 0 1 0 1 1 1 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n839, new_n840, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202));
  INV_X1    g001(.A(G71gat), .ZN(new_n203));
  INV_X1    g002(.A(G78gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g005(.A1(G71gat), .A2(G78gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT9), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n202), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT9), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n206), .B1(new_n202), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT94), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n207), .A2(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT94), .B1(G71gat), .B2(G78gat), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NOR3_X1   g015(.A1(new_n212), .A2(new_n216), .A3(KEYINPUT95), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT95), .ZN(new_n218));
  INV_X1    g017(.A(G64gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G57gat), .ZN(new_n220));
  INV_X1    g019(.A(G57gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G64gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n205), .B1(new_n223), .B2(KEYINPUT9), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n214), .A2(new_n215), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n218), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n210), .B1(new_n217), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT96), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT95), .B1(new_n212), .B2(new_n216), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n224), .A2(new_n218), .A3(new_n225), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n209), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT96), .ZN(new_n233));
  NAND2_X1  g032(.A1(G99gat), .A2(G106gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT99), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(KEYINPUT99), .A2(G99gat), .A3(G106gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(KEYINPUT8), .A3(new_n237), .ZN(new_n238));
  AND2_X1   g037(.A1(G85gat), .A2(G92gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT98), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n239), .A2(KEYINPUT97), .A3(new_n240), .A4(KEYINPUT7), .ZN(new_n241));
  INV_X1    g040(.A(G85gat), .ZN(new_n242));
  INV_X1    g041(.A(G92gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(G85gat), .A2(G92gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(KEYINPUT97), .A2(KEYINPUT7), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT7), .ZN(new_n247));
  AOI22_X1  g046(.A1(new_n245), .A2(new_n246), .B1(new_n247), .B2(KEYINPUT98), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n238), .A2(new_n241), .A3(new_n244), .A4(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G99gat), .B(G106gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n229), .A2(new_n233), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT10), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n251), .A2(new_n232), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT101), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT101), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n251), .A2(new_n232), .A3(new_n257), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n253), .A2(new_n254), .A3(new_n256), .A4(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT102), .ZN(new_n260));
  INV_X1    g059(.A(new_n258), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n257), .B1(new_n251), .B2(new_n232), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT102), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n263), .A2(new_n264), .A3(new_n254), .A4(new_n253), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n260), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n229), .A2(new_n233), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n267), .A2(KEYINPUT10), .A3(new_n251), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G230gat), .A2(G233gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n263), .A2(new_n253), .ZN(new_n272));
  INV_X1    g071(.A(new_n270), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G120gat), .B(G148gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(G176gat), .B(G204gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n271), .A2(new_n274), .A3(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n268), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n280), .B1(new_n260), .B2(new_n265), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n274), .B1(new_n281), .B2(new_n273), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(new_n277), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT27), .B(G183gat), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT28), .B1(new_n286), .B2(G190gat), .ZN(new_n287));
  INV_X1    g086(.A(G169gat), .ZN(new_n288));
  INV_X1    g087(.A(G176gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT26), .ZN(new_n291));
  OR3_X1    g090(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n291), .B(new_n292), .C1(new_n288), .C2(new_n289), .ZN(new_n293));
  NAND2_X1  g092(.A1(G183gat), .A2(G190gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT28), .ZN(new_n295));
  INV_X1    g094(.A(G190gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n285), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n287), .A2(new_n293), .A3(new_n294), .A4(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT24), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(G183gat), .A2(G190gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n294), .A2(new_n299), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  XOR2_X1   g103(.A(KEYINPUT64), .B(G169gat), .Z(new_n305));
  NAND3_X1  g104(.A1(new_n305), .A2(KEYINPUT23), .A3(new_n289), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT25), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT23), .B1(new_n288), .B2(new_n289), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(new_n290), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n304), .A2(new_n306), .A3(new_n307), .A4(new_n309), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n298), .A2(new_n310), .ZN(new_n311));
  AND2_X1   g110(.A1(KEYINPUT65), .A2(KEYINPUT24), .ZN(new_n312));
  NOR2_X1   g111(.A1(KEYINPUT65), .A2(KEYINPUT24), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n294), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT66), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI211_X1 g115(.A(KEYINPUT66), .B(new_n294), .C1(new_n312), .C2(new_n313), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(new_n302), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT23), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n318), .B(new_n309), .C1(new_n319), .C2(new_n290), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT25), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n311), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G113gat), .B(G120gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n323), .A2(KEYINPUT1), .ZN(new_n324));
  XOR2_X1   g123(.A(G127gat), .B(G134gat), .Z(new_n325));
  XNOR2_X1  g124(.A(new_n324), .B(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n322), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G227gat), .ZN(new_n329));
  INV_X1    g128(.A(G233gat), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n311), .A2(new_n321), .A3(new_n326), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n328), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT70), .ZN(new_n335));
  AND3_X1   g134(.A1(new_n334), .A2(new_n335), .A3(KEYINPUT34), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n335), .B1(new_n334), .B2(KEYINPUT34), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n334), .A2(KEYINPUT34), .ZN(new_n338));
  NOR3_X1   g137(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G15gat), .B(G43gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n341), .B(G99gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT68), .B(G71gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n342), .B(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n333), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n326), .B1(new_n311), .B2(new_n321), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n331), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT67), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI211_X1 g149(.A(KEYINPUT67), .B(new_n331), .C1(new_n346), .C2(new_n347), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT32), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT33), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n345), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n345), .A2(KEYINPUT69), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT69), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT33), .B1(new_n344), .B2(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  AOI211_X1 g158(.A(new_n353), .B(new_n359), .C1(new_n350), .C2(new_n351), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n340), .B1(new_n355), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n351), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n328), .A2(new_n333), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT67), .B1(new_n363), .B2(new_n331), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n354), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n344), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n352), .B(KEYINPUT32), .C1(new_n356), .C2(new_n358), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n366), .A2(new_n367), .A3(new_n339), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n361), .A2(KEYINPUT71), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT71), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n340), .B(new_n370), .C1(new_n355), .C2(new_n360), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(G8gat), .B(G36gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(G64gat), .B(G92gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  XOR2_X1   g174(.A(G197gat), .B(G204gat), .Z(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT73), .B(G211gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(G218gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(KEYINPUT72), .B(KEYINPUT22), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n376), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT74), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT74), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(G211gat), .B(G218gat), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n382), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n384), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n385), .B1(new_n380), .B2(new_n383), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(G226gat), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n391), .A2(new_n330), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n322), .A2(KEYINPUT75), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT75), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n311), .A2(new_n321), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n393), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n392), .A2(KEYINPUT29), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n322), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n390), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT76), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n394), .A2(new_n396), .A3(new_n398), .ZN(new_n403));
  INV_X1    g202(.A(new_n390), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n311), .A2(new_n321), .A3(new_n392), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n401), .A2(new_n402), .A3(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n402), .B1(new_n401), .B2(new_n406), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n375), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n401), .A2(new_n406), .ZN(new_n411));
  INV_X1    g210(.A(new_n375), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT30), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n403), .A2(new_n405), .A3(new_n404), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n311), .A2(new_n321), .A3(new_n395), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n395), .B1(new_n311), .B2(new_n321), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n392), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n404), .B1(new_n419), .B2(new_n399), .ZN(new_n420));
  OAI211_X1 g219(.A(KEYINPUT30), .B(new_n412), .C1(new_n416), .C2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT77), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n411), .A2(KEYINPUT77), .A3(KEYINPUT30), .A4(new_n412), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n410), .A2(new_n415), .A3(new_n423), .A4(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT85), .ZN(new_n427));
  NAND2_X1  g226(.A1(G225gat), .A2(G233gat), .ZN(new_n428));
  XNOR2_X1  g227(.A(G155gat), .B(G162gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(G141gat), .B(G148gat), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT2), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n429), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n429), .ZN(new_n434));
  XOR2_X1   g233(.A(KEYINPUT80), .B(G155gat), .Z(new_n435));
  XNOR2_X1  g234(.A(KEYINPUT81), .B(G162gat), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n434), .B1(new_n437), .B2(KEYINPUT2), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n430), .B(KEYINPUT79), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n433), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n441), .A2(new_n327), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT4), .ZN(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT82), .B(KEYINPUT4), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT3), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n438), .A2(new_n439), .ZN(new_n446));
  INV_X1    g245(.A(new_n433), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AOI211_X1 g247(.A(KEYINPUT3), .B(new_n433), .C1(new_n438), .C2(new_n439), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n444), .B1(new_n450), .B2(new_n327), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n428), .B(new_n443), .C1(new_n451), .C2(new_n442), .ZN(new_n452));
  INV_X1    g251(.A(new_n442), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n441), .A2(new_n327), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n455), .A2(G225gat), .A3(G233gat), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n452), .A2(KEYINPUT5), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n448), .ZN(new_n458));
  INV_X1    g257(.A(new_n449), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n458), .A2(new_n459), .A3(new_n327), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n460), .A2(KEYINPUT4), .A3(new_n453), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n442), .A2(new_n444), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT5), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n463), .A2(new_n464), .A3(new_n428), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n457), .A2(new_n465), .ZN(new_n466));
  XOR2_X1   g265(.A(G57gat), .B(G85gat), .Z(new_n467));
  XNOR2_X1  g266(.A(G1gat), .B(G29gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n467), .B(new_n468), .ZN(new_n469));
  XOR2_X1   g268(.A(KEYINPUT83), .B(KEYINPUT0), .Z(new_n470));
  XNOR2_X1  g269(.A(new_n470), .B(KEYINPUT84), .ZN(new_n471));
  XOR2_X1   g270(.A(new_n469), .B(new_n471), .Z(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n466), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT6), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n427), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n472), .B1(new_n457), .B2(new_n465), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n477), .A2(KEYINPUT85), .A3(KEYINPUT6), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n457), .A2(new_n472), .A3(new_n465), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n474), .A2(new_n475), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n476), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT29), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n386), .A2(new_n389), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n445), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(new_n441), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n459), .A2(new_n482), .B1(new_n389), .B2(new_n386), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(G228gat), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n488), .A2(new_n330), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT86), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT86), .B1(new_n488), .B2(new_n330), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n485), .A2(new_n487), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n440), .B1(new_n483), .B2(new_n445), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n490), .B(new_n489), .C1(new_n494), .C2(new_n486), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(new_n495), .A3(G22gat), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT87), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(G78gat), .B(G106gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n499), .B(KEYINPUT31), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(G50gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n493), .A2(new_n495), .ZN(new_n503));
  INV_X1    g302(.A(G22gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n496), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n505), .A2(KEYINPUT87), .A3(new_n496), .A4(new_n501), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT35), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n372), .A2(new_n426), .A3(new_n481), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT88), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n425), .B1(new_n369), .B2(new_n371), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT88), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n512), .A2(new_n513), .A3(new_n481), .A4(new_n509), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT78), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n423), .A2(new_n424), .ZN(new_n516));
  INV_X1    g315(.A(new_n409), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n412), .B1(new_n517), .B2(new_n407), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n515), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n410), .A2(KEYINPUT78), .A3(new_n423), .A4(new_n424), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n481), .A2(new_n519), .A3(new_n415), .A4(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n361), .A2(new_n368), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n508), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NOR3_X1   g323(.A1(new_n521), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT35), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n511), .B(new_n514), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n463), .A2(new_n428), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n453), .A2(new_n428), .A3(new_n454), .ZN(new_n529));
  AND3_X1   g328(.A1(new_n528), .A2(KEYINPUT39), .A3(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n472), .B1(new_n528), .B2(KEYINPUT39), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT40), .ZN(new_n532));
  OR3_X1    g331(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n532), .B1(new_n530), .B2(new_n531), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n533), .A2(new_n425), .A3(new_n474), .A4(new_n534), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n477), .A2(KEYINPUT85), .A3(KEYINPUT6), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT85), .B1(new_n477), .B2(KEYINPUT6), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n404), .B1(new_n397), .B2(new_n400), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n403), .A2(new_n390), .A3(new_n405), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n539), .A2(KEYINPUT37), .A3(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n541), .B1(new_n411), .B2(KEYINPUT37), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT38), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n542), .A2(new_n543), .A3(new_n375), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n538), .A2(new_n480), .A3(new_n413), .A4(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n517), .A2(KEYINPUT37), .A3(new_n407), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n546), .B1(KEYINPUT37), .B2(new_n411), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n543), .B1(new_n547), .B2(new_n375), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n523), .B(new_n535), .C1(new_n545), .C2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n521), .A2(new_n524), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT36), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n551), .B1(new_n361), .B2(new_n368), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n552), .B1(new_n372), .B2(new_n551), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n549), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n284), .B1(new_n527), .B2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G127gat), .B(G155gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(G211gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n267), .A2(KEYINPUT21), .ZN(new_n558));
  XNOR2_X1  g357(.A(G15gat), .B(G22gat), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT16), .ZN(new_n560));
  AOI21_X1  g359(.A(G1gat), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(G8gat), .ZN(new_n562));
  OR2_X1    g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n559), .A2(KEYINPUT92), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n561), .A2(new_n562), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n563), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n565), .B1(new_n563), .B2(new_n566), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n558), .A2(new_n571), .ZN(new_n572));
  OR2_X1    g371(.A1(new_n572), .A2(G183gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(G183gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n267), .A2(KEYINPUT21), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G231gat), .A2(G233gat), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n573), .B(new_n574), .C1(KEYINPUT21), .C2(new_n267), .ZN(new_n580));
  AND3_X1   g379(.A1(new_n577), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n579), .B1(new_n577), .B2(new_n580), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n557), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n577), .A2(new_n580), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(new_n578), .ZN(new_n585));
  INV_X1    g384(.A(new_n557), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n577), .A2(new_n579), .A3(new_n580), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n583), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n589), .B1(new_n583), .B2(new_n588), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(G29gat), .ZN(new_n594));
  INV_X1    g393(.A(G36gat), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n594), .A2(new_n595), .A3(KEYINPUT14), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT14), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n597), .B1(G29gat), .B2(G36gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(G29gat), .A2(G36gat), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n596), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G43gat), .B(G50gat), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n600), .A2(KEYINPUT15), .A3(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT89), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n600), .A2(KEYINPUT89), .A3(KEYINPUT15), .A4(new_n601), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(G43gat), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT90), .B1(new_n607), .B2(G50gat), .ZN(new_n608));
  OR3_X1    g407(.A1(new_n601), .A2(KEYINPUT15), .A3(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n600), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n601), .B1(KEYINPUT15), .B2(new_n608), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n606), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(KEYINPUT91), .A2(KEYINPUT17), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT91), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT17), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n613), .A2(new_n614), .A3(new_n617), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n606), .A2(new_n612), .A3(new_n615), .A4(new_n616), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n570), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n569), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n621), .A2(new_n613), .A3(new_n567), .ZN(new_n622));
  NAND2_X1  g421(.A1(G229gat), .A2(G233gat), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NOR3_X1   g423(.A1(new_n620), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(KEYINPUT18), .B1(new_n625), .B2(KEYINPUT93), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n570), .B(new_n613), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n623), .B(KEYINPUT13), .Z(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n618), .A2(new_n619), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n571), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n622), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n631), .A2(new_n632), .A3(new_n623), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT93), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT18), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n626), .A2(new_n629), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G113gat), .B(G141gat), .ZN(new_n638));
  INV_X1    g437(.A(G197gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT11), .B(G169gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT12), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n637), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n626), .A2(new_n643), .A3(new_n629), .A4(new_n636), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  AND2_X1   g447(.A1(G232gat), .A2(G233gat), .ZN(new_n649));
  AOI22_X1  g448(.A1(new_n630), .A2(new_n252), .B1(KEYINPUT41), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n613), .A2(new_n251), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g451(.A(G190gat), .B(G218gat), .Z(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n650), .A2(new_n653), .A3(new_n651), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n649), .A2(KEYINPUT41), .ZN(new_n658));
  XNOR2_X1  g457(.A(G134gat), .B(G162gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n657), .A2(KEYINPUT100), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(KEYINPUT100), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n663), .B(new_n656), .C1(new_n655), .C2(new_n661), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n593), .A2(new_n648), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n555), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n667), .A2(new_n481), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT103), .B(G1gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(G1324gat));
  INV_X1    g469(.A(new_n667), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n425), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(G8gat), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(KEYINPUT42), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT104), .B(KEYINPUT16), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(G8gat), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  MUX2_X1   g476(.A(new_n674), .B(KEYINPUT42), .S(new_n677), .Z(G1325gat));
  INV_X1    g477(.A(new_n553), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n671), .A2(G15gat), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(G15gat), .B1(new_n671), .B2(new_n372), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n680), .A2(new_n681), .ZN(G1326gat));
  NAND2_X1  g481(.A1(new_n671), .A2(new_n524), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(G22gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1327gat));
  INV_X1    g485(.A(new_n665), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n687), .B1(new_n527), .B2(new_n554), .ZN(new_n688));
  INV_X1    g487(.A(new_n284), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n593), .A2(new_n689), .A3(new_n647), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n481), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n693), .A2(new_n594), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT45), .ZN(new_n696));
  AOI211_X1 g495(.A(KEYINPUT44), .B(new_n687), .C1(new_n527), .C2(new_n554), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n521), .A2(new_n524), .ZN(new_n699));
  INV_X1    g498(.A(new_n522), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n526), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n511), .A2(new_n514), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n554), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n698), .B1(new_n703), .B2(new_n665), .ZN(new_n704));
  OR2_X1    g503(.A1(new_n697), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(new_n691), .ZN(new_n706));
  OAI21_X1  g505(.A(G29gat), .B1(new_n706), .B2(new_n481), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n696), .A2(new_n707), .ZN(G1328gat));
  NOR3_X1   g507(.A1(new_n692), .A2(G36gat), .A3(new_n426), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT46), .ZN(new_n710));
  OAI21_X1  g509(.A(G36gat), .B1(new_n706), .B2(new_n426), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(G1329gat));
  AND3_X1   g511(.A1(new_n693), .A2(new_n607), .A3(new_n372), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n705), .A2(new_n679), .A3(new_n691), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n713), .B1(new_n714), .B2(G43gat), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT47), .ZN(G1330gat));
  OR2_X1    g515(.A1(new_n692), .A2(KEYINPUT106), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n692), .A2(KEYINPUT106), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n717), .A2(new_n524), .A3(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(G50gat), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n524), .A2(G50gat), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n721), .B1(new_n706), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(KEYINPUT48), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT48), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n721), .B(new_n725), .C1(new_n706), .C2(new_n722), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(G1331gat));
  NAND2_X1  g526(.A1(new_n583), .A2(new_n588), .ZN(new_n728));
  INV_X1    g527(.A(new_n589), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n583), .A2(new_n588), .A3(new_n589), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n730), .A2(new_n648), .A3(new_n731), .A4(new_n687), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n732), .B1(new_n527), .B2(new_n554), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n284), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n734), .A2(new_n481), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(new_n221), .ZN(G1332gat));
  AOI21_X1  g535(.A(new_n426), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n737));
  XOR2_X1   g536(.A(new_n737), .B(KEYINPUT107), .Z(new_n738));
  NAND3_X1  g537(.A1(new_n733), .A2(new_n284), .A3(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  XOR2_X1   g539(.A(new_n739), .B(new_n740), .Z(G1333gat));
  OAI21_X1  g540(.A(G71gat), .B1(new_n734), .B2(new_n553), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n733), .A2(new_n203), .A3(new_n284), .A4(new_n372), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT108), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT108), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n742), .A2(new_n746), .A3(new_n743), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g548(.A1(new_n734), .A2(new_n523), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(new_n204), .ZN(G1335gat));
  NOR2_X1   g550(.A1(new_n592), .A2(new_n647), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n284), .B(new_n752), .C1(new_n697), .C2(new_n704), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n481), .A2(new_n242), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT109), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n703), .A2(new_n665), .ZN(new_n758));
  INV_X1    g557(.A(new_n752), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n757), .B(KEYINPUT51), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n757), .A2(KEYINPUT51), .ZN(new_n761));
  OR2_X1    g560(.A1(new_n757), .A2(KEYINPUT51), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n688), .A2(new_n761), .A3(new_n752), .A4(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n760), .A2(new_n694), .A3(new_n284), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n242), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n756), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n766), .B(new_n767), .ZN(G1336gat));
  AOI21_X1  g567(.A(new_n243), .B1(new_n754), .B2(new_n425), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n760), .A2(new_n243), .A3(new_n284), .A4(new_n763), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n770), .A2(new_n426), .ZN(new_n771));
  OAI21_X1  g570(.A(KEYINPUT52), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n773), .B1(new_n754), .B2(new_n425), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n753), .A2(KEYINPUT111), .A3(new_n426), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n774), .A2(new_n243), .A3(new_n775), .ZN(new_n776));
  OR2_X1    g575(.A1(new_n771), .A2(KEYINPUT52), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n772), .B1(new_n776), .B2(new_n777), .ZN(G1337gat));
  OAI21_X1  g577(.A(G99gat), .B1(new_n753), .B2(new_n553), .ZN(new_n779));
  AOI21_X1  g578(.A(G99gat), .B1(new_n369), .B2(new_n371), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n760), .A2(new_n284), .A3(new_n763), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n779), .A2(new_n781), .ZN(G1338gat));
  NOR2_X1   g581(.A1(new_n523), .A2(G106gat), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n760), .A2(new_n284), .A3(new_n763), .A4(new_n783), .ZN(new_n784));
  OR2_X1    g583(.A1(new_n784), .A2(KEYINPUT114), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n786));
  XNOR2_X1  g585(.A(KEYINPUT112), .B(G106gat), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n787), .B1(new_n753), .B2(new_n523), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n784), .A2(KEYINPUT114), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n785), .A2(new_n786), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n784), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT113), .B1(new_n791), .B2(KEYINPUT53), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT113), .ZN(new_n793));
  AOI211_X1 g592(.A(new_n793), .B(new_n786), .C1(new_n788), .C2(new_n784), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n790), .B1(new_n792), .B2(new_n794), .ZN(G1339gat));
  NOR2_X1   g594(.A1(new_n732), .A2(new_n284), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n627), .A2(new_n628), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n623), .B1(new_n631), .B2(new_n632), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n642), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n284), .A2(new_n646), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n801), .B1(new_n281), .B2(new_n273), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n271), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n273), .B1(new_n266), .B2(new_n268), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n278), .B1(new_n804), .B2(new_n801), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n803), .A2(new_n805), .A3(KEYINPUT55), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n806), .A2(new_n279), .A3(new_n647), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT55), .B1(new_n803), .B2(new_n805), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n800), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n806), .A2(new_n279), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n810), .A2(new_n808), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n646), .A2(new_n799), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n687), .A2(new_n812), .ZN(new_n813));
  AOI22_X1  g612(.A1(new_n809), .A2(new_n687), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n592), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817));
  AOI211_X1 g616(.A(new_n270), .B(new_n280), .C1(new_n260), .C2(new_n265), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n804), .A2(new_n818), .A3(new_n801), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n269), .A2(new_n801), .A3(new_n270), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n277), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n817), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n822), .A2(new_n279), .A3(new_n647), .A4(new_n806), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n665), .B1(new_n823), .B2(new_n800), .ZN(new_n824));
  NOR4_X1   g623(.A1(new_n810), .A2(new_n808), .A3(new_n687), .A4(new_n812), .ZN(new_n825));
  OAI21_X1  g624(.A(KEYINPUT115), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n796), .B1(new_n816), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n827), .A2(new_n524), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n828), .A2(new_n694), .A3(new_n512), .ZN(new_n829));
  OAI21_X1  g628(.A(G113gat), .B1(new_n829), .B2(new_n648), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n827), .A2(new_n524), .A3(new_n522), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n481), .A2(new_n425), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n648), .A2(G113gat), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n830), .B1(new_n833), .B2(new_n834), .ZN(G1340gat));
  OAI21_X1  g634(.A(G120gat), .B1(new_n829), .B2(new_n689), .ZN(new_n836));
  OR2_X1    g635(.A1(new_n689), .A2(G120gat), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n836), .B1(new_n833), .B2(new_n837), .ZN(G1341gat));
  INV_X1    g637(.A(G127gat), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n829), .A2(new_n839), .A3(new_n593), .ZN(new_n840));
  INV_X1    g639(.A(new_n833), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n592), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n840), .B1(new_n842), .B2(new_n839), .ZN(G1342gat));
  OR3_X1    g642(.A1(new_n833), .A2(G134gat), .A3(new_n687), .ZN(new_n844));
  OR2_X1    g643(.A1(new_n844), .A2(KEYINPUT56), .ZN(new_n845));
  OAI21_X1  g644(.A(G134gat), .B1(new_n829), .B2(new_n687), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n844), .A2(KEYINPUT56), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(G1343gat));
  INV_X1    g647(.A(KEYINPUT117), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n809), .A2(new_n687), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n811), .A2(new_n813), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n850), .A2(new_n815), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n826), .A2(new_n852), .A3(new_n593), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n732), .A2(new_n284), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n523), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  XOR2_X1   g654(.A(KEYINPUT116), .B(KEYINPUT57), .Z(new_n856));
  OAI21_X1  g655(.A(new_n849), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n807), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT118), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n859), .B1(new_n819), .B2(new_n821), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n803), .A2(new_n805), .A3(KEYINPUT118), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(new_n817), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n858), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n800), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n825), .B1(new_n864), .B2(new_n687), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n854), .B1(new_n865), .B2(new_n592), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(KEYINPUT57), .A3(new_n524), .ZN(new_n867));
  INV_X1    g666(.A(new_n856), .ZN(new_n868));
  OAI211_X1 g667(.A(KEYINPUT117), .B(new_n868), .C1(new_n827), .C2(new_n523), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n857), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n553), .A2(new_n832), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n870), .A2(new_n647), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(G141gat), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n853), .A2(new_n854), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n524), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n876), .A2(new_n871), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  OR3_X1    g677(.A1(new_n878), .A2(G141gat), .A3(new_n648), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n874), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT58), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT58), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n874), .A2(new_n882), .A3(new_n879), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n881), .A2(new_n883), .ZN(G1344gat));
  XNOR2_X1  g683(.A(new_n871), .B(KEYINPUT121), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n876), .A2(new_n868), .ZN(new_n886));
  AOI21_X1  g685(.A(KEYINPUT57), .B1(new_n866), .B2(new_n524), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n284), .B(new_n885), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n888), .A2(G148gat), .ZN(new_n889));
  XNOR2_X1  g688(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n870), .A2(new_n284), .A3(new_n872), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(G148gat), .ZN(new_n892));
  OAI22_X1  g691(.A1(new_n889), .A2(new_n890), .B1(new_n892), .B2(KEYINPUT59), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n878), .A2(G148gat), .A3(new_n689), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(KEYINPUT119), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(new_n895), .ZN(G1345gat));
  AOI21_X1  g695(.A(new_n435), .B1(new_n877), .B2(new_n592), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n870), .A2(new_n872), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n592), .A2(new_n435), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n899), .B(KEYINPUT122), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n897), .B1(new_n898), .B2(new_n900), .ZN(G1346gat));
  AOI21_X1  g700(.A(new_n436), .B1(new_n877), .B2(new_n665), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n665), .A2(new_n436), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(new_n898), .B2(new_n903), .ZN(G1347gat));
  NOR2_X1   g703(.A1(new_n694), .A2(new_n426), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n905), .A2(new_n372), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n906), .A2(KEYINPUT123), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(KEYINPUT123), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n828), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(G169gat), .B1(new_n909), .B2(new_n648), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n831), .A2(new_n905), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n647), .A2(new_n305), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(G1348gat));
  NOR3_X1   g712(.A1(new_n909), .A2(new_n289), .A3(new_n689), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n831), .A2(new_n284), .A3(new_n905), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n914), .B1(new_n289), .B2(new_n915), .ZN(G1349gat));
  OAI21_X1  g715(.A(G183gat), .B1(new_n909), .B2(new_n593), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n592), .A2(new_n285), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n911), .B2(new_n918), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT60), .ZN(G1350gat));
  NAND4_X1  g719(.A1(new_n828), .A2(new_n665), .A3(new_n907), .A4(new_n908), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT61), .ZN(new_n922));
  AND3_X1   g721(.A1(new_n921), .A2(new_n922), .A3(G190gat), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n922), .B1(new_n921), .B2(G190gat), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n665), .A2(new_n296), .ZN(new_n925));
  OAI22_X1  g724(.A1(new_n923), .A2(new_n924), .B1(new_n911), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(KEYINPUT124), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT124), .ZN(new_n928));
  OAI221_X1 g727(.A(new_n928), .B1(new_n911), .B2(new_n925), .C1(new_n923), .C2(new_n924), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(G1351gat));
  AND2_X1   g729(.A1(new_n866), .A2(new_n524), .ZN(new_n931));
  OAI22_X1  g730(.A1(new_n931), .A2(KEYINPUT57), .B1(new_n876), .B2(new_n868), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n553), .A2(new_n905), .ZN(new_n933));
  XOR2_X1   g732(.A(new_n933), .B(KEYINPUT125), .Z(new_n934));
  NAND3_X1  g733(.A1(new_n932), .A2(new_n647), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(KEYINPUT126), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT126), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n932), .A2(new_n937), .A3(new_n647), .A4(new_n934), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n936), .A2(G197gat), .A3(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(new_n933), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n855), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n647), .A2(new_n639), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(G1352gat));
  NOR3_X1   g742(.A1(new_n941), .A2(G204gat), .A3(new_n689), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT62), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n886), .A2(new_n887), .ZN(new_n946));
  INV_X1    g745(.A(new_n934), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n946), .A2(new_n689), .A3(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(G204gat), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(G1353gat));
  OR3_X1    g749(.A1(new_n941), .A2(new_n377), .A3(new_n593), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n932), .A2(new_n592), .A3(new_n940), .ZN(new_n952));
  AND3_X1   g751(.A1(new_n952), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n953));
  AOI21_X1  g752(.A(KEYINPUT63), .B1(new_n952), .B2(G211gat), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n951), .B1(new_n953), .B2(new_n954), .ZN(G1354gat));
  INV_X1    g754(.A(KEYINPUT127), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n956), .B1(new_n946), .B2(new_n947), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n932), .A2(KEYINPUT127), .A3(new_n934), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n957), .A2(new_n665), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(G218gat), .ZN(new_n960));
  OR3_X1    g759(.A1(new_n941), .A2(G218gat), .A3(new_n687), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(G1355gat));
endmodule


