

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U555 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U556 ( .A1(n706), .A2(n969), .ZN(n687) );
  INV_X1 U557 ( .A(KEYINPUT28), .ZN(n523) );
  NOR2_X1 U558 ( .A1(n624), .A2(n623), .ZN(n654) );
  XNOR2_X1 U559 ( .A(n622), .B(KEYINPUT27), .ZN(n624) );
  NOR2_X1 U560 ( .A1(n591), .A2(G651), .ZN(n802) );
  XNOR2_X1 U561 ( .A(n521), .B(KEYINPUT23), .ZN(n540) );
  XNOR2_X1 U562 ( .A(n536), .B(n535), .ZN(n551) );
  NAND2_X1 U563 ( .A1(n534), .A2(G2104), .ZN(n536) );
  NAND2_X1 U564 ( .A1(n551), .A2(G101), .ZN(n521) );
  NAND2_X1 U565 ( .A1(n657), .A2(n522), .ZN(n659) );
  XNOR2_X1 U566 ( .A(n625), .B(n523), .ZN(n522) );
  NOR2_X2 U567 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X2 U568 ( .A1(G2105), .A2(G2104), .ZN(n542) );
  NOR2_X2 U569 ( .A1(G543), .A2(G651), .ZN(n796) );
  BUF_X1 U570 ( .A(n721), .Z(n524) );
  XNOR2_X1 U571 ( .A(n538), .B(KEYINPUT65), .ZN(n721) );
  OR2_X1 U572 ( .A1(n650), .A2(n649), .ZN(n653) );
  AND2_X1 U573 ( .A1(n638), .A2(n637), .ZN(n650) );
  AND2_X2 U574 ( .A1(G2104), .A2(G2105), .ZN(n884) );
  AND2_X1 U575 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U576 ( .A1(n646), .A2(G1961), .ZN(n610) );
  AND2_X1 U577 ( .A1(n694), .A2(n711), .ZN(n695) );
  XNOR2_X1 U578 ( .A(n542), .B(n541), .ZN(n550) );
  INV_X1 U579 ( .A(KEYINPUT17), .ZN(n541) );
  INV_X1 U580 ( .A(n688), .ZN(n667) );
  AND2_X1 U581 ( .A1(n636), .A2(n770), .ZN(n637) );
  NOR2_X1 U582 ( .A1(G171), .A2(n660), .ZN(n620) );
  NAND2_X1 U583 ( .A1(n614), .A2(G8), .ZN(n615) );
  XNOR2_X1 U584 ( .A(n615), .B(KEYINPUT93), .ZN(n688) );
  BUF_X1 U585 ( .A(n688), .Z(n711) );
  NAND2_X1 U586 ( .A1(n550), .A2(G137), .ZN(n545) );
  INV_X1 U587 ( .A(KEYINPUT66), .ZN(n535) );
  NOR2_X2 U588 ( .A1(n591), .A2(n528), .ZN(n797) );
  BUF_X1 U589 ( .A(n550), .Z(n879) );
  XNOR2_X1 U590 ( .A(n549), .B(KEYINPUT64), .ZN(n608) );
  BUF_X1 U591 ( .A(n608), .Z(G160) );
  INV_X1 U592 ( .A(G651), .ZN(n528) );
  NOR2_X1 U593 ( .A1(G543), .A2(n528), .ZN(n525) );
  XOR2_X2 U594 ( .A(KEYINPUT1), .B(n525), .Z(n801) );
  NAND2_X1 U595 ( .A1(G64), .A2(n801), .ZN(n527) );
  XOR2_X1 U596 ( .A(KEYINPUT0), .B(G543), .Z(n591) );
  NAND2_X1 U597 ( .A1(G52), .A2(n802), .ZN(n526) );
  NAND2_X1 U598 ( .A1(n527), .A2(n526), .ZN(n533) );
  NAND2_X1 U599 ( .A1(G90), .A2(n796), .ZN(n530) );
  NAND2_X1 U600 ( .A1(G77), .A2(n797), .ZN(n529) );
  NAND2_X1 U601 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U602 ( .A(KEYINPUT9), .B(n531), .Z(n532) );
  NOR2_X1 U603 ( .A1(n533), .A2(n532), .ZN(G171) );
  INV_X1 U604 ( .A(G2105), .ZN(n534) );
  INV_X1 U605 ( .A(G2104), .ZN(n543) );
  NAND2_X1 U606 ( .A1(n543), .A2(G2105), .ZN(n538) );
  AND2_X1 U607 ( .A1(G125), .A2(n721), .ZN(n539) );
  NOR2_X1 U608 ( .A1(n540), .A2(n539), .ZN(n548) );
  NAND2_X1 U609 ( .A1(G113), .A2(n884), .ZN(n544) );
  NAND2_X1 U610 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n546), .B(KEYINPUT67), .ZN(n547) );
  NAND2_X1 U612 ( .A1(G138), .A2(n879), .ZN(n553) );
  BUF_X1 U613 ( .A(n551), .Z(n880) );
  NAND2_X1 U614 ( .A1(G102), .A2(n880), .ZN(n552) );
  NAND2_X1 U615 ( .A1(n553), .A2(n552), .ZN(n557) );
  NAND2_X1 U616 ( .A1(G114), .A2(n884), .ZN(n555) );
  NAND2_X1 U617 ( .A1(G126), .A2(n524), .ZN(n554) );
  NAND2_X1 U618 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U619 ( .A1(n557), .A2(n556), .ZN(G164) );
  NAND2_X1 U620 ( .A1(G63), .A2(n801), .ZN(n559) );
  NAND2_X1 U621 ( .A1(G51), .A2(n802), .ZN(n558) );
  NAND2_X1 U622 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U623 ( .A(KEYINPUT6), .B(n560), .Z(n568) );
  NAND2_X1 U624 ( .A1(G76), .A2(n797), .ZN(n564) );
  XOR2_X1 U625 ( .A(KEYINPUT4), .B(KEYINPUT71), .Z(n562) );
  NAND2_X1 U626 ( .A1(G89), .A2(n796), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(n563) );
  NAND2_X1 U628 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U629 ( .A(n565), .B(KEYINPUT5), .ZN(n566) );
  XNOR2_X1 U630 ( .A(KEYINPUT72), .B(n566), .ZN(n567) );
  NAND2_X1 U631 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U632 ( .A(KEYINPUT7), .B(n569), .ZN(G168) );
  NAND2_X1 U633 ( .A1(G91), .A2(n796), .ZN(n571) );
  NAND2_X1 U634 ( .A1(G78), .A2(n797), .ZN(n570) );
  NAND2_X1 U635 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U636 ( .A(KEYINPUT68), .B(n572), .ZN(n575) );
  NAND2_X1 U637 ( .A1(G53), .A2(n802), .ZN(n573) );
  XNOR2_X1 U638 ( .A(KEYINPUT69), .B(n573), .ZN(n574) );
  NOR2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U640 ( .A1(n801), .A2(G65), .ZN(n576) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(G299) );
  XOR2_X1 U642 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U643 ( .A1(G62), .A2(n801), .ZN(n579) );
  NAND2_X1 U644 ( .A1(G50), .A2(n802), .ZN(n578) );
  NAND2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(KEYINPUT81), .B(n580), .ZN(n585) );
  NAND2_X1 U647 ( .A1(G88), .A2(n796), .ZN(n582) );
  NAND2_X1 U648 ( .A1(G75), .A2(n797), .ZN(n581) );
  NAND2_X1 U649 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U650 ( .A(KEYINPUT82), .B(n583), .Z(n584) );
  NAND2_X1 U651 ( .A1(n585), .A2(n584), .ZN(G303) );
  INV_X1 U652 ( .A(G303), .ZN(G166) );
  NAND2_X1 U653 ( .A1(G49), .A2(n802), .ZN(n587) );
  NAND2_X1 U654 ( .A1(G74), .A2(G651), .ZN(n586) );
  NAND2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U656 ( .A(KEYINPUT78), .B(n588), .ZN(n589) );
  NOR2_X1 U657 ( .A1(n801), .A2(n589), .ZN(n590) );
  XOR2_X1 U658 ( .A(KEYINPUT79), .B(n590), .Z(n593) );
  NAND2_X1 U659 ( .A1(n591), .A2(G87), .ZN(n592) );
  NAND2_X1 U660 ( .A1(n593), .A2(n592), .ZN(G288) );
  XOR2_X1 U661 ( .A(KEYINPUT2), .B(KEYINPUT80), .Z(n595) );
  NAND2_X1 U662 ( .A1(G73), .A2(n797), .ZN(n594) );
  XNOR2_X1 U663 ( .A(n595), .B(n594), .ZN(n599) );
  NAND2_X1 U664 ( .A1(G61), .A2(n801), .ZN(n597) );
  NAND2_X1 U665 ( .A1(G86), .A2(n796), .ZN(n596) );
  NAND2_X1 U666 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U667 ( .A1(n599), .A2(n598), .ZN(n601) );
  NAND2_X1 U668 ( .A1(n802), .A2(G48), .ZN(n600) );
  NAND2_X1 U669 ( .A1(n601), .A2(n600), .ZN(G305) );
  NAND2_X1 U670 ( .A1(G85), .A2(n796), .ZN(n603) );
  NAND2_X1 U671 ( .A1(G72), .A2(n797), .ZN(n602) );
  NAND2_X1 U672 ( .A1(n603), .A2(n602), .ZN(n607) );
  NAND2_X1 U673 ( .A1(G60), .A2(n801), .ZN(n605) );
  NAND2_X1 U674 ( .A1(G47), .A2(n802), .ZN(n604) );
  NAND2_X1 U675 ( .A1(n605), .A2(n604), .ZN(n606) );
  OR2_X1 U676 ( .A1(n607), .A2(n606), .ZN(G290) );
  NAND2_X1 U677 ( .A1(n608), .A2(G40), .ZN(n716) );
  INV_X1 U678 ( .A(n716), .ZN(n609) );
  NOR2_X1 U679 ( .A1(G164), .A2(G1384), .ZN(n717) );
  NAND2_X1 U680 ( .A1(n609), .A2(n717), .ZN(n614) );
  INV_X2 U681 ( .A(n614), .ZN(n646) );
  XNOR2_X1 U682 ( .A(n610), .B(KEYINPUT95), .ZN(n612) );
  XNOR2_X1 U683 ( .A(G2078), .B(KEYINPUT25), .ZN(n1026) );
  NAND2_X1 U684 ( .A1(n646), .A2(n1026), .ZN(n611) );
  NAND2_X1 U685 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U686 ( .A(KEYINPUT96), .B(n613), .ZN(n660) );
  NOR2_X2 U687 ( .A1(G1966), .A2(n667), .ZN(n682) );
  INV_X1 U688 ( .A(n646), .ZN(n668) );
  NOR2_X1 U689 ( .A1(G2084), .A2(n668), .ZN(n677) );
  NOR2_X1 U690 ( .A1(n682), .A2(n677), .ZN(n616) );
  NAND2_X1 U691 ( .A1(G8), .A2(n616), .ZN(n617) );
  XNOR2_X1 U692 ( .A(n617), .B(KEYINPUT30), .ZN(n618) );
  NOR2_X1 U693 ( .A1(n618), .A2(G168), .ZN(n619) );
  XNOR2_X1 U694 ( .A(n621), .B(KEYINPUT31), .ZN(n664) );
  INV_X1 U695 ( .A(G299), .ZN(n964) );
  NAND2_X1 U696 ( .A1(n646), .A2(G2072), .ZN(n622) );
  INV_X1 U697 ( .A(G1956), .ZN(n942) );
  NOR2_X1 U698 ( .A1(n942), .A2(n646), .ZN(n623) );
  NOR2_X1 U699 ( .A1(n964), .A2(n654), .ZN(n625) );
  AND2_X1 U700 ( .A1(n646), .A2(G1996), .ZN(n626) );
  XOR2_X1 U701 ( .A(n626), .B(KEYINPUT26), .Z(n638) );
  NAND2_X1 U702 ( .A1(n668), .A2(G1341), .ZN(n636) );
  NAND2_X1 U703 ( .A1(G56), .A2(n801), .ZN(n627) );
  XOR2_X1 U704 ( .A(KEYINPUT14), .B(n627), .Z(n633) );
  NAND2_X1 U705 ( .A1(n796), .A2(G81), .ZN(n628) );
  XNOR2_X1 U706 ( .A(n628), .B(KEYINPUT12), .ZN(n630) );
  NAND2_X1 U707 ( .A1(G68), .A2(n797), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U709 ( .A(KEYINPUT13), .B(n631), .Z(n632) );
  NOR2_X1 U710 ( .A1(n633), .A2(n632), .ZN(n635) );
  NAND2_X1 U711 ( .A1(n802), .A2(G43), .ZN(n634) );
  NAND2_X1 U712 ( .A1(n635), .A2(n634), .ZN(n977) );
  INV_X1 U713 ( .A(n977), .ZN(n770) );
  NAND2_X1 U714 ( .A1(G79), .A2(n797), .ZN(n640) );
  NAND2_X1 U715 ( .A1(G54), .A2(n802), .ZN(n639) );
  NAND2_X1 U716 ( .A1(n640), .A2(n639), .ZN(n644) );
  NAND2_X1 U717 ( .A1(G66), .A2(n801), .ZN(n642) );
  NAND2_X1 U718 ( .A1(G92), .A2(n796), .ZN(n641) );
  NAND2_X1 U719 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U720 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U721 ( .A(n645), .B(KEYINPUT15), .ZN(n961) );
  NAND2_X1 U722 ( .A1(G1348), .A2(n668), .ZN(n648) );
  NAND2_X1 U723 ( .A1(G2067), .A2(n646), .ZN(n647) );
  NAND2_X1 U724 ( .A1(n648), .A2(n647), .ZN(n651) );
  NOR2_X1 U725 ( .A1(n961), .A2(n651), .ZN(n649) );
  NAND2_X1 U726 ( .A1(n961), .A2(n651), .ZN(n652) );
  NAND2_X1 U727 ( .A1(n653), .A2(n652), .ZN(n656) );
  NAND2_X1 U728 ( .A1(n964), .A2(n654), .ZN(n655) );
  NAND2_X1 U729 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U730 ( .A(n659), .B(KEYINPUT29), .ZN(n662) );
  AND2_X1 U731 ( .A1(G171), .A2(n660), .ZN(n661) );
  NOR2_X1 U732 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U733 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U734 ( .A(n665), .B(KEYINPUT97), .ZN(n679) );
  NAND2_X1 U735 ( .A1(n679), .A2(G286), .ZN(n666) );
  XNOR2_X1 U736 ( .A(n666), .B(KEYINPUT98), .ZN(n673) );
  NOR2_X1 U737 ( .A1(G1971), .A2(n667), .ZN(n670) );
  NOR2_X1 U738 ( .A1(G2090), .A2(n668), .ZN(n669) );
  NOR2_X1 U739 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U740 ( .A1(n671), .A2(G303), .ZN(n672) );
  NAND2_X1 U741 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U742 ( .A1(n674), .A2(G8), .ZN(n676) );
  INV_X1 U743 ( .A(KEYINPUT32), .ZN(n675) );
  XNOR2_X1 U744 ( .A(n676), .B(n675), .ZN(n684) );
  NAND2_X1 U745 ( .A1(G8), .A2(n677), .ZN(n678) );
  XNOR2_X1 U746 ( .A(n678), .B(KEYINPUT94), .ZN(n680) );
  NAND2_X1 U747 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U748 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X2 U749 ( .A1(n684), .A2(n683), .ZN(n706) );
  INV_X1 U750 ( .A(G1971), .ZN(n967) );
  NAND2_X1 U751 ( .A1(G166), .A2(n967), .ZN(n686) );
  NOR2_X1 U752 ( .A1(G1976), .A2(G288), .ZN(n689) );
  INV_X1 U753 ( .A(n689), .ZN(n685) );
  NAND2_X1 U754 ( .A1(n686), .A2(n685), .ZN(n969) );
  INV_X1 U755 ( .A(n687), .ZN(n696) );
  NAND2_X1 U756 ( .A1(G1976), .A2(G288), .ZN(n971) );
  INV_X1 U757 ( .A(KEYINPUT33), .ZN(n698) );
  NAND2_X1 U758 ( .A1(n711), .A2(n689), .ZN(n690) );
  NOR2_X1 U759 ( .A1(n698), .A2(n690), .ZN(n691) );
  XNOR2_X1 U760 ( .A(n691), .B(KEYINPUT99), .ZN(n697) );
  AND2_X1 U761 ( .A1(n971), .A2(n697), .ZN(n693) );
  XNOR2_X1 U762 ( .A(G1981), .B(G305), .ZN(n959) );
  INV_X1 U763 ( .A(n959), .ZN(n692) );
  AND2_X1 U764 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U765 ( .A1(n696), .A2(n695), .ZN(n702) );
  INV_X1 U766 ( .A(n697), .ZN(n699) );
  OR2_X1 U767 ( .A1(n699), .A2(n698), .ZN(n700) );
  OR2_X1 U768 ( .A1(n959), .A2(n700), .ZN(n701) );
  NAND2_X1 U769 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U770 ( .A(n703), .B(KEYINPUT100), .ZN(n715) );
  NAND2_X1 U771 ( .A1(G166), .A2(G8), .ZN(n704) );
  NOR2_X1 U772 ( .A1(G2090), .A2(n704), .ZN(n705) );
  NOR2_X1 U773 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U774 ( .A(KEYINPUT101), .B(n707), .ZN(n708) );
  NAND2_X1 U775 ( .A1(n708), .A2(n667), .ZN(n713) );
  NOR2_X1 U776 ( .A1(G1981), .A2(G305), .ZN(n709) );
  XNOR2_X1 U777 ( .A(n709), .B(KEYINPUT24), .ZN(n710) );
  NAND2_X1 U778 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U779 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U780 ( .A1(n715), .A2(n714), .ZN(n748) );
  NOR2_X1 U781 ( .A1(n717), .A2(n716), .ZN(n763) );
  NAND2_X1 U782 ( .A1(G140), .A2(n879), .ZN(n719) );
  NAND2_X1 U783 ( .A1(G104), .A2(n880), .ZN(n718) );
  NAND2_X1 U784 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U785 ( .A(KEYINPUT34), .B(n720), .ZN(n727) );
  NAND2_X1 U786 ( .A1(G116), .A2(n884), .ZN(n723) );
  NAND2_X1 U787 ( .A1(G128), .A2(n524), .ZN(n722) );
  NAND2_X1 U788 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U789 ( .A(KEYINPUT89), .B(n724), .ZN(n725) );
  XNOR2_X1 U790 ( .A(KEYINPUT35), .B(n725), .ZN(n726) );
  NOR2_X1 U791 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U792 ( .A(n728), .B(KEYINPUT36), .ZN(n729) );
  XNOR2_X1 U793 ( .A(n729), .B(KEYINPUT90), .ZN(n891) );
  XNOR2_X1 U794 ( .A(KEYINPUT37), .B(G2067), .ZN(n761) );
  NOR2_X1 U795 ( .A1(n891), .A2(n761), .ZN(n990) );
  NAND2_X1 U796 ( .A1(n763), .A2(n990), .ZN(n759) );
  NAND2_X1 U797 ( .A1(G131), .A2(n879), .ZN(n731) );
  NAND2_X1 U798 ( .A1(G107), .A2(n884), .ZN(n730) );
  NAND2_X1 U799 ( .A1(n731), .A2(n730), .ZN(n734) );
  NAND2_X1 U800 ( .A1(G95), .A2(n880), .ZN(n732) );
  XNOR2_X1 U801 ( .A(KEYINPUT91), .B(n732), .ZN(n733) );
  NOR2_X1 U802 ( .A1(n734), .A2(n733), .ZN(n736) );
  NAND2_X1 U803 ( .A1(n524), .A2(G119), .ZN(n735) );
  NAND2_X1 U804 ( .A1(n736), .A2(n735), .ZN(n897) );
  NAND2_X1 U805 ( .A1(G1991), .A2(n897), .ZN(n746) );
  NAND2_X1 U806 ( .A1(G117), .A2(n884), .ZN(n738) );
  NAND2_X1 U807 ( .A1(G129), .A2(n524), .ZN(n737) );
  NAND2_X1 U808 ( .A1(n738), .A2(n737), .ZN(n741) );
  NAND2_X1 U809 ( .A1(G105), .A2(n880), .ZN(n739) );
  XOR2_X1 U810 ( .A(KEYINPUT38), .B(n739), .Z(n740) );
  NOR2_X1 U811 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U812 ( .A(n742), .B(KEYINPUT92), .ZN(n744) );
  NAND2_X1 U813 ( .A1(G141), .A2(n879), .ZN(n743) );
  NAND2_X1 U814 ( .A1(n744), .A2(n743), .ZN(n901) );
  NAND2_X1 U815 ( .A1(G1996), .A2(n901), .ZN(n745) );
  NAND2_X1 U816 ( .A1(n746), .A2(n745), .ZN(n996) );
  NAND2_X1 U817 ( .A1(n763), .A2(n996), .ZN(n754) );
  NAND2_X1 U818 ( .A1(n759), .A2(n754), .ZN(n747) );
  XNOR2_X1 U819 ( .A(n749), .B(KEYINPUT102), .ZN(n751) );
  XNOR2_X1 U820 ( .A(G1986), .B(G290), .ZN(n963) );
  NAND2_X1 U821 ( .A1(n963), .A2(n763), .ZN(n750) );
  NAND2_X1 U822 ( .A1(n751), .A2(n750), .ZN(n766) );
  NOR2_X1 U823 ( .A1(G1986), .A2(G290), .ZN(n752) );
  NOR2_X1 U824 ( .A1(G1991), .A2(n897), .ZN(n992) );
  NOR2_X1 U825 ( .A1(n752), .A2(n992), .ZN(n753) );
  XNOR2_X1 U826 ( .A(n753), .B(KEYINPUT103), .ZN(n755) );
  NAND2_X1 U827 ( .A1(n755), .A2(n754), .ZN(n756) );
  OR2_X1 U828 ( .A1(n901), .A2(G1996), .ZN(n1003) );
  NAND2_X1 U829 ( .A1(n756), .A2(n1003), .ZN(n758) );
  XOR2_X1 U830 ( .A(KEYINPUT39), .B(KEYINPUT104), .Z(n757) );
  XNOR2_X1 U831 ( .A(n758), .B(n757), .ZN(n760) );
  NAND2_X1 U832 ( .A1(n760), .A2(n759), .ZN(n762) );
  NAND2_X1 U833 ( .A1(n891), .A2(n761), .ZN(n993) );
  NAND2_X1 U834 ( .A1(n762), .A2(n993), .ZN(n764) );
  NAND2_X1 U835 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U836 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U837 ( .A(n767), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U838 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U839 ( .A(G120), .ZN(G236) );
  INV_X1 U840 ( .A(G69), .ZN(G235) );
  INV_X1 U841 ( .A(G108), .ZN(G238) );
  INV_X1 U842 ( .A(G132), .ZN(G219) );
  INV_X1 U843 ( .A(G82), .ZN(G220) );
  NAND2_X1 U844 ( .A1(G7), .A2(G661), .ZN(n768) );
  XNOR2_X1 U845 ( .A(n768), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U846 ( .A(G223), .ZN(n851) );
  AND2_X1 U847 ( .A1(G567), .A2(n851), .ZN(n769) );
  XNOR2_X1 U848 ( .A(n769), .B(KEYINPUT11), .ZN(G234) );
  NAND2_X1 U849 ( .A1(n770), .A2(G860), .ZN(G153) );
  INV_X1 U850 ( .A(G171), .ZN(G301) );
  NOR2_X1 U851 ( .A1(G868), .A2(n961), .ZN(n772) );
  INV_X1 U852 ( .A(G868), .ZN(n817) );
  NOR2_X1 U853 ( .A1(n817), .A2(G301), .ZN(n771) );
  NOR2_X1 U854 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U855 ( .A(KEYINPUT70), .B(n773), .ZN(G284) );
  NOR2_X1 U856 ( .A1(G286), .A2(n817), .ZN(n775) );
  NOR2_X1 U857 ( .A1(G868), .A2(G299), .ZN(n774) );
  NOR2_X1 U858 ( .A1(n775), .A2(n774), .ZN(G297) );
  INV_X1 U859 ( .A(G559), .ZN(n776) );
  NOR2_X1 U860 ( .A1(G860), .A2(n776), .ZN(n777) );
  XNOR2_X1 U861 ( .A(KEYINPUT73), .B(n777), .ZN(n778) );
  INV_X1 U862 ( .A(n961), .ZN(n793) );
  NAND2_X1 U863 ( .A1(n778), .A2(n793), .ZN(n779) );
  XNOR2_X1 U864 ( .A(n779), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U865 ( .A1(G868), .A2(n977), .ZN(n782) );
  NAND2_X1 U866 ( .A1(G868), .A2(n793), .ZN(n780) );
  NOR2_X1 U867 ( .A1(G559), .A2(n780), .ZN(n781) );
  NOR2_X1 U868 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U869 ( .A(KEYINPUT74), .B(n783), .ZN(G282) );
  NAND2_X1 U870 ( .A1(G135), .A2(n879), .ZN(n785) );
  NAND2_X1 U871 ( .A1(G111), .A2(n884), .ZN(n784) );
  NAND2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n790) );
  NAND2_X1 U873 ( .A1(G123), .A2(n524), .ZN(n786) );
  XNOR2_X1 U874 ( .A(n786), .B(KEYINPUT18), .ZN(n788) );
  NAND2_X1 U875 ( .A1(G99), .A2(n880), .ZN(n787) );
  NAND2_X1 U876 ( .A1(n788), .A2(n787), .ZN(n789) );
  NOR2_X1 U877 ( .A1(n790), .A2(n789), .ZN(n991) );
  XNOR2_X1 U878 ( .A(n991), .B(G2096), .ZN(n792) );
  INV_X1 U879 ( .A(G2100), .ZN(n791) );
  NAND2_X1 U880 ( .A1(n792), .A2(n791), .ZN(G156) );
  NAND2_X1 U881 ( .A1(G559), .A2(n793), .ZN(n794) );
  XOR2_X1 U882 ( .A(KEYINPUT75), .B(n794), .Z(n795) );
  XNOR2_X1 U883 ( .A(n977), .B(n795), .ZN(n815) );
  NOR2_X1 U884 ( .A1(n815), .A2(G860), .ZN(n808) );
  NAND2_X1 U885 ( .A1(G93), .A2(n796), .ZN(n799) );
  NAND2_X1 U886 ( .A1(G80), .A2(n797), .ZN(n798) );
  NAND2_X1 U887 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U888 ( .A(KEYINPUT76), .B(n800), .ZN(n807) );
  NAND2_X1 U889 ( .A1(G67), .A2(n801), .ZN(n804) );
  NAND2_X1 U890 ( .A1(G55), .A2(n802), .ZN(n803) );
  NAND2_X1 U891 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U892 ( .A(KEYINPUT77), .B(n805), .Z(n806) );
  OR2_X1 U893 ( .A1(n807), .A2(n806), .ZN(n818) );
  XOR2_X1 U894 ( .A(n808), .B(n818), .Z(G145) );
  XOR2_X1 U895 ( .A(KEYINPUT83), .B(KEYINPUT19), .Z(n809) );
  XNOR2_X1 U896 ( .A(G305), .B(n809), .ZN(n810) );
  XNOR2_X1 U897 ( .A(G166), .B(n810), .ZN(n812) );
  XNOR2_X1 U898 ( .A(G290), .B(n964), .ZN(n811) );
  XNOR2_X1 U899 ( .A(n812), .B(n811), .ZN(n813) );
  XOR2_X1 U900 ( .A(n818), .B(n813), .Z(n814) );
  XNOR2_X1 U901 ( .A(n814), .B(G288), .ZN(n858) );
  XNOR2_X1 U902 ( .A(n815), .B(n858), .ZN(n816) );
  NAND2_X1 U903 ( .A1(n816), .A2(G868), .ZN(n820) );
  NAND2_X1 U904 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U905 ( .A1(n820), .A2(n819), .ZN(G295) );
  NAND2_X1 U906 ( .A1(G2078), .A2(G2084), .ZN(n822) );
  XOR2_X1 U907 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n821) );
  XNOR2_X1 U908 ( .A(n822), .B(n821), .ZN(n823) );
  NAND2_X1 U909 ( .A1(G2090), .A2(n823), .ZN(n824) );
  XNOR2_X1 U910 ( .A(KEYINPUT21), .B(n824), .ZN(n825) );
  NAND2_X1 U911 ( .A1(n825), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U912 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U913 ( .A1(G220), .A2(G219), .ZN(n826) );
  XOR2_X1 U914 ( .A(KEYINPUT22), .B(n826), .Z(n827) );
  NOR2_X1 U915 ( .A1(G218), .A2(n827), .ZN(n828) );
  NAND2_X1 U916 ( .A1(G96), .A2(n828), .ZN(n856) );
  NAND2_X1 U917 ( .A1(G2106), .A2(n856), .ZN(n829) );
  XNOR2_X1 U918 ( .A(n829), .B(KEYINPUT85), .ZN(n835) );
  NOR2_X1 U919 ( .A1(G235), .A2(G236), .ZN(n830) );
  XOR2_X1 U920 ( .A(KEYINPUT86), .B(n830), .Z(n831) );
  NOR2_X1 U921 ( .A1(G238), .A2(n831), .ZN(n832) );
  NAND2_X1 U922 ( .A1(n832), .A2(G57), .ZN(n833) );
  XOR2_X1 U923 ( .A(n833), .B(KEYINPUT87), .Z(n857) );
  AND2_X1 U924 ( .A1(G567), .A2(n857), .ZN(n834) );
  NOR2_X1 U925 ( .A1(n835), .A2(n834), .ZN(G319) );
  NAND2_X1 U926 ( .A1(G661), .A2(G483), .ZN(n837) );
  INV_X1 U927 ( .A(G319), .ZN(n836) );
  NOR2_X1 U928 ( .A1(n837), .A2(n836), .ZN(n838) );
  XNOR2_X1 U929 ( .A(n838), .B(KEYINPUT88), .ZN(n854) );
  NAND2_X1 U930 ( .A1(G36), .A2(n854), .ZN(G176) );
  XOR2_X1 U931 ( .A(KEYINPUT107), .B(G2446), .Z(n840) );
  XNOR2_X1 U932 ( .A(G2454), .B(G2451), .ZN(n839) );
  XNOR2_X1 U933 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U934 ( .A(n841), .B(G2430), .Z(n843) );
  XNOR2_X1 U935 ( .A(G1341), .B(G1348), .ZN(n842) );
  XNOR2_X1 U936 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U937 ( .A(KEYINPUT105), .B(G2435), .Z(n845) );
  XNOR2_X1 U938 ( .A(KEYINPUT106), .B(G2438), .ZN(n844) );
  XNOR2_X1 U939 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U940 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U941 ( .A(G2443), .B(G2427), .ZN(n848) );
  XNOR2_X1 U942 ( .A(n849), .B(n848), .ZN(n850) );
  NAND2_X1 U943 ( .A1(n850), .A2(G14), .ZN(n926) );
  XOR2_X1 U944 ( .A(KEYINPUT108), .B(n926), .Z(G401) );
  NAND2_X1 U945 ( .A1(G2106), .A2(n851), .ZN(G217) );
  AND2_X1 U946 ( .A1(G15), .A2(G2), .ZN(n852) );
  NAND2_X1 U947 ( .A1(G661), .A2(n852), .ZN(G259) );
  NAND2_X1 U948 ( .A1(G3), .A2(G1), .ZN(n853) );
  XOR2_X1 U949 ( .A(KEYINPUT109), .B(n853), .Z(n855) );
  NAND2_X1 U950 ( .A1(n855), .A2(n854), .ZN(G188) );
  INV_X1 U952 ( .A(G96), .ZN(G221) );
  NOR2_X1 U953 ( .A1(n857), .A2(n856), .ZN(G325) );
  INV_X1 U954 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U955 ( .A(G286), .B(n977), .ZN(n859) );
  XNOR2_X1 U956 ( .A(n859), .B(n858), .ZN(n861) );
  XNOR2_X1 U957 ( .A(n961), .B(G171), .ZN(n860) );
  XNOR2_X1 U958 ( .A(n861), .B(n860), .ZN(n862) );
  NOR2_X1 U959 ( .A1(G37), .A2(n862), .ZN(n863) );
  XOR2_X1 U960 ( .A(KEYINPUT115), .B(n863), .Z(G397) );
  NAND2_X1 U961 ( .A1(G124), .A2(n524), .ZN(n864) );
  XNOR2_X1 U962 ( .A(n864), .B(KEYINPUT112), .ZN(n865) );
  XNOR2_X1 U963 ( .A(n865), .B(KEYINPUT44), .ZN(n867) );
  NAND2_X1 U964 ( .A1(G112), .A2(n884), .ZN(n866) );
  NAND2_X1 U965 ( .A1(n867), .A2(n866), .ZN(n871) );
  NAND2_X1 U966 ( .A1(G136), .A2(n879), .ZN(n869) );
  NAND2_X1 U967 ( .A1(G100), .A2(n880), .ZN(n868) );
  NAND2_X1 U968 ( .A1(n869), .A2(n868), .ZN(n870) );
  NOR2_X1 U969 ( .A1(n871), .A2(n870), .ZN(G162) );
  NAND2_X1 U970 ( .A1(G139), .A2(n879), .ZN(n873) );
  NAND2_X1 U971 ( .A1(G103), .A2(n880), .ZN(n872) );
  NAND2_X1 U972 ( .A1(n873), .A2(n872), .ZN(n878) );
  NAND2_X1 U973 ( .A1(G115), .A2(n884), .ZN(n875) );
  NAND2_X1 U974 ( .A1(G127), .A2(n524), .ZN(n874) );
  NAND2_X1 U975 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U976 ( .A(KEYINPUT47), .B(n876), .Z(n877) );
  NOR2_X1 U977 ( .A1(n878), .A2(n877), .ZN(n999) );
  NAND2_X1 U978 ( .A1(G142), .A2(n879), .ZN(n882) );
  NAND2_X1 U979 ( .A1(G106), .A2(n880), .ZN(n881) );
  NAND2_X1 U980 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U981 ( .A(n883), .B(KEYINPUT45), .ZN(n886) );
  NAND2_X1 U982 ( .A1(G118), .A2(n884), .ZN(n885) );
  NAND2_X1 U983 ( .A1(n886), .A2(n885), .ZN(n889) );
  NAND2_X1 U984 ( .A1(G130), .A2(n524), .ZN(n887) );
  XNOR2_X1 U985 ( .A(KEYINPUT113), .B(n887), .ZN(n888) );
  NOR2_X1 U986 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U987 ( .A(n999), .B(n890), .ZN(n893) );
  XNOR2_X1 U988 ( .A(G160), .B(n891), .ZN(n892) );
  XNOR2_X1 U989 ( .A(n893), .B(n892), .ZN(n903) );
  XOR2_X1 U990 ( .A(KEYINPUT48), .B(KEYINPUT114), .Z(n895) );
  XNOR2_X1 U991 ( .A(G164), .B(KEYINPUT46), .ZN(n894) );
  XNOR2_X1 U992 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n991), .B(n896), .ZN(n899) );
  XNOR2_X1 U994 ( .A(n897), .B(G162), .ZN(n898) );
  XNOR2_X1 U995 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U996 ( .A(n901), .B(n900), .Z(n902) );
  XNOR2_X1 U997 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U998 ( .A1(G37), .A2(n904), .ZN(G395) );
  XOR2_X1 U999 ( .A(KEYINPUT110), .B(G1986), .Z(n906) );
  XNOR2_X1 U1000 ( .A(G1996), .B(G1991), .ZN(n905) );
  XNOR2_X1 U1001 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1002 ( .A(n907), .B(KEYINPUT41), .Z(n909) );
  XNOR2_X1 U1003 ( .A(G1966), .B(G1981), .ZN(n908) );
  XNOR2_X1 U1004 ( .A(n909), .B(n908), .ZN(n913) );
  XOR2_X1 U1005 ( .A(G1976), .B(G1971), .Z(n911) );
  XNOR2_X1 U1006 ( .A(G1961), .B(G1956), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(n911), .B(n910), .ZN(n912) );
  XOR2_X1 U1008 ( .A(n913), .B(n912), .Z(n915) );
  XNOR2_X1 U1009 ( .A(KEYINPUT111), .B(G2474), .ZN(n914) );
  XNOR2_X1 U1010 ( .A(n915), .B(n914), .ZN(G229) );
  XOR2_X1 U1011 ( .A(G2100), .B(G2096), .Z(n917) );
  XNOR2_X1 U1012 ( .A(KEYINPUT42), .B(G2678), .ZN(n916) );
  XNOR2_X1 U1013 ( .A(n917), .B(n916), .ZN(n921) );
  XOR2_X1 U1014 ( .A(KEYINPUT43), .B(G2090), .Z(n919) );
  XNOR2_X1 U1015 ( .A(G2067), .B(G2072), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(n919), .B(n918), .ZN(n920) );
  XOR2_X1 U1017 ( .A(n921), .B(n920), .Z(n923) );
  XNOR2_X1 U1018 ( .A(G2078), .B(G2084), .ZN(n922) );
  XNOR2_X1 U1019 ( .A(n923), .B(n922), .ZN(G227) );
  NOR2_X1 U1020 ( .A1(G397), .A2(G395), .ZN(n924) );
  XNOR2_X1 U1021 ( .A(n924), .B(KEYINPUT116), .ZN(n925) );
  NAND2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n929) );
  NOR2_X1 U1023 ( .A1(G229), .A2(G227), .ZN(n927) );
  XNOR2_X1 U1024 ( .A(KEYINPUT49), .B(n927), .ZN(n928) );
  NOR2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1026 ( .A1(G319), .A2(n930), .ZN(G225) );
  INV_X1 U1027 ( .A(G225), .ZN(G308) );
  INV_X1 U1028 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1029 ( .A(G1971), .B(G22), .ZN(n932) );
  XNOR2_X1 U1030 ( .A(G1976), .B(G23), .ZN(n931) );
  NOR2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1032 ( .A(KEYINPUT126), .B(n933), .ZN(n936) );
  XNOR2_X1 U1033 ( .A(G1986), .B(KEYINPUT127), .ZN(n934) );
  XNOR2_X1 U1034 ( .A(n934), .B(G24), .ZN(n935) );
  NAND2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1036 ( .A(n937), .B(KEYINPUT58), .ZN(n955) );
  XNOR2_X1 U1037 ( .A(KEYINPUT124), .B(KEYINPUT125), .ZN(n938) );
  XNOR2_X1 U1038 ( .A(n938), .B(KEYINPUT60), .ZN(n949) );
  XNOR2_X1 U1039 ( .A(G1341), .B(G19), .ZN(n940) );
  XNOR2_X1 U1040 ( .A(G1981), .B(G6), .ZN(n939) );
  NOR2_X1 U1041 ( .A1(n940), .A2(n939), .ZN(n947) );
  XOR2_X1 U1042 ( .A(G1348), .B(KEYINPUT59), .Z(n941) );
  XNOR2_X1 U1043 ( .A(G4), .B(n941), .ZN(n945) );
  XNOR2_X1 U1044 ( .A(KEYINPUT123), .B(G20), .ZN(n943) );
  XNOR2_X1 U1045 ( .A(n943), .B(n942), .ZN(n944) );
  NOR2_X1 U1046 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1047 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1048 ( .A(n949), .B(n948), .ZN(n953) );
  XNOR2_X1 U1049 ( .A(G1966), .B(G21), .ZN(n951) );
  XNOR2_X1 U1050 ( .A(G1961), .B(G5), .ZN(n950) );
  NOR2_X1 U1051 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1052 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1053 ( .A1(n955), .A2(n954), .ZN(n956) );
  XOR2_X1 U1054 ( .A(KEYINPUT61), .B(n956), .Z(n957) );
  NOR2_X1 U1055 ( .A1(G16), .A2(n957), .ZN(n988) );
  XOR2_X1 U1056 ( .A(G1966), .B(G168), .Z(n958) );
  NOR2_X1 U1057 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1058 ( .A(KEYINPUT57), .B(n960), .ZN(n983) );
  XNOR2_X1 U1059 ( .A(G1348), .B(n961), .ZN(n962) );
  NOR2_X1 U1060 ( .A1(n963), .A2(n962), .ZN(n976) );
  XNOR2_X1 U1061 ( .A(n964), .B(G1956), .ZN(n966) );
  XNOR2_X1 U1062 ( .A(G171), .B(G1961), .ZN(n965) );
  NAND2_X1 U1063 ( .A1(n966), .A2(n965), .ZN(n974) );
  NOR2_X1 U1064 ( .A1(G166), .A2(n967), .ZN(n968) );
  NOR2_X1 U1065 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n972) );
  XOR2_X1 U1067 ( .A(KEYINPUT119), .B(n972), .Z(n973) );
  NOR2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n980) );
  XNOR2_X1 U1070 ( .A(n977), .B(G1341), .ZN(n978) );
  XNOR2_X1 U1071 ( .A(KEYINPUT120), .B(n978), .ZN(n979) );
  NOR2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1073 ( .A(KEYINPUT121), .B(n981), .ZN(n982) );
  NOR2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n985) );
  XOR2_X1 U1075 ( .A(KEYINPUT56), .B(G16), .Z(n984) );
  NOR2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1077 ( .A(KEYINPUT122), .B(n986), .ZN(n987) );
  NOR2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n1015) );
  XOR2_X1 U1079 ( .A(G160), .B(G2084), .Z(n989) );
  NOR2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n998) );
  NOR2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n994) );
  NAND2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1084 ( .A1(n998), .A2(n997), .ZN(n1009) );
  XOR2_X1 U1085 ( .A(G2072), .B(n999), .Z(n1001) );
  XOR2_X1 U1086 ( .A(G164), .B(G2078), .Z(n1000) );
  NOR2_X1 U1087 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1088 ( .A(KEYINPUT50), .B(n1002), .ZN(n1007) );
  XNOR2_X1 U1089 ( .A(G2090), .B(G162), .ZN(n1004) );
  NAND2_X1 U1090 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1091 ( .A(n1005), .B(KEYINPUT51), .ZN(n1006) );
  NAND2_X1 U1092 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1093 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1094 ( .A(KEYINPUT52), .B(n1010), .ZN(n1012) );
  INV_X1 U1095 ( .A(KEYINPUT55), .ZN(n1011) );
  NAND2_X1 U1096 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1097 ( .A1(n1013), .A2(G29), .ZN(n1014) );
  NAND2_X1 U1098 ( .A1(n1015), .A2(n1014), .ZN(n1038) );
  XOR2_X1 U1099 ( .A(G2090), .B(G35), .Z(n1018) );
  XOR2_X1 U1100 ( .A(KEYINPUT54), .B(G34), .Z(n1016) );
  XNOR2_X1 U1101 ( .A(G2084), .B(n1016), .ZN(n1017) );
  NAND2_X1 U1102 ( .A1(n1018), .A2(n1017), .ZN(n1031) );
  XNOR2_X1 U1103 ( .A(G1996), .B(G32), .ZN(n1020) );
  XNOR2_X1 U1104 ( .A(G33), .B(G2072), .ZN(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1025) );
  XOR2_X1 U1106 ( .A(G1991), .B(G25), .Z(n1021) );
  NAND2_X1 U1107 ( .A1(n1021), .A2(G28), .ZN(n1023) );
  XNOR2_X1 U1108 ( .A(G26), .B(G2067), .ZN(n1022) );
  NOR2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1028) );
  XOR2_X1 U1111 ( .A(G27), .B(n1026), .Z(n1027) );
  NOR2_X1 U1112 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1113 ( .A(n1029), .B(KEYINPUT53), .ZN(n1030) );
  NOR2_X1 U1114 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XOR2_X1 U1115 ( .A(KEYINPUT55), .B(n1032), .Z(n1033) );
  NOR2_X1 U1116 ( .A1(G29), .A2(n1033), .ZN(n1034) );
  XNOR2_X1 U1117 ( .A(KEYINPUT117), .B(n1034), .ZN(n1035) );
  NAND2_X1 U1118 ( .A1(n1035), .A2(G11), .ZN(n1036) );
  XNOR2_X1 U1119 ( .A(n1036), .B(KEYINPUT118), .ZN(n1037) );
  NOR2_X1 U1120 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  XNOR2_X1 U1121 ( .A(n1039), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1122 ( .A(G311), .ZN(G150) );
endmodule

