//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1 0 1 1 1 1 0 1 0 1 1 1 1 0 0 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G20), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n202), .A2(G50), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G68), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n210), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n213), .B1(new_n216), .B2(new_n217), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT64), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G87), .B(G97), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT65), .ZN(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  XNOR2_X1  g0046(.A(KEYINPUT8), .B(G58), .ZN(new_n247));
  AOI21_X1  g0047(.A(new_n247), .B1(new_n207), .B2(G20), .ZN(new_n248));
  INV_X1    g0048(.A(G13), .ZN(new_n249));
  NOR3_X1   g0049(.A1(new_n249), .A2(new_n208), .A3(G1), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n214), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  AOI22_X1  g0053(.A1(new_n248), .A2(new_n253), .B1(new_n250), .B2(new_n247), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n252), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT3), .B(G33), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT7), .ZN(new_n258));
  NOR3_X1   g0058(.A1(new_n257), .A2(new_n258), .A3(G20), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT3), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(KEYINPUT7), .B1(new_n264), .B2(new_n208), .ZN(new_n265));
  OAI21_X1  g0065(.A(G68), .B1(new_n259), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n208), .A2(new_n260), .A3(KEYINPUT66), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT66), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n268), .B1(G20), .B2(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G159), .ZN(new_n271));
  INV_X1    g0071(.A(G58), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(new_n219), .ZN(new_n273));
  OAI21_X1  g0073(.A(G20), .B1(new_n273), .B2(new_n201), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n266), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT16), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n256), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AND3_X1   g0079(.A1(new_n260), .A2(KEYINPUT70), .A3(KEYINPUT3), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT70), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n280), .B1(new_n257), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n258), .B1(new_n282), .B2(new_n208), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n261), .A2(new_n263), .A3(new_n281), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n260), .A2(KEYINPUT70), .A3(KEYINPUT3), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n284), .A2(new_n258), .A3(new_n208), .A4(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G68), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n276), .B(KEYINPUT16), .C1(new_n283), .C2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n255), .B1(new_n279), .B2(new_n288), .ZN(new_n289));
  XOR2_X1   g0089(.A(KEYINPUT73), .B(KEYINPUT17), .Z(new_n290));
  AOI21_X1  g0090(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n291));
  INV_X1    g0091(.A(G274), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G232), .ZN(new_n297));
  INV_X1    g0097(.A(new_n291), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n294), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n296), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT71), .ZN(new_n301));
  INV_X1    g0101(.A(G1698), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G223), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n301), .B1(new_n282), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(G33), .A2(G87), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n284), .A2(new_n285), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n306), .A2(G226), .A3(G1698), .ZN(new_n307));
  INV_X1    g0107(.A(new_n303), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n306), .A2(KEYINPUT71), .A3(new_n308), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n304), .A2(new_n305), .A3(new_n307), .A4(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n300), .B1(new_n310), .B2(new_n291), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n311), .A2(G200), .ZN(new_n312));
  AOI211_X1 g0112(.A(G190), .B(new_n300), .C1(new_n310), .C2(new_n291), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n289), .B(new_n290), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n258), .B1(new_n257), .B2(G20), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n264), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n219), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n278), .B1(new_n317), .B2(new_n275), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n288), .A2(new_n252), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n254), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n310), .A2(new_n291), .ZN(new_n321));
  INV_X1    g0121(.A(new_n300), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G200), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G190), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n311), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n320), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT17), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n314), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT74), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n289), .B1(new_n312), .B2(new_n313), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT17), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n334), .A2(KEYINPUT74), .A3(new_n314), .ZN(new_n335));
  INV_X1    g0135(.A(G169), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n311), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G179), .ZN(new_n338));
  AOI211_X1 g0138(.A(new_n338), .B(new_n300), .C1(new_n310), .C2(new_n291), .ZN(new_n339));
  OAI211_X1 g0139(.A(KEYINPUT18), .B(new_n320), .C1(new_n337), .C2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n321), .A2(G179), .A3(new_n322), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(new_n336), .B2(new_n311), .ZN(new_n343));
  AOI21_X1  g0143(.A(KEYINPUT18), .B1(new_n343), .B2(new_n320), .ZN(new_n344));
  OAI21_X1  g0144(.A(KEYINPUT72), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n320), .B1(new_n337), .B2(new_n339), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT18), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT72), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n332), .A2(new_n335), .B1(new_n345), .B2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(G222), .A2(G1698), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n302), .A2(G223), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n257), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n354), .B(new_n291), .C1(G77), .C2(new_n257), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n291), .A2(new_n295), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(G226), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n355), .A2(new_n296), .A3(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n358), .A2(G179), .ZN(new_n359));
  OAI21_X1  g0159(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n208), .A2(G33), .ZN(new_n361));
  INV_X1    g0161(.A(new_n270), .ZN(new_n362));
  INV_X1    g0162(.A(G150), .ZN(new_n363));
  OAI221_X1 g0163(.A(new_n360), .B1(new_n247), .B2(new_n361), .C1(new_n362), .C2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n252), .ZN(new_n365));
  INV_X1    g0165(.A(G50), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n366), .B1(new_n207), .B2(G20), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n253), .A2(new_n367), .B1(new_n366), .B2(new_n250), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  AOI211_X1 g0170(.A(new_n359), .B(new_n370), .C1(new_n336), .C2(new_n358), .ZN(new_n371));
  AOI21_X1  g0171(.A(KEYINPUT68), .B1(new_n358), .B2(G200), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(new_n326), .B2(new_n358), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n373), .B1(KEYINPUT9), .B2(new_n370), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT67), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n370), .B2(KEYINPUT9), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT9), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n369), .A2(KEYINPUT67), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n374), .A2(new_n379), .ZN(new_n380));
  OR2_X1    g0180(.A1(new_n380), .A2(KEYINPUT10), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(KEYINPUT10), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n371), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n362), .A2(new_n366), .ZN(new_n384));
  INV_X1    g0184(.A(G77), .ZN(new_n385));
  OAI22_X1  g0185(.A1(new_n361), .A2(new_n385), .B1(new_n208), .B2(G68), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n252), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT11), .ZN(new_n388));
  AND2_X1   g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n250), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT12), .B1(new_n390), .B2(G68), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT12), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n250), .A2(new_n392), .A3(new_n219), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n219), .B1(new_n207), .B2(G20), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n391), .A2(new_n393), .B1(new_n253), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n387), .B2(new_n388), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n389), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n297), .A2(G1698), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n257), .B(new_n398), .C1(G226), .C2(G1698), .ZN(new_n399));
  NAND2_X1  g0199(.A1(G33), .A2(G97), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n298), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NOR3_X1   g0202(.A1(new_n291), .A2(new_n292), .A3(new_n294), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n403), .B1(G238), .B2(new_n356), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT13), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n402), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n296), .B1(new_n220), .B2(new_n299), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT13), .B1(new_n407), .B2(new_n401), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n397), .B1(new_n409), .B2(new_n326), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT69), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n406), .A2(new_n408), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n411), .B1(new_n412), .B2(new_n324), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n409), .A2(KEYINPUT69), .A3(G200), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n410), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT14), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n416), .B1(new_n409), .B2(G169), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n409), .A2(new_n416), .A3(G169), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n418), .B(new_n419), .C1(new_n338), .C2(new_n409), .ZN(new_n420));
  OR2_X1    g0220(.A1(new_n389), .A2(new_n396), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n415), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  XOR2_X1   g0222(.A(KEYINPUT15), .B(G87), .Z(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  OAI22_X1  g0224(.A1(new_n424), .A2(new_n361), .B1(new_n208), .B2(new_n385), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n362), .A2(new_n247), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n252), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n385), .B1(new_n207), .B2(G20), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n253), .A2(new_n428), .B1(new_n385), .B2(new_n250), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n257), .A2(G232), .A3(new_n302), .ZN(new_n432));
  INV_X1    g0232(.A(G107), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n257), .A2(G1698), .ZN(new_n434));
  OAI221_X1 g0234(.A(new_n432), .B1(new_n433), .B2(new_n257), .C1(new_n434), .C2(new_n220), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n291), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n403), .B1(G244), .B2(new_n356), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n431), .B1(new_n336), .B2(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n438), .A2(G179), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n438), .A2(G200), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n443), .B(new_n431), .C1(new_n326), .C2(new_n438), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n351), .A2(new_n383), .A3(new_n422), .A4(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(G1698), .B1(new_n284), .B2(new_n285), .ZN(new_n448));
  AOI21_X1  g0248(.A(KEYINPUT4), .B1(new_n448), .B2(G244), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n257), .A2(KEYINPUT4), .A3(G244), .A4(new_n302), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G33), .A2(G283), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n450), .B(new_n451), .C1(new_n434), .C2(new_n222), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n291), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  XNOR2_X1  g0253(.A(KEYINPUT5), .B(G41), .ZN(new_n454));
  INV_X1    g0254(.A(G45), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n455), .A2(G1), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n298), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(G257), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n293), .A2(new_n456), .A3(new_n454), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n453), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  OR2_X1    g0262(.A1(new_n462), .A2(new_n326), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT6), .ZN(new_n464));
  INV_X1    g0264(.A(G97), .ZN(new_n465));
  NOR3_X1   g0265(.A1(new_n464), .A2(new_n465), .A3(G107), .ZN(new_n466));
  XNOR2_X1  g0266(.A(G97), .B(G107), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n466), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  OAI22_X1  g0268(.A1(new_n468), .A2(new_n208), .B1(new_n385), .B2(new_n362), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n433), .B1(new_n315), .B2(new_n316), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n252), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n390), .A2(G97), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n260), .A2(G1), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n250), .A2(new_n252), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n472), .B1(new_n474), .B2(G97), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n476), .B1(new_n462), .B2(G200), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n462), .A2(new_n336), .B1(new_n471), .B2(new_n475), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n453), .A2(new_n338), .A3(new_n460), .A4(new_n461), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n463), .A2(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n390), .A2(new_n423), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n208), .A2(G33), .A3(G97), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT77), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT19), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n483), .B1(new_n482), .B2(new_n484), .ZN(new_n486));
  NAND3_X1  g0286(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n208), .A2(new_n487), .B1(new_n204), .B2(new_n221), .ZN(new_n488));
  NOR3_X1   g0288(.A1(new_n485), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(G20), .B1(new_n284), .B2(new_n285), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT76), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n490), .A2(new_n491), .A3(G68), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n491), .B1(new_n490), .B2(G68), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n489), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n481), .B1(new_n495), .B2(new_n252), .ZN(new_n496));
  INV_X1    g0296(.A(new_n474), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n497), .A2(new_n221), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n293), .A2(new_n456), .ZN(new_n500));
  OAI21_X1  g0300(.A(G250), .B1(new_n455), .B2(G1), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n500), .B1(new_n291), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n306), .A2(G244), .A3(G1698), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n306), .A2(G238), .A3(new_n302), .ZN(new_n504));
  OR2_X1    g0304(.A1(KEYINPUT75), .A2(G116), .ZN(new_n505));
  NAND2_X1  g0305(.A1(KEYINPUT75), .A2(G116), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G33), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n503), .A2(new_n504), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n502), .B1(new_n509), .B2(new_n291), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n510), .A2(G200), .ZN(new_n511));
  AOI211_X1 g0311(.A(G190), .B(new_n502), .C1(new_n509), .C2(new_n291), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n496), .B(new_n499), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n481), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n474), .A2(new_n423), .ZN(new_n515));
  INV_X1    g0315(.A(new_n489), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n306), .A2(new_n208), .A3(G68), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(KEYINPUT76), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n516), .B1(new_n518), .B2(new_n492), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n514), .B(new_n515), .C1(new_n519), .C2(new_n256), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n510), .A2(new_n338), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n448), .A2(G238), .B1(G33), .B2(new_n507), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n298), .B1(new_n522), .B2(new_n503), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n336), .B1(new_n523), .B2(new_n502), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n520), .A2(new_n521), .A3(new_n524), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n513), .A2(new_n525), .A3(KEYINPUT78), .ZN(new_n526));
  AOI21_X1  g0326(.A(KEYINPUT78), .B1(new_n513), .B2(new_n525), .ZN(new_n527));
  OAI211_X1 g0327(.A(KEYINPUT79), .B(new_n480), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n480), .B1(new_n526), .B2(new_n527), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT79), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(G264), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n461), .B1(new_n532), .B2(new_n458), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n448), .A2(G250), .B1(G33), .B2(G294), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n306), .A2(G257), .A3(G1698), .ZN(new_n536));
  AOI211_X1 g0336(.A(KEYINPUT82), .B(new_n298), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT82), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n306), .A2(G250), .A3(new_n302), .ZN(new_n539));
  NAND2_X1  g0339(.A1(G33), .A2(G294), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n536), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n538), .B1(new_n541), .B2(new_n291), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n534), .B1(new_n537), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G169), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n533), .B1(new_n541), .B2(new_n291), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G179), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(KEYINPUT25), .B1(new_n250), .B2(new_n433), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n250), .A2(KEYINPUT25), .A3(new_n433), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n549), .A2(new_n550), .B1(new_n474), .B2(G107), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT22), .ZN(new_n553));
  NOR4_X1   g0353(.A1(new_n282), .A2(new_n553), .A3(G20), .A4(new_n221), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n208), .A2(G87), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n553), .B1(new_n264), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n433), .A2(G20), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT23), .ZN(new_n558));
  XNOR2_X1  g0358(.A(new_n557), .B(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n556), .B(new_n559), .C1(G20), .C2(new_n508), .ZN(new_n560));
  OR3_X1    g0360(.A1(new_n554), .A2(new_n560), .A3(KEYINPUT24), .ZN(new_n561));
  OAI21_X1  g0361(.A(KEYINPUT24), .B1(new_n554), .B2(new_n560), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n552), .B1(new_n563), .B2(new_n252), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n547), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n326), .B(new_n534), .C1(new_n537), .C2(new_n542), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT83), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(new_n545), .B2(G200), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n298), .B1(new_n535), .B2(new_n536), .ZN(new_n570));
  OAI211_X1 g0370(.A(KEYINPUT83), .B(new_n324), .C1(new_n570), .C2(new_n533), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n567), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n564), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n306), .A2(G257), .A3(new_n302), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n306), .A2(G264), .A3(G1698), .ZN(new_n575));
  XOR2_X1   g0375(.A(KEYINPUT80), .B(G303), .Z(new_n576));
  OAI211_X1 g0376(.A(new_n574), .B(new_n575), .C1(new_n257), .C2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n291), .ZN(new_n578));
  INV_X1    g0378(.A(G270), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n461), .B1(new_n579), .B2(new_n458), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(KEYINPUT81), .A2(KEYINPUT21), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n451), .B(new_n208), .C1(G33), .C2(new_n465), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n252), .B(new_n585), .C1(new_n507), .C2(new_n208), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT20), .ZN(new_n587));
  XNOR2_X1  g0387(.A(new_n586), .B(new_n587), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n505), .A2(new_n506), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n474), .A2(G116), .B1(new_n250), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n336), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n582), .A2(new_n584), .A3(new_n591), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n586), .A2(new_n587), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n586), .A2(new_n587), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n590), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(G169), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n580), .B1(new_n577), .B2(new_n291), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n583), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n597), .A2(G179), .A3(new_n595), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n592), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n595), .B1(new_n582), .B2(G200), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n326), .B2(new_n582), .ZN(new_n602));
  AND4_X1   g0402(.A1(new_n566), .A2(new_n573), .A3(new_n600), .A4(new_n602), .ZN(new_n603));
  AND4_X1   g0403(.A1(new_n447), .A2(new_n528), .A3(new_n531), .A4(new_n603), .ZN(G372));
  NAND2_X1  g0404(.A1(new_n413), .A2(new_n414), .ZN(new_n605));
  INV_X1    g0405(.A(new_n410), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n438), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n430), .B1(new_n608), .B2(G169), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n609), .A2(new_n440), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n419), .B1(new_n338), .B2(new_n409), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n421), .B1(new_n612), .B2(new_n417), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT85), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n332), .A2(new_n335), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n611), .A2(KEYINPUT85), .A3(new_n613), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n348), .A2(new_n340), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n381), .A2(new_n382), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n371), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n478), .A2(new_n479), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n624), .B1(new_n526), .B2(new_n527), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(KEYINPUT26), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT84), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n521), .A2(new_n524), .ZN(new_n628));
  AOI211_X1 g0428(.A(new_n481), .B(new_n498), .C1(new_n495), .C2(new_n252), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n510), .A2(new_n326), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n324), .B1(new_n523), .B2(new_n502), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n628), .A2(new_n520), .B1(new_n629), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n573), .A2(new_n633), .A3(new_n480), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n592), .A2(new_n598), .A3(new_n599), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n635), .B1(new_n547), .B2(new_n565), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n627), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT26), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n633), .A2(new_n638), .A3(new_n624), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n639), .A2(new_n525), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n463), .A2(new_n477), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n478), .A2(new_n479), .ZN(new_n642));
  AND4_X1   g0442(.A1(new_n525), .A2(new_n641), .A3(new_n642), .A4(new_n513), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n543), .A2(G169), .B1(G179), .B2(new_n545), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n600), .B1(new_n644), .B2(new_n564), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n643), .A2(new_n645), .A3(KEYINPUT84), .A4(new_n573), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n626), .A2(new_n637), .A3(new_n640), .A4(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n447), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n623), .A2(new_n648), .ZN(G369));
  AND2_X1   g0449(.A1(new_n566), .A2(new_n573), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(new_n653), .A3(G213), .ZN(new_n654));
  INV_X1    g0454(.A(G343), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n650), .B1(new_n564), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n566), .B2(new_n657), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n657), .B1(new_n588), .B2(new_n590), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n635), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n600), .A2(new_n602), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n661), .B1(new_n662), .B2(new_n660), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(G330), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n547), .A2(new_n565), .A3(new_n657), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n600), .A2(new_n656), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n650), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n666), .A2(new_n667), .A3(new_n669), .ZN(G399));
  INV_X1    g0470(.A(G41), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n211), .A2(new_n671), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n205), .A2(G87), .A3(G116), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(G1), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n674), .B1(new_n217), .B2(new_n672), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT28), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT29), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n647), .A2(new_n677), .A3(new_n657), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n643), .A2(new_n573), .A3(new_n645), .ZN(new_n679));
  OAI211_X1 g0479(.A(new_n638), .B(new_n624), .C1(new_n526), .C2(new_n527), .ZN(new_n680));
  INV_X1    g0480(.A(new_n525), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n624), .A2(new_n525), .A3(new_n513), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n681), .B1(new_n682), .B2(KEYINPUT26), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n679), .A2(new_n680), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n657), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(KEYINPUT29), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n678), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(G330), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n510), .A2(new_n453), .A3(new_n460), .ZN(new_n689));
  AOI211_X1 g0489(.A(new_n338), .B(new_n580), .C1(new_n577), .C2(new_n291), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n689), .A2(KEYINPUT30), .A3(new_n545), .A4(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT30), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n545), .A2(new_n510), .A3(new_n453), .A4(new_n460), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n597), .A2(G179), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n597), .A2(new_n545), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n510), .A2(G179), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(new_n462), .A3(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n691), .A2(new_n695), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(KEYINPUT31), .B1(new_n699), .B2(new_n656), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT86), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n699), .A2(KEYINPUT31), .A3(new_n656), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n699), .A2(new_n656), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n704), .A2(KEYINPUT86), .A3(KEYINPUT31), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n531), .A2(new_n603), .A3(new_n528), .A4(new_n657), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n688), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n687), .A2(new_n708), .ZN(new_n709));
  OR2_X1    g0509(.A1(new_n709), .A2(KEYINPUT87), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(KEYINPUT87), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n676), .B1(new_n712), .B2(G1), .ZN(G364));
  INV_X1    g0513(.A(new_n672), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n249), .A2(G20), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n207), .B1(new_n715), .B2(G45), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  OR2_X1    g0518(.A1(G355), .A2(KEYINPUT88), .ZN(new_n719));
  NAND2_X1  g0519(.A1(G355), .A2(KEYINPUT88), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n719), .A2(new_n211), .A3(new_n257), .A4(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(G116), .B2(new_n211), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n282), .A2(new_n211), .ZN(new_n723));
  XOR2_X1   g0523(.A(new_n723), .B(KEYINPUT89), .Z(new_n724));
  NOR2_X1   g0524(.A1(new_n217), .A2(G45), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n725), .B1(new_n245), .B2(G45), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n722), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(G13), .A2(G33), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G20), .ZN(new_n730));
  XOR2_X1   g0530(.A(new_n730), .B(KEYINPUT90), .Z(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n214), .B1(G20), .B2(new_n336), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n718), .B1(new_n727), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n338), .A2(new_n324), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT91), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n738), .A2(new_n208), .A3(G190), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G159), .ZN(new_n740));
  XOR2_X1   g0540(.A(new_n740), .B(KEYINPUT32), .Z(new_n741));
  NOR2_X1   g0541(.A1(new_n208), .A2(new_n338), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n743), .A2(new_n326), .A3(G200), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n743), .A2(G190), .A3(G200), .ZN(new_n745));
  AOI22_X1  g0545(.A1(G58), .A2(new_n744), .B1(new_n745), .B2(G77), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n743), .A2(new_n324), .A3(G190), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n746), .B1(new_n219), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n326), .A2(new_n324), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n208), .A2(G179), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n221), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n750), .A2(new_n742), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n751), .A2(new_n326), .A3(G200), .ZN(new_n755));
  OAI22_X1  g0555(.A1(new_n366), .A2(new_n754), .B1(new_n755), .B2(new_n433), .ZN(new_n756));
  NOR4_X1   g0556(.A1(new_n749), .A2(new_n264), .A3(new_n753), .A4(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(G20), .B1(new_n738), .B2(new_n326), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G97), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n741), .A2(new_n757), .A3(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n754), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n745), .A2(G311), .B1(new_n761), .B2(G326), .ZN(new_n762));
  INV_X1    g0562(.A(new_n758), .ZN(new_n763));
  INV_X1    g0563(.A(G294), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT92), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n739), .A2(G329), .ZN(new_n767));
  XNOR2_X1  g0567(.A(KEYINPUT33), .B(G317), .ZN(new_n768));
  OR2_X1    g0568(.A1(new_n768), .A2(KEYINPUT93), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(KEYINPUT93), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n747), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n752), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n744), .A2(G322), .B1(G303), .B2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n755), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n257), .B1(new_n774), .B2(G283), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n767), .A2(new_n771), .A3(new_n773), .A4(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n760), .B1(new_n766), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n736), .B1(new_n777), .B2(new_n733), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(new_n663), .B2(new_n731), .ZN(new_n779));
  INV_X1    g0579(.A(new_n718), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n664), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n663), .A2(G330), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n779), .B1(new_n781), .B2(new_n782), .ZN(G396));
  NAND2_X1  g0583(.A1(new_n647), .A2(new_n657), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT96), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n609), .A2(new_n440), .A3(new_n656), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n430), .A2(new_n656), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n444), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(new_n442), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n785), .B1(new_n787), .B2(new_n790), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n444), .A2(new_n788), .B1(new_n439), .B2(new_n441), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n792), .A2(KEYINPUT96), .A3(new_n786), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n784), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n647), .A2(new_n657), .A3(new_n794), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n708), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n718), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n796), .A2(new_n708), .A3(new_n797), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n744), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n802), .A2(new_n764), .B1(new_n221), .B2(new_n755), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n257), .B(new_n803), .C1(G107), .C2(new_n772), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n739), .A2(G311), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n761), .A2(G303), .ZN(new_n806));
  INV_X1    g0606(.A(G283), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n806), .B1(new_n748), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(new_n507), .B2(new_n745), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n804), .A2(new_n759), .A3(new_n805), .A4(new_n809), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n747), .A2(G150), .B1(new_n761), .B2(G137), .ZN(new_n811));
  INV_X1    g0611(.A(G143), .ZN(new_n812));
  INV_X1    g0612(.A(G159), .ZN(new_n813));
  INV_X1    g0613(.A(new_n745), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n811), .B1(new_n812), .B2(new_n802), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(KEYINPUT34), .Z(new_n816));
  OAI22_X1  g0616(.A1(new_n755), .A2(new_n219), .B1(new_n752), .B2(new_n366), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n282), .B(new_n817), .C1(new_n739), .C2(G132), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n272), .B2(new_n763), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n810), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  OR2_X1    g0620(.A1(new_n820), .A2(KEYINPUT95), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(KEYINPUT95), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n821), .A2(new_n733), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n733), .A2(new_n728), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT94), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n780), .B1(new_n826), .B2(new_n385), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n823), .B(new_n827), .C1(new_n794), .C2(new_n729), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n801), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(G384));
  NOR2_X1   g0630(.A1(new_n715), .A2(new_n207), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n421), .B(new_n656), .C1(new_n420), .C2(new_n415), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n421), .A2(new_n656), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n613), .A2(new_n607), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n794), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT102), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n702), .B1(new_n700), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n704), .A2(KEYINPUT102), .A3(KEYINPUT31), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI211_X1 g0640(.A(KEYINPUT40), .B(new_n836), .C1(new_n840), .C2(new_n707), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT99), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT38), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n276), .B1(new_n283), .B2(new_n287), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n278), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n845), .A2(new_n288), .A3(new_n252), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n254), .ZN(new_n847));
  INV_X1    g0647(.A(new_n654), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n345), .A2(new_n350), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n849), .B1(new_n617), .B2(new_n850), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n654), .B(KEYINPUT98), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n320), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n333), .A2(new_n346), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n854), .A2(KEYINPUT37), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n343), .A2(new_n847), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n856), .A2(new_n333), .A3(new_n849), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n855), .B1(KEYINPUT37), .B2(new_n857), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n842), .B(new_n843), .C1(new_n851), .C2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n843), .B1(new_n851), .B2(new_n858), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n857), .A2(KEYINPUT37), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(KEYINPUT37), .B2(new_n854), .ZN(new_n862));
  OAI211_X1 g0662(.A(KEYINPUT38), .B(new_n862), .C1(new_n351), .C2(new_n849), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n860), .A2(KEYINPUT99), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n841), .A2(new_n859), .A3(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n836), .ZN(new_n866));
  AND4_X1   g0666(.A1(new_n528), .A2(new_n531), .A3(new_n603), .A4(new_n657), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n838), .A2(new_n839), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n854), .B(KEYINPUT37), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n620), .A2(new_n330), .ZN(new_n871));
  INV_X1    g0671(.A(new_n853), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT38), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n335), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT74), .B1(new_n334), .B2(new_n314), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n349), .B1(new_n348), .B2(new_n340), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n344), .A2(KEYINPUT72), .ZN(new_n878));
  OAI22_X1  g0678(.A1(new_n875), .A2(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n849), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n858), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n874), .B1(new_n881), .B2(KEYINPUT38), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT40), .B1(new_n869), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n865), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n446), .B1(new_n707), .B2(new_n840), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n688), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n885), .B2(new_n884), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n887), .B(KEYINPUT103), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n687), .A2(new_n447), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n623), .ZN(new_n891));
  XOR2_X1   g0691(.A(new_n891), .B(KEYINPUT101), .Z(new_n892));
  NAND3_X1  g0692(.A1(new_n864), .A2(KEYINPUT39), .A3(new_n859), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT100), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT39), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n894), .B1(new_n882), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n420), .A2(new_n421), .A3(new_n657), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n864), .A2(new_n894), .A3(KEYINPUT39), .A4(new_n859), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n897), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n797), .A2(new_n787), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n864), .A2(new_n902), .A3(new_n835), .A4(new_n859), .ZN(new_n903));
  OR2_X1    g0703(.A1(new_n620), .A2(new_n852), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n901), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n892), .B(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n831), .B1(new_n889), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n889), .B2(new_n907), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT35), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n468), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n911), .A2(G20), .A3(G116), .A4(new_n215), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT97), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n912), .A2(new_n913), .B1(new_n910), .B2(new_n468), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n913), .B2(new_n912), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n915), .B(KEYINPUT36), .Z(new_n916));
  NOR3_X1   g0716(.A1(new_n217), .A2(new_n385), .A3(new_n273), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n219), .A2(G50), .ZN(new_n918));
  OAI211_X1 g0718(.A(G1), .B(new_n249), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n909), .A2(new_n916), .A3(new_n919), .ZN(G367));
  NOR2_X1   g0720(.A1(new_n755), .A2(new_n465), .ZN(new_n921));
  AND2_X1   g0721(.A1(KEYINPUT46), .A2(G116), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n921), .B1(new_n772), .B2(new_n922), .ZN(new_n923));
  OAI221_X1 g0723(.A(new_n923), .B1(new_n814), .B2(new_n807), .C1(new_n764), .C2(new_n748), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(G317), .B2(new_n739), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n761), .A2(G311), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n802), .B2(new_n576), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT46), .B1(new_n772), .B2(new_n507), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n927), .A2(new_n306), .A3(new_n928), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n925), .B(new_n929), .C1(new_n433), .C2(new_n763), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n763), .A2(new_n219), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n774), .A2(G77), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n272), .B2(new_n752), .ZN(new_n933));
  AOI211_X1 g0733(.A(new_n264), .B(new_n933), .C1(G150), .C2(new_n744), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n748), .A2(new_n813), .B1(new_n754), .B2(new_n812), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(G50), .B2(new_n745), .ZN(new_n936));
  INV_X1    g0736(.A(G137), .ZN(new_n937));
  INV_X1    g0737(.A(new_n739), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n934), .B(new_n936), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n930), .B1(new_n931), .B2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT47), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n733), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n724), .A2(new_n237), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n943), .B(new_n734), .C1(new_n211), .C2(new_n424), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n942), .A2(new_n718), .A3(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n629), .A2(new_n657), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT104), .Z(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n681), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT105), .ZN(new_n949));
  INV_X1    g0749(.A(new_n633), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n948), .B(new_n949), .C1(new_n950), .C2(new_n947), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n949), .B2(new_n948), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n945), .B1(new_n952), .B2(new_n732), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT108), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n642), .A2(new_n657), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n955), .A2(KEYINPUT106), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(KEYINPUT106), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n476), .A2(new_n656), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n956), .A2(new_n957), .B1(new_n480), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n959), .A2(new_n669), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT107), .Z(new_n961));
  OR2_X1    g0761(.A1(new_n961), .A2(KEYINPUT42), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n959), .A2(new_n566), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n656), .B1(new_n963), .B2(new_n642), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(new_n961), .B2(KEYINPUT42), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT43), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n952), .A2(new_n967), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n952), .A2(new_n967), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n966), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n962), .A2(new_n965), .A3(new_n967), .A4(new_n952), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n666), .A2(new_n959), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n972), .B(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n669), .A2(new_n667), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n959), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT44), .Z(new_n977));
  NOR2_X1   g0777(.A1(new_n975), .A2(new_n959), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT45), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n980), .A2(new_n665), .A3(new_n659), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n977), .A2(new_n666), .A3(new_n979), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n669), .B1(new_n659), .B2(new_n668), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(new_n665), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n983), .A2(new_n985), .B1(new_n710), .B2(new_n711), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n672), .B(KEYINPUT41), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n716), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n954), .B1(new_n974), .B2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(G387));
  AND2_X1   g0790(.A1(new_n712), .A2(new_n985), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n991), .A2(new_n672), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n712), .B2(new_n985), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n659), .A2(new_n731), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n211), .A2(new_n257), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n995), .A2(new_n673), .B1(G107), .B2(new_n211), .ZN(new_n996));
  INV_X1    g0796(.A(new_n724), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n673), .B(new_n455), .C1(new_n219), .C2(new_n385), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT50), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n247), .B2(G50), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n247), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n1001), .A2(KEYINPUT50), .A3(new_n366), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n998), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n997), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n234), .A2(G45), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n996), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n718), .B1(new_n1006), .B2(new_n735), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n748), .A2(new_n247), .B1(new_n814), .B2(new_n219), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n802), .A2(new_n366), .B1(new_n754), .B2(new_n813), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n758), .A2(new_n423), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n739), .A2(G150), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n282), .B(new_n921), .C1(G77), .C2(new_n772), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT109), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n747), .A2(G311), .B1(new_n761), .B2(G322), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n1016), .A2(KEYINPUT110), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(KEYINPUT110), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n576), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n1019), .A2(new_n745), .B1(new_n744), .B2(G317), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1017), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT48), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n763), .A2(new_n807), .B1(new_n764), .B2(new_n752), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1023), .A2(KEYINPUT49), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n739), .A2(G326), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n306), .B1(new_n507), .B2(new_n774), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(KEYINPUT49), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1015), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1007), .B1(new_n1031), .B2(new_n733), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n985), .A2(new_n717), .B1(new_n994), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n993), .A2(new_n1033), .ZN(G393));
  OAI22_X1  g0834(.A1(new_n748), .A2(new_n576), .B1(new_n814), .B2(new_n764), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n257), .B(new_n1035), .C1(G107), .C2(new_n774), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n744), .A2(G311), .B1(new_n761), .B2(G317), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT52), .Z(new_n1038));
  OAI211_X1 g0838(.A(new_n1036), .B(new_n1038), .C1(new_n589), .C2(new_n763), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n739), .A2(G322), .B1(G283), .B2(new_n772), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT112), .Z(new_n1041));
  NAND2_X1  g0841(.A1(new_n758), .A2(G77), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n747), .A2(G50), .B1(G87), .B2(new_n774), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n745), .A2(new_n1001), .B1(G68), .B2(new_n772), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .A4(new_n306), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n744), .A2(G159), .B1(new_n761), .B2(G150), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT51), .Z(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n812), .B2(new_n938), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n1039), .A2(new_n1041), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n733), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n734), .B1(new_n465), .B2(new_n211), .C1(new_n997), .C2(new_n242), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1050), .A2(new_n718), .A3(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n959), .B2(new_n732), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n981), .A2(KEYINPUT111), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(new_n982), .Z(new_n1055));
  AOI21_X1  g0855(.A(new_n1053), .B1(new_n1055), .B2(new_n717), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1055), .A2(new_n991), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n991), .A2(new_n983), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n714), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1056), .B1(new_n1057), .B2(new_n1059), .ZN(G390));
  NAND2_X1  g0860(.A1(new_n897), .A2(new_n900), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n902), .A2(new_n835), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n898), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n685), .A2(new_n795), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1065), .A2(new_n786), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n835), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NOR3_X1   g0868(.A1(new_n1068), .A2(new_n882), .A3(new_n899), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n706), .A2(new_n707), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1071), .A2(G330), .A3(new_n794), .A4(new_n835), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1064), .A2(new_n1070), .A3(new_n1072), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n688), .B(new_n836), .C1(new_n840), .C2(new_n707), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n897), .A2(new_n900), .B1(new_n898), .B2(new_n1062), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1074), .B1(new_n1075), .B2(new_n1069), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n447), .B(G330), .C1(new_n867), .C2(new_n868), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n890), .A2(new_n623), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n835), .B1(new_n708), .B2(new_n794), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n902), .B1(new_n1080), .B2(new_n1074), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n688), .B(new_n795), .C1(new_n840), .C2(new_n707), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1072), .B(new_n1066), .C1(new_n1082), .C2(new_n835), .ZN(new_n1083));
  AOI211_X1 g0883(.A(KEYINPUT113), .B(new_n1079), .C1(new_n1081), .C2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT113), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1079), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1084), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n672), .B1(new_n1077), .B2(new_n1089), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1088), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1086), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1091), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1090), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1061), .A2(new_n728), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n718), .B1(new_n825), .B2(new_n1001), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT53), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n752), .A2(new_n363), .ZN(new_n1100));
  INV_X1    g0900(.A(G132), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n257), .B1(new_n1099), .B2(new_n1100), .C1(new_n802), .C2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n758), .A2(G159), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n739), .A2(G125), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n748), .A2(new_n937), .B1(new_n366), .B2(new_n755), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(KEYINPUT54), .B(G143), .ZN(new_n1107));
  INV_X1    g0907(.A(G128), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n814), .A2(new_n1107), .B1(new_n1108), .B2(new_n754), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .A4(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n753), .A2(new_n257), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(G107), .A2(new_n747), .B1(new_n744), .B2(G116), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n745), .A2(G97), .B1(new_n761), .B2(G283), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1042), .A2(new_n1112), .A3(new_n1113), .A4(new_n1114), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n739), .A2(G294), .B1(G68), .B2(new_n774), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT114), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1111), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1098), .B1(new_n1118), .B2(new_n733), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1091), .A2(new_n717), .B1(new_n1097), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1096), .A2(new_n1120), .ZN(G378));
  NAND2_X1  g0921(.A1(new_n369), .A2(new_n848), .ZN(new_n1122));
  XOR2_X1   g0922(.A(new_n1122), .B(KEYINPUT55), .Z(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n383), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n383), .A2(new_n1124), .ZN(new_n1127));
  XOR2_X1   g0927(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n1126), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  OR2_X1    g0930(.A1(new_n383), .A2(new_n1124), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1128), .B1(new_n1131), .B2(new_n1125), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n728), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n718), .B1(new_n825), .B2(G50), .ZN(new_n1135));
  AOI211_X1 g0935(.A(G41), .B(new_n306), .C1(new_n739), .C2(G283), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n755), .A2(new_n272), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G116), .B2(new_n761), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n1139), .B1(new_n748), .B2(new_n465), .C1(new_n433), .C2(new_n802), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n814), .A2(new_n424), .B1(new_n385), .B2(new_n752), .ZN(new_n1141));
  NOR4_X1   g0941(.A1(new_n1137), .A2(new_n1140), .A3(new_n931), .A4(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1142), .A2(KEYINPUT58), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n260), .A2(new_n671), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT115), .ZN(new_n1145));
  AOI211_X1 g0945(.A(G50), .B(new_n1145), .C1(new_n671), .C2(new_n282), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1147));
  XOR2_X1   g0947(.A(new_n1147), .B(KEYINPUT116), .Z(new_n1148));
  NOR2_X1   g0948(.A1(new_n752), .A2(new_n1107), .ZN(new_n1149));
  XOR2_X1   g0949(.A(new_n1149), .B(KEYINPUT117), .Z(new_n1150));
  NAND2_X1  g0950(.A1(new_n758), .A2(G150), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n747), .A2(G132), .B1(new_n761), .B2(G125), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(G128), .A2(new_n744), .B1(new_n745), .B2(G137), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  OR2_X1    g0954(.A1(new_n1154), .A2(KEYINPUT59), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n739), .A2(G124), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1156), .B(new_n1145), .C1(new_n813), .C2(new_n755), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n1154), .B2(KEYINPUT59), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n1142), .A2(KEYINPUT58), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1148), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1135), .B1(new_n1160), .B2(new_n733), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1134), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n884), .A2(G330), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n1133), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1133), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n884), .A2(G330), .A3(new_n1166), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1165), .A2(new_n901), .A3(new_n905), .A4(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1166), .B1(new_n884), .B2(G330), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n688), .B(new_n1133), .C1(new_n865), .C2(new_n883), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n906), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1168), .A2(new_n1171), .A3(KEYINPUT119), .ZN(new_n1172));
  NOR3_X1   g0972(.A1(new_n906), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT119), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  AND2_X1   g0975(.A1(new_n1172), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1163), .B1(new_n1176), .B2(new_n717), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1087), .B1(new_n1077), .B2(new_n1089), .ZN(new_n1178));
  AOI21_X1  g0978(.A(KEYINPUT57), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1079), .B1(new_n1091), .B2(new_n1094), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(KEYINPUT57), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n714), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1177), .B1(new_n1179), .B2(new_n1183), .ZN(G375));
  NAND2_X1  g0984(.A1(new_n1067), .A2(new_n728), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n718), .B1(new_n825), .B2(G68), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n748), .A2(new_n1107), .B1(new_n814), .B2(new_n363), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n802), .A2(new_n937), .B1(new_n754), .B2(new_n1101), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n306), .B1(new_n272), .B2(new_n755), .C1(new_n813), .C2(new_n752), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1190), .B1(new_n366), .B2(new_n763), .C1(new_n1108), .C2(new_n938), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n802), .A2(new_n807), .B1(new_n754), .B2(new_n764), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(G97), .B2(new_n772), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1193), .A2(new_n264), .A3(new_n932), .A4(new_n1011), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n507), .A2(new_n747), .B1(new_n745), .B2(G107), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT120), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n1195), .A2(new_n1196), .B1(new_n739), .B2(G303), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n1196), .B2(new_n1195), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1191), .B1(new_n1194), .B2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1186), .B1(new_n1199), .B2(new_n733), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n1086), .A2(new_n717), .B1(new_n1185), .B2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1081), .A2(new_n1079), .A3(new_n1083), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n987), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1201), .B1(new_n1094), .B2(new_n1204), .ZN(G381));
  OR2_X1    g1005(.A1(G390), .A2(G384), .ZN(new_n1206));
  OR2_X1    g1006(.A1(G393), .A2(G396), .ZN(new_n1207));
  OR4_X1    g1007(.A1(G387), .A2(new_n1206), .A3(G381), .A4(new_n1207), .ZN(new_n1208));
  XOR2_X1   g1008(.A(G375), .B(KEYINPUT121), .Z(new_n1209));
  OR3_X1    g1009(.A1(new_n1208), .A2(new_n1209), .A3(G378), .ZN(G407));
  AND2_X1   g1010(.A1(new_n1096), .A2(new_n1120), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n655), .A2(G213), .ZN(new_n1212));
  XOR2_X1   g1012(.A(new_n1212), .B(KEYINPUT122), .Z(new_n1213));
  NAND2_X1  g1013(.A1(new_n1211), .A2(new_n1213), .ZN(new_n1214));
  OAI211_X1 g1014(.A(G407), .B(G213), .C1(new_n1209), .C2(new_n1214), .ZN(G409));
  NOR2_X1   g1015(.A1(G390), .A2(new_n989), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(G393), .B(G396), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(G390), .A2(new_n989), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1217), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1220), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1218), .B1(new_n1222), .B2(new_n1216), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1221), .A2(new_n1223), .ZN(new_n1224));
  OAI211_X1 g1024(.A(G378), .B(new_n1177), .C1(new_n1179), .C2(new_n1183), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1178), .A2(new_n1203), .A3(new_n1175), .A4(new_n1172), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT123), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n716), .B1(new_n1168), .B2(new_n1171), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1227), .B1(new_n1228), .B2(new_n1163), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1181), .A2(new_n717), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1230), .A2(KEYINPUT123), .A3(new_n1162), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1226), .A2(new_n1229), .A3(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n1211), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1213), .B1(new_n1225), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT60), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1202), .B1(new_n1094), .B2(new_n1235), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1081), .A2(new_n1079), .A3(new_n1083), .A4(KEYINPUT60), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT125), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n672), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1236), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n1201), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n829), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1242), .A2(G384), .A3(new_n1201), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT62), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  AND2_X1   g1048(.A1(new_n1234), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1225), .A2(new_n1233), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT124), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1246), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1225), .A2(new_n1233), .A3(KEYINPUT124), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1252), .A2(new_n1212), .A3(new_n1253), .A4(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1249), .B1(new_n1255), .B2(new_n1247), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT61), .ZN(new_n1257));
  INV_X1    g1057(.A(G2897), .ZN(new_n1258));
  NOR3_X1   g1058(.A1(new_n1246), .A2(new_n1258), .A3(new_n1212), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n1244), .A2(new_n1245), .B1(G2897), .B2(new_n1213), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1257), .B1(new_n1261), .B2(new_n1234), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1224), .B1(new_n1256), .B2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1252), .A2(new_n1212), .A3(new_n1254), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n1260), .B2(new_n1259), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT63), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1255), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1234), .A2(KEYINPUT63), .A3(new_n1253), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1224), .A2(KEYINPUT61), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1265), .A2(new_n1267), .A3(new_n1268), .A4(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1263), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(KEYINPUT126), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT126), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1263), .A2(new_n1273), .A3(new_n1270), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1272), .A2(new_n1274), .ZN(G405));
  INV_X1    g1075(.A(KEYINPUT127), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1246), .A2(new_n1276), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(new_n1224), .B(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(G375), .A2(new_n1211), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n1279), .B(new_n1225), .C1(new_n1276), .C2(new_n1246), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(new_n1278), .B(new_n1280), .ZN(G402));
endmodule


