//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 0 1 1 0 1 1 1 0 0 0 1 0 0 1 1 1 1 1 1 1 0 1 0 0 0 0 0 0 1 0 0 1 1 0 0 0 1 1 0 1 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n210));
  NAND4_X1  g0010(.A1(new_n207), .A2(new_n208), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G1), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n211), .A2(new_n215), .ZN(new_n216));
  OR2_X1    g0016(.A1(new_n216), .A2(KEYINPUT1), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT65), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n215), .A2(G13), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n219), .B(G250), .C1(G257), .C2(G264), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT0), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(KEYINPUT64), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT64), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n224), .A2(G1), .A3(G13), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n227), .A2(new_n213), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n202), .A2(new_n203), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n221), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n218), .B(new_n232), .C1(KEYINPUT1), .C2(new_n216), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n242), .B(new_n243), .Z(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n223), .A2(new_n225), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(KEYINPUT66), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT66), .ZN(new_n252));
  NAND4_X1  g0052(.A1(new_n223), .A2(new_n225), .A3(new_n252), .A4(new_n249), .ZN(new_n253));
  AND2_X1   g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(G20), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n256), .A2(G77), .B1(G20), .B2(new_n203), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n257), .B1(new_n201), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n254), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(new_n261), .B(KEYINPUT11), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n212), .A2(G13), .A3(G20), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT69), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT69), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n254), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n213), .A2(G1), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(new_n203), .ZN(new_n272));
  OAI21_X1  g0072(.A(KEYINPUT12), .B1(new_n268), .B2(G68), .ZN(new_n273));
  INV_X1    g0073(.A(G13), .ZN(new_n274));
  NOR3_X1   g0074(.A1(new_n274), .A2(KEYINPUT12), .A3(G1), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(G20), .A3(new_n203), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n270), .A2(new_n272), .B1(new_n273), .B2(new_n276), .ZN(new_n277));
  AND2_X1   g0077(.A1(new_n262), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT3), .B(G33), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G232), .A3(G1698), .ZN(new_n280));
  INV_X1    g0080(.A(G1698), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(G226), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G97), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n280), .B(new_n282), .C1(new_n255), .C2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G33), .A2(G41), .ZN(new_n285));
  AND2_X1   g0085(.A1(new_n226), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n212), .B1(G41), .B2(G45), .ZN(new_n288));
  INV_X1    g0088(.A(G274), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OR2_X1    g0090(.A1(new_n290), .A2(KEYINPUT70), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(KEYINPUT70), .ZN(new_n292));
  INV_X1    g0092(.A(new_n222), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n285), .ZN(new_n294));
  AND2_X1   g0094(.A1(new_n294), .A2(new_n288), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n291), .A2(new_n292), .B1(G238), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT13), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n287), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n297), .B1(new_n287), .B2(new_n296), .ZN(new_n300));
  OAI21_X1  g0100(.A(G200), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n300), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n302), .A2(G190), .A3(new_n298), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n278), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT71), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n304), .B(new_n305), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n258), .ZN(new_n307));
  XOR2_X1   g0107(.A(KEYINPUT8), .B(G58), .Z(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n256), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n307), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n254), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n251), .A2(new_n253), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n271), .A2(new_n201), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n313), .A2(new_n263), .A3(new_n314), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n312), .B(new_n315), .C1(G50), .C2(new_n263), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n316), .B(KEYINPUT9), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n279), .A2(G222), .A3(new_n281), .ZN(new_n318));
  INV_X1    g0118(.A(G77), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n279), .A2(G1698), .ZN(new_n320));
  INV_X1    g0120(.A(G223), .ZN(new_n321));
  OAI221_X1 g0121(.A(new_n318), .B1(new_n319), .B2(new_n279), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n286), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n290), .B1(new_n295), .B2(G226), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G190), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G200), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n328), .B1(new_n323), .B2(new_n324), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n317), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT10), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT10), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n317), .A2(new_n330), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n262), .A2(new_n277), .ZN(new_n336));
  XNOR2_X1  g0136(.A(new_n336), .B(KEYINPUT72), .ZN(new_n337));
  OAI21_X1  g0137(.A(G169), .B1(new_n299), .B2(new_n300), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT14), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT14), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n340), .B(G169), .C1(new_n299), .C2(new_n300), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n302), .A2(G179), .A3(new_n298), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n339), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n337), .A2(new_n343), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n308), .A2(new_n258), .B1(G20), .B2(G77), .ZN(new_n345));
  XNOR2_X1  g0145(.A(KEYINPUT15), .B(G87), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n347), .A2(KEYINPUT67), .A3(new_n256), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT67), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(new_n346), .B2(new_n310), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n345), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n254), .ZN(new_n352));
  XNOR2_X1  g0152(.A(new_n352), .B(KEYINPUT68), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n271), .A2(new_n319), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n270), .A2(new_n354), .B1(new_n319), .B2(new_n269), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n279), .A2(G232), .A3(new_n281), .ZN(new_n357));
  INV_X1    g0157(.A(G107), .ZN(new_n358));
  INV_X1    g0158(.A(G238), .ZN(new_n359));
  OAI221_X1 g0159(.A(new_n357), .B1(new_n358), .B2(new_n279), .C1(new_n320), .C2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n286), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n290), .B1(new_n295), .B2(G244), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n363), .A2(G179), .ZN(new_n364));
  AOI21_X1  g0164(.A(G169), .B1(new_n361), .B2(new_n362), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n356), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G169), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n325), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(G179), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n323), .A2(new_n371), .A3(new_n324), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n370), .A2(new_n316), .A3(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n363), .A2(G200), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n326), .B2(new_n363), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n356), .A2(new_n376), .ZN(new_n377));
  NOR3_X1   g0177(.A1(new_n368), .A2(new_n374), .A3(new_n377), .ZN(new_n378));
  AND4_X1   g0178(.A1(new_n306), .A2(new_n335), .A3(new_n344), .A4(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT74), .ZN(new_n380));
  AND3_X1   g0180(.A1(KEYINPUT73), .A2(G58), .A3(G68), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT73), .B1(G58), .B2(G68), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n213), .B1(new_n383), .B2(new_n230), .ZN(new_n384));
  INV_X1    g0184(.A(G159), .ZN(new_n385));
  NOR3_X1   g0185(.A1(new_n385), .A2(G20), .A3(G33), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n380), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(G58), .A2(G68), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT73), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(KEYINPUT73), .A2(G58), .A3(G68), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(new_n230), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(G20), .ZN(new_n393));
  INV_X1    g0193(.A(new_n386), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n393), .A2(KEYINPUT74), .A3(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(KEYINPUT7), .B1(new_n279), .B2(G20), .ZN(new_n396));
  AND2_X1   g0196(.A1(KEYINPUT3), .A2(G33), .ZN(new_n397));
  NOR2_X1   g0197(.A1(KEYINPUT3), .A2(G33), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT7), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(new_n400), .A3(new_n213), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n396), .A2(new_n401), .A3(G68), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n387), .A2(new_n395), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT75), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n387), .A2(new_n395), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT16), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n403), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(KEYINPUT74), .B1(new_n393), .B2(new_n394), .ZN(new_n408));
  AOI211_X1 g0208(.A(new_n380), .B(new_n386), .C1(new_n392), .C2(G20), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n410), .B(new_n402), .C1(new_n404), .C2(KEYINPUT16), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n407), .A2(new_n411), .A3(new_n254), .ZN(new_n412));
  NOR4_X1   g0212(.A1(new_n254), .A2(new_n264), .A3(new_n309), .A4(new_n271), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n413), .B1(new_n264), .B2(new_n309), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n290), .B1(new_n295), .B2(G232), .ZN(new_n415));
  INV_X1    g0215(.A(G226), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(G1698), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(G223), .B2(G1698), .ZN(new_n418));
  INV_X1    g0218(.A(G87), .ZN(new_n419));
  OAI22_X1  g0219(.A1(new_n418), .A2(new_n399), .B1(new_n255), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n286), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n415), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n328), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(G190), .B2(new_n422), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n412), .A2(new_n414), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT17), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n412), .A2(KEYINPUT17), .A3(new_n414), .A4(new_n424), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n412), .A2(new_n414), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n422), .A2(new_n371), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n369), .B1(new_n421), .B2(new_n415), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT18), .B1(new_n430), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT76), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n430), .A2(KEYINPUT18), .A3(new_n434), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n430), .A2(KEYINPUT76), .A3(KEYINPUT18), .A4(new_n434), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n429), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n379), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(G45), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n442), .A2(G1), .ZN(new_n443));
  AND2_X1   g0243(.A1(KEYINPUT5), .A2(G41), .ZN(new_n444));
  NOR2_X1   g0244(.A1(KEYINPUT5), .A2(G41), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n222), .B1(G33), .B2(G41), .ZN(new_n447));
  NOR3_X1   g0247(.A1(new_n446), .A2(new_n447), .A3(new_n289), .ZN(new_n448));
  XNOR2_X1  g0248(.A(KEYINPUT5), .B(G41), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n449), .A2(new_n443), .B1(new_n293), .B2(new_n285), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n448), .B1(G270), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n279), .A2(G264), .A3(G1698), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n279), .A2(G257), .A3(new_n281), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n399), .A2(G303), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n286), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n369), .B1(new_n451), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT85), .ZN(new_n458));
  AOI21_X1  g0258(.A(G20), .B1(G33), .B2(G283), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n255), .A2(G97), .ZN(new_n460));
  INV_X1    g0260(.A(G116), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n459), .A2(new_n460), .B1(G20), .B2(new_n461), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n462), .A2(new_n250), .A3(KEYINPUT20), .ZN(new_n463));
  AOI21_X1  g0263(.A(KEYINPUT20), .B1(new_n462), .B2(new_n250), .ZN(new_n464));
  OAI22_X1  g0264(.A1(new_n463), .A2(new_n464), .B1(G116), .B2(new_n268), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT84), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n255), .A2(G1), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(new_n461), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n313), .A2(new_n268), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n465), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n313), .A2(KEYINPUT84), .A3(new_n268), .A4(new_n468), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n458), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n469), .A2(new_n466), .ZN(new_n473));
  INV_X1    g0273(.A(new_n464), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n462), .A2(new_n250), .A3(KEYINPUT20), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n474), .A2(new_n475), .B1(new_n269), .B2(new_n461), .ZN(new_n476));
  AND4_X1   g0276(.A1(new_n458), .A2(new_n473), .A3(new_n476), .A4(new_n471), .ZN(new_n477));
  OAI211_X1 g0277(.A(KEYINPUT21), .B(new_n457), .C1(new_n472), .C2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n451), .A2(new_n456), .A3(G179), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n480), .B1(new_n472), .B2(new_n477), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n470), .A2(new_n458), .A3(new_n471), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n473), .A2(new_n476), .A3(new_n471), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT85), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(KEYINPUT21), .B1(new_n486), .B2(new_n457), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n451), .A2(new_n456), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G200), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n489), .B1(new_n326), .B2(new_n488), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  NOR3_X1   g0291(.A1(new_n482), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT83), .ZN(new_n493));
  OAI211_X1 g0293(.A(G244), .B(new_n281), .C1(new_n397), .C2(new_n398), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n279), .A2(KEYINPUT4), .A3(G244), .A4(new_n281), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G33), .A2(G283), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n279), .A2(G250), .A3(G1698), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n496), .A2(new_n497), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n286), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n294), .A2(new_n449), .A3(G274), .A4(new_n443), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n446), .A2(new_n294), .ZN(new_n503));
  INV_X1    g0303(.A(G257), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT79), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n505), .B1(new_n500), .B2(new_n286), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(KEYINPUT79), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n509), .A2(G190), .A3(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n467), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n313), .A2(G97), .A3(new_n263), .A4(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n263), .A2(G97), .ZN(new_n515));
  XNOR2_X1  g0315(.A(new_n515), .B(KEYINPUT78), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  AND3_X1   g0317(.A1(new_n396), .A2(new_n401), .A3(G107), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n358), .A2(KEYINPUT6), .A3(G97), .ZN(new_n519));
  XNOR2_X1  g0319(.A(G97), .B(G107), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT6), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OAI22_X1  g0322(.A1(new_n522), .A2(new_n213), .B1(new_n319), .B2(new_n259), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n254), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT77), .ZN(new_n525));
  AND2_X1   g0325(.A1(G97), .A2(G107), .ZN(new_n526));
  NOR2_X1   g0326(.A1(G97), .A2(G107), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n521), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n358), .A2(KEYINPUT6), .A3(G97), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n530), .A2(G20), .B1(G77), .B2(new_n258), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n396), .A2(new_n401), .A3(G107), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT77), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n533), .A2(new_n534), .A3(new_n254), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n517), .B1(new_n525), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n507), .A2(G200), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n512), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n501), .A2(KEYINPUT79), .A3(new_n506), .ZN(new_n539));
  AOI21_X1  g0339(.A(KEYINPUT79), .B1(new_n501), .B2(new_n506), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n369), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n507), .A2(G179), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n517), .ZN(new_n544));
  AOI211_X1 g0344(.A(KEYINPUT77), .B(new_n313), .C1(new_n531), .C2(new_n532), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n534), .B1(new_n533), .B2(new_n254), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n541), .A2(new_n543), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n538), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n443), .A2(G274), .ZN(new_n550));
  OAI21_X1  g0350(.A(G250), .B1(new_n442), .B2(G1), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n550), .B1(new_n447), .B2(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(G244), .B(G1698), .C1(new_n397), .C2(new_n398), .ZN(new_n553));
  OAI211_X1 g0353(.A(G238), .B(new_n281), .C1(new_n397), .C2(new_n398), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G33), .A2(G116), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n552), .B1(new_n556), .B2(new_n286), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n557), .A2(new_n369), .ZN(new_n558));
  AOI211_X1 g0358(.A(new_n371), .B(new_n552), .C1(new_n556), .C2(new_n286), .ZN(new_n559));
  OAI21_X1  g0359(.A(KEYINPUT80), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AOI211_X1 g0360(.A(new_n264), .B(new_n467), .C1(new_n251), .C2(new_n253), .ZN(new_n561));
  XNOR2_X1  g0361(.A(new_n346), .B(KEYINPUT82), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT19), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n310), .B2(new_n283), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n279), .A2(new_n213), .A3(G68), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n568));
  AND2_X1   g0368(.A1(new_n568), .A2(new_n213), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n419), .A2(new_n283), .A3(new_n358), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(KEYINPUT81), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT81), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n572), .A2(new_n419), .A3(new_n283), .A4(new_n358), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n569), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n251), .B(new_n253), .C1(new_n567), .C2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n269), .A2(new_n346), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n563), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n557), .A2(G179), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT80), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n578), .B(new_n579), .C1(new_n369), .C2(new_n557), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n560), .A2(new_n577), .A3(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n557), .A2(new_n328), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n582), .B1(G190), .B2(new_n557), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n313), .A2(G87), .A3(new_n263), .A4(new_n513), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n575), .A2(new_n584), .A3(new_n576), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n493), .B1(new_n549), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n557), .A2(G190), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(new_n328), .B2(new_n557), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n591), .A2(new_n585), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n578), .B1(new_n369), .B2(new_n557), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n571), .A2(new_n573), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n566), .B(new_n565), .C1(new_n594), .C2(new_n569), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n595), .A2(new_n254), .B1(new_n269), .B2(new_n346), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n593), .A2(KEYINPUT80), .B1(new_n596), .B2(new_n563), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n592), .B1(new_n597), .B2(new_n580), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n598), .A2(new_n538), .A3(new_n548), .A4(KEYINPUT83), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n213), .B(G87), .C1(new_n397), .C2(new_n398), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT22), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT22), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n279), .A2(new_n602), .A3(new_n213), .A4(G87), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT24), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n555), .A2(G20), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT23), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n607), .B1(new_n213), .B2(G107), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n358), .A2(KEYINPUT23), .A3(G20), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n606), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n604), .A2(new_n605), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n605), .B1(new_n604), .B2(new_n610), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n254), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n264), .A2(new_n358), .ZN(new_n614));
  XNOR2_X1  g0414(.A(new_n614), .B(KEYINPUT25), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n615), .B1(new_n561), .B2(G107), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  OAI211_X1 g0417(.A(G250), .B(new_n281), .C1(new_n397), .C2(new_n398), .ZN(new_n618));
  OAI211_X1 g0418(.A(G257), .B(G1698), .C1(new_n397), .C2(new_n398), .ZN(new_n619));
  NAND2_X1  g0419(.A1(G33), .A2(G294), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n621), .A2(new_n286), .B1(new_n450), .B2(G264), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n622), .A2(new_n371), .A3(new_n502), .ZN(new_n623));
  AOI21_X1  g0423(.A(G169), .B1(new_n622), .B2(new_n502), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n617), .A2(KEYINPUT86), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(KEYINPUT86), .B1(new_n617), .B2(new_n625), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n622), .A2(new_n502), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(G200), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n622), .A2(G190), .A3(new_n502), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n617), .A2(new_n631), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n626), .A2(new_n627), .A3(new_n632), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n599), .A2(new_n633), .ZN(new_n634));
  AND4_X1   g0434(.A1(new_n441), .A2(new_n492), .A3(new_n589), .A4(new_n634), .ZN(G372));
  INV_X1    g0435(.A(KEYINPUT87), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n335), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n332), .A2(KEYINPUT87), .A3(new_n334), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n430), .A2(new_n434), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT18), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n437), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n337), .A2(new_n343), .B1(new_n368), .B2(new_n304), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n643), .B1(new_n644), .B2(new_n429), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n374), .B1(new_n639), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n441), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n457), .B1(new_n472), .B2(new_n477), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT21), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n617), .A2(new_n625), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n650), .A2(new_n478), .A3(new_n481), .A4(new_n651), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n583), .A2(new_n586), .B1(new_n577), .B2(new_n593), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n653), .B1(new_n617), .B2(new_n631), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n549), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(KEYINPUT26), .B1(new_n548), .B2(new_n588), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n577), .A2(new_n593), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n536), .A2(new_n542), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT26), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n659), .A2(new_n653), .A3(new_n660), .A4(new_n541), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n657), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n646), .B1(new_n647), .B2(new_n663), .ZN(G369));
  OR3_X1    g0464(.A1(new_n482), .A2(new_n487), .A3(new_n491), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n665), .A2(KEYINPUT89), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n274), .A2(G20), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n212), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n668), .B(KEYINPUT88), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n670), .A2(G213), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(G343), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n486), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n665), .B2(KEYINPUT89), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n482), .A2(new_n487), .ZN(new_n677));
  OAI22_X1  g0477(.A1(new_n666), .A2(new_n676), .B1(new_n677), .B2(new_n675), .ZN(new_n678));
  XNOR2_X1  g0478(.A(KEYINPUT90), .B(G330), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n674), .A2(new_n617), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n633), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n674), .A2(new_n617), .A3(new_n625), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n677), .A2(new_n674), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n633), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n673), .A2(new_n617), .A3(new_n625), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n686), .A2(new_n690), .ZN(G399));
  INV_X1    g0491(.A(new_n219), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G41), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n594), .A2(new_n461), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n694), .A2(G1), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n231), .B2(new_n694), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n626), .A2(new_n627), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n700), .A2(new_n650), .A3(new_n478), .A4(new_n481), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n655), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n598), .A2(new_n660), .A3(new_n541), .A4(new_n659), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n587), .A2(new_n658), .ZN(new_n704));
  OAI21_X1  g0504(.A(KEYINPUT26), .B1(new_n548), .B2(new_n704), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n703), .A2(new_n658), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n674), .B1(new_n702), .B2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT29), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n674), .B1(new_n656), .B2(new_n662), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n708), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n634), .A2(new_n492), .A3(new_n589), .A4(new_n673), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n622), .A2(new_n557), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n479), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n715), .A2(new_n509), .A3(new_n511), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT30), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n557), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n488), .A2(new_n371), .A3(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT91), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n628), .ZN(new_n723));
  OAI21_X1  g0523(.A(KEYINPUT92), .B1(new_n723), .B2(new_n510), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT92), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n507), .A2(new_n725), .A3(new_n628), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n488), .A2(new_n719), .A3(KEYINPUT91), .A4(new_n371), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n722), .A2(new_n724), .A3(new_n726), .A4(new_n727), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n715), .A2(new_n509), .A3(KEYINPUT30), .A4(new_n511), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n718), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(new_n674), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT31), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n673), .A2(new_n732), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n718), .A2(new_n728), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n729), .B1(new_n735), .B2(KEYINPUT93), .ZN(new_n736));
  AND3_X1   g0536(.A1(new_n718), .A2(new_n728), .A3(KEYINPUT93), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n734), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n713), .A2(new_n733), .A3(new_n738), .ZN(new_n739));
  AOI211_X1 g0539(.A(new_n709), .B(new_n712), .C1(new_n679), .C2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n699), .B1(new_n740), .B2(G1), .ZN(G364));
  AOI21_X1  g0541(.A(new_n212), .B1(new_n667), .B2(G45), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n693), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n681), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n745), .B1(new_n679), .B2(new_n678), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n219), .A2(new_n279), .ZN(new_n747));
  INV_X1    g0547(.A(G355), .ZN(new_n748));
  OAI22_X1  g0548(.A1(new_n747), .A2(new_n748), .B1(G116), .B2(new_n219), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n219), .A2(new_n399), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT94), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n231), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n752), .B1(new_n442), .B2(new_n753), .ZN(new_n754));
  OR2_X1    g0554(.A1(new_n244), .A2(new_n442), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n749), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n227), .B1(G20), .B2(new_n369), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G13), .A2(G33), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G20), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n744), .B1(new_n756), .B2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n757), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n213), .A2(new_n326), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n371), .A2(G200), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  XOR2_X1   g0567(.A(new_n767), .B(KEYINPUT95), .Z(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n371), .A2(G200), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT96), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(new_n765), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n769), .A2(G58), .B1(G87), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n371), .A2(new_n328), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n765), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n279), .B1(new_n776), .B2(new_n201), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n213), .A2(G190), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n766), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n779), .A2(new_n203), .B1(new_n780), .B2(new_n319), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G179), .A2(G200), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n213), .B1(new_n782), .B2(G190), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n777), .B(new_n781), .C1(G97), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n771), .A2(new_n778), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G107), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n778), .A2(new_n782), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n385), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT32), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n774), .A2(new_n785), .A3(new_n788), .A4(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G294), .ZN(new_n793));
  INV_X1    g0593(.A(G326), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n399), .B1(new_n783), .B2(new_n793), .C1(new_n776), .C2(new_n794), .ZN(new_n795));
  XOR2_X1   g0595(.A(KEYINPUT33), .B(G317), .Z(new_n796));
  INV_X1    g0596(.A(G322), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n796), .A2(new_n779), .B1(new_n767), .B2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G311), .ZN(new_n799));
  INV_X1    g0599(.A(G329), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n780), .A2(new_n799), .B1(new_n789), .B2(new_n800), .ZN(new_n801));
  NOR3_X1   g0601(.A1(new_n795), .A2(new_n798), .A3(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G283), .ZN(new_n803));
  INV_X1    g0603(.A(G303), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n802), .B1(new_n803), .B2(new_n786), .C1(new_n804), .C2(new_n772), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n764), .B1(new_n792), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n763), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n760), .B(KEYINPUT97), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n807), .B1(new_n678), .B2(new_n808), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n746), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(G396));
  AOI21_X1  g0611(.A(new_n673), .B1(new_n353), .B2(new_n355), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n367), .B1(new_n377), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n356), .A2(new_n366), .A3(new_n673), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n710), .B(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n739), .A2(new_n679), .ZN(new_n818));
  OR3_X1    g0618(.A1(new_n817), .A2(KEYINPUT101), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(KEYINPUT101), .B1(new_n817), .B2(new_n818), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n744), .B1(new_n817), .B2(new_n818), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n744), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n757), .A2(new_n758), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n823), .B1(new_n824), .B2(new_n319), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n780), .A2(new_n385), .ZN(new_n826));
  INV_X1    g0626(.A(G137), .ZN(new_n827));
  INV_X1    g0627(.A(G150), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n776), .A2(new_n827), .B1(new_n779), .B2(new_n828), .ZN(new_n829));
  XOR2_X1   g0629(.A(KEYINPUT99), .B(G143), .Z(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n826), .B(new_n829), .C1(new_n769), .C2(new_n831), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(KEYINPUT34), .ZN(new_n833));
  INV_X1    g0633(.A(G132), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n279), .B1(new_n789), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(G58), .B2(new_n784), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n836), .B1(new_n201), .B2(new_n772), .C1(new_n203), .C2(new_n786), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n787), .A2(G87), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n799), .B2(new_n789), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n839), .B(KEYINPUT98), .Z(new_n840));
  OAI22_X1  g0640(.A1(new_n776), .A2(new_n804), .B1(new_n779), .B2(new_n803), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n399), .B1(new_n783), .B2(new_n283), .C1(new_n793), .C2(new_n767), .ZN(new_n842));
  INV_X1    g0642(.A(new_n780), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n841), .B(new_n842), .C1(G116), .C2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n358), .B2(new_n772), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n833), .A2(new_n837), .B1(new_n840), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(KEYINPUT100), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n757), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n846), .A2(KEYINPUT100), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n825), .B1(new_n816), .B2(new_n759), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n822), .A2(new_n850), .ZN(G384));
  NOR2_X1   g0651(.A1(new_n667), .A2(new_n212), .ZN(new_n852));
  INV_X1    g0652(.A(new_n343), .ZN(new_n853));
  AND3_X1   g0653(.A1(new_n303), .A2(new_n262), .A3(new_n277), .ZN(new_n854));
  AOI21_X1  g0654(.A(KEYINPUT71), .B1(new_n854), .B2(new_n301), .ZN(new_n855));
  AND4_X1   g0655(.A1(KEYINPUT71), .A2(new_n278), .A3(new_n301), .A4(new_n303), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n853), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n337), .A2(new_n674), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n344), .A2(new_n858), .A3(new_n304), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n815), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n730), .A2(KEYINPUT31), .A3(new_n674), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT105), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n730), .A2(KEYINPUT105), .A3(KEYINPUT31), .A4(new_n674), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n713), .A2(new_n733), .A3(new_n867), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n862), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n430), .A2(new_n672), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT37), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n640), .A2(new_n870), .A3(new_n871), .A4(new_n425), .ZN(new_n872));
  INV_X1    g0672(.A(new_n425), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n403), .A2(new_n406), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n410), .A2(KEYINPUT16), .A3(new_n402), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n874), .A2(new_n875), .A3(new_n254), .ZN(new_n876));
  INV_X1    g0676(.A(new_n672), .ZN(new_n877));
  AOI22_X1  g0677(.A1(new_n414), .A2(new_n876), .B1(new_n877), .B2(new_n433), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT37), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n872), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n414), .A2(new_n876), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n672), .ZN(new_n882));
  OAI211_X1 g0682(.A(KEYINPUT38), .B(new_n880), .C1(new_n440), .C2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT104), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n429), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n427), .A2(KEYINPUT104), .A3(new_n428), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n885), .A2(new_n643), .A3(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n870), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n640), .A2(new_n870), .A3(new_n425), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT37), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n887), .A2(new_n888), .B1(new_n872), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n883), .B1(new_n891), .B2(KEYINPUT38), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n869), .A2(KEYINPUT40), .A3(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT38), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n437), .A2(new_n436), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n896), .A2(new_n439), .A3(new_n642), .ZN(new_n897));
  INV_X1    g0697(.A(new_n429), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n882), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n880), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n895), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n883), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT40), .B1(new_n869), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n894), .A2(new_n903), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n441), .A2(new_n868), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n679), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT106), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n906), .A2(new_n907), .ZN(new_n909));
  AOI211_X1 g0709(.A(new_n908), .B(new_n909), .C1(new_n905), .C2(new_n904), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT39), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n887), .A2(new_n888), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n890), .A2(new_n872), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT38), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n899), .A2(new_n900), .A3(new_n895), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n912), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n344), .A2(new_n674), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n901), .A2(new_n883), .A3(KEYINPUT39), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n643), .A2(new_n672), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n814), .B(KEYINPUT103), .Z(new_n922));
  AOI21_X1  g0722(.A(new_n922), .B1(new_n710), .B2(new_n816), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n860), .A2(new_n861), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n921), .B1(new_n926), .B2(new_n902), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n920), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n441), .B1(new_n712), .B2(new_n709), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n646), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n928), .B(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n852), .B1(new_n911), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n931), .B2(new_n911), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n228), .B(G116), .C1(KEYINPUT35), .C2(new_n530), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n934), .A2(KEYINPUT102), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(KEYINPUT102), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n530), .A2(KEYINPUT35), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT36), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n753), .A2(G77), .A3(new_n383), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(G50), .B2(new_n203), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n941), .A2(G1), .A3(new_n274), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n933), .A2(new_n939), .A3(new_n942), .ZN(G367));
  OAI211_X1 g0743(.A(new_n538), .B(new_n548), .C1(new_n536), .C2(new_n673), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT108), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n659), .A2(new_n541), .A3(new_n674), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n947), .A2(new_n633), .A3(new_n687), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n948), .A2(KEYINPUT42), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(KEYINPUT42), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n548), .B1(new_n945), .B2(new_n700), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n673), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n949), .A2(new_n950), .A3(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n673), .A2(new_n586), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n954), .A2(new_n593), .A3(new_n577), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n704), .B2(new_n954), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT107), .Z(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT109), .Z(new_n961));
  AND3_X1   g0761(.A1(new_n953), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n959), .B1(new_n953), .B2(new_n961), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n680), .B1(new_n683), .B2(new_n684), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n947), .ZN(new_n965));
  OR3_X1    g0765(.A1(new_n962), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n965), .B1(new_n962), .B2(new_n963), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n693), .B(KEYINPUT41), .Z(new_n968));
  AOI21_X1  g0768(.A(KEYINPUT45), .B1(new_n690), .B2(new_n947), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n688), .A2(new_n689), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n945), .A2(new_n946), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT45), .ZN(new_n972));
  NOR3_X1   g0772(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n969), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(KEYINPUT44), .B1(new_n970), .B2(new_n971), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT44), .ZN(new_n976));
  NOR3_X1   g0776(.A1(new_n690), .A2(new_n976), .A3(new_n947), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n974), .B(new_n686), .C1(new_n975), .C2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n688), .B1(new_n687), .B2(new_n685), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n680), .B(new_n979), .Z(new_n980));
  OAI22_X1  g0780(.A1(new_n975), .A2(new_n977), .B1(new_n969), .B2(new_n973), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n964), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n978), .A2(new_n740), .A3(new_n980), .A4(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n968), .B1(new_n983), .B2(new_n740), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n966), .B(new_n967), .C1(new_n984), .C2(new_n743), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n762), .B1(new_n692), .B2(new_n347), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n751), .A2(new_n240), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n823), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n787), .A2(G97), .ZN(new_n989));
  INV_X1    g0789(.A(G317), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n989), .B(new_n399), .C1(new_n990), .C2(new_n789), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT111), .ZN(new_n992));
  AOI21_X1  g0792(.A(KEYINPUT46), .B1(new_n773), .B2(G116), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT110), .Z(new_n994));
  NAND3_X1  g0794(.A1(new_n773), .A2(KEYINPUT46), .A3(G116), .ZN(new_n995));
  INV_X1    g0795(.A(new_n776), .ZN(new_n996));
  INV_X1    g0796(.A(new_n779), .ZN(new_n997));
  AOI22_X1  g0797(.A1(G311), .A2(new_n996), .B1(new_n997), .B2(G294), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(new_n358), .B2(new_n783), .C1(new_n803), .C2(new_n780), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(G303), .B2(new_n769), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n992), .A2(new_n994), .A3(new_n995), .A4(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT112), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n279), .B1(new_n783), .B2(new_n203), .C1(new_n828), .C2(new_n767), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n776), .A2(new_n830), .B1(new_n827), .B2(new_n789), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n779), .A2(new_n385), .B1(new_n780), .B2(new_n201), .ZN(new_n1005));
  NOR3_X1   g0805(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n787), .A2(G77), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1006), .B(new_n1007), .C1(new_n202), .C2(new_n772), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1002), .A2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT47), .Z(new_n1010));
  OAI221_X1 g0810(.A(new_n988), .B1(new_n808), .B2(new_n956), .C1(new_n1010), .C2(new_n764), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n985), .A2(new_n1011), .ZN(G387));
  OR2_X1    g0812(.A1(new_n685), .A2(new_n808), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n751), .B1(new_n237), .B2(new_n442), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n696), .B2(new_n747), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n442), .B1(new_n203), .B2(new_n319), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n308), .A2(new_n201), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1016), .B1(new_n1017), .B2(KEYINPUT50), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n696), .B(new_n1018), .C1(KEYINPUT50), .C2(new_n1017), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n1015), .A2(new_n1019), .B1(new_n358), .B2(new_n692), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n744), .B1(new_n1020), .B2(new_n762), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n309), .A2(new_n779), .B1(new_n203), .B2(new_n780), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n767), .A2(new_n201), .B1(new_n789), .B2(new_n828), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n279), .B1(new_n776), .B2(new_n385), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n773), .A2(G77), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n562), .A2(new_n784), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1025), .A2(new_n989), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n776), .A2(new_n797), .B1(new_n779), .B2(new_n799), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT113), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n804), .B2(new_n780), .C1(new_n990), .C2(new_n768), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT48), .ZN(new_n1032));
  AND2_X1   g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n772), .A2(new_n793), .B1(new_n803), .B2(new_n783), .ZN(new_n1035));
  NOR3_X1   g0835(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(KEYINPUT49), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n789), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n279), .B1(new_n1038), .B2(G326), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1037), .B(new_n1039), .C1(new_n461), .C2(new_n786), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1036), .A2(KEYINPUT49), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1028), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1021), .B1(new_n1042), .B2(new_n757), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n980), .A2(new_n743), .B1(new_n1013), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n980), .A2(new_n740), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n693), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n980), .A2(new_n740), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1044), .B1(new_n1046), .B2(new_n1047), .ZN(G393));
  NAND2_X1  g0848(.A1(new_n971), .A2(new_n760), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n1038), .A2(new_n831), .B1(new_n997), .B2(G50), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n399), .B1(new_n843), .B2(new_n308), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1050), .B(new_n1051), .C1(new_n319), .C2(new_n783), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT51), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n776), .A2(new_n828), .B1(new_n767), .B2(new_n385), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n773), .A2(G68), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1055), .B(new_n838), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n776), .A2(new_n990), .B1(new_n767), .B2(new_n799), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1057), .B(new_n1058), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1059), .B(new_n788), .C1(new_n803), .C2(new_n772), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G303), .A2(new_n997), .B1(new_n843), .B2(G294), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n279), .B1(new_n1038), .B2(G322), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1061), .B(new_n1062), .C1(new_n461), .C2(new_n783), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n1052), .A2(new_n1056), .B1(new_n1060), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n757), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n761), .B1(new_n283), .B2(new_n219), .C1(new_n752), .C2(new_n247), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1049), .A2(new_n744), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n978), .A2(new_n982), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1067), .B1(new_n1068), .B2(new_n742), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n983), .A2(new_n693), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1068), .A2(new_n1045), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1069), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(G390));
  NAND3_X1  g0873(.A1(new_n441), .A2(G330), .A3(new_n868), .ZN(new_n1074));
  AND3_X1   g0874(.A1(new_n929), .A2(new_n1074), .A3(new_n646), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n868), .A2(G330), .A3(new_n816), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n925), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n674), .B(new_n815), .C1(new_n702), .C2(new_n706), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1078), .A2(new_n922), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n739), .A2(new_n679), .A3(new_n924), .A4(new_n816), .ZN(new_n1080));
  AND3_X1   g0880(.A1(new_n1077), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n739), .A2(new_n679), .A3(new_n816), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n925), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n862), .A2(new_n868), .A3(G330), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n923), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1075), .B1(new_n1081), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n918), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n674), .B(new_n815), .C1(new_n656), .C2(new_n662), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n924), .B1(new_n1088), .B2(new_n922), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n917), .A2(new_n919), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n924), .B1(new_n1078), .B2(new_n922), .ZN(new_n1091));
  AND3_X1   g0891(.A1(new_n1091), .A2(new_n892), .A3(new_n1087), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1080), .ZN(new_n1093));
  NOR3_X1   g0893(.A1(new_n1090), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1087), .B1(new_n923), .B2(new_n925), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n429), .A2(new_n884), .B1(new_n642), .B2(new_n437), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n870), .B1(new_n1096), .B2(new_n886), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n914), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n895), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(KEYINPUT39), .B1(new_n1099), .B2(new_n883), .ZN(new_n1100));
  AND3_X1   g0900(.A1(new_n901), .A2(new_n883), .A3(KEYINPUT39), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1095), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1091), .A2(new_n892), .A3(new_n1087), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1084), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1086), .B1(new_n1094), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1084), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1102), .A2(new_n1103), .A3(new_n1080), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1077), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n869), .A2(G330), .B1(new_n1082), .B2(new_n925), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1109), .B1(new_n1110), .B2(new_n923), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1107), .A2(new_n1108), .A3(new_n1075), .A4(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1105), .A2(new_n693), .A3(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1107), .A2(new_n1108), .A3(new_n743), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n758), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n779), .A2(new_n358), .B1(new_n780), .B2(new_n283), .ZN(new_n1116));
  XOR2_X1   g0916(.A(new_n1116), .B(KEYINPUT115), .Z(new_n1117));
  OAI221_X1 g0917(.A(new_n1117), .B1(new_n203), .B2(new_n786), .C1(new_n419), .C2(new_n772), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n767), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(G283), .A2(new_n996), .B1(new_n1119), .B2(G116), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n279), .B1(new_n1038), .B2(G294), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1120), .B(new_n1121), .C1(new_n319), .C2(new_n783), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n773), .A2(G150), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT53), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n787), .A2(G50), .ZN(new_n1125));
  XOR2_X1   g0925(.A(KEYINPUT54), .B(G143), .Z(new_n1126));
  AOI22_X1  g0926(.A1(new_n996), .A2(G128), .B1(new_n843), .B2(new_n1126), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n997), .A2(G137), .B1(new_n1038), .B2(G125), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n279), .B1(new_n767), .B2(new_n834), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(G159), .B2(new_n784), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1125), .A2(new_n1127), .A3(new_n1128), .A4(new_n1130), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n1118), .A2(new_n1122), .B1(new_n1124), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n757), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n823), .B1(new_n824), .B2(new_n309), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1115), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  AND2_X1   g0935(.A1(new_n1114), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1113), .A2(new_n1136), .ZN(G378));
  NAND2_X1  g0937(.A1(new_n862), .A2(new_n868), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n883), .B2(new_n901), .ZN(new_n1139));
  OAI211_X1 g0939(.A(G330), .B(new_n893), .C1(new_n1139), .C2(KEYINPUT40), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n672), .A2(new_n316), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n639), .A2(new_n373), .A3(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n637), .A2(new_n373), .A3(new_n638), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1143), .A2(new_n316), .A3(new_n672), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1142), .A2(new_n1144), .A3(new_n1146), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  AND3_X1   g0950(.A1(new_n1150), .A2(new_n920), .A3(new_n927), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1150), .B1(new_n920), .B2(new_n927), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1140), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1150), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n928), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(G330), .ZN(new_n1156));
  NOR3_X1   g0956(.A1(new_n894), .A2(new_n903), .A3(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1150), .A2(new_n920), .A3(new_n927), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1155), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1153), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n743), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1150), .A2(new_n759), .ZN(new_n1162));
  INV_X1    g0962(.A(G41), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1163), .B(new_n399), .C1(new_n789), .C2(new_n803), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(G116), .A2(new_n996), .B1(new_n997), .B2(G97), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n358), .B2(new_n767), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1164), .B(new_n1166), .C1(G68), .C2(new_n784), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n562), .A2(new_n843), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n787), .A2(G58), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1167), .A2(new_n1026), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT58), .ZN(new_n1171));
  OR2_X1    g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n201), .B1(new_n397), .B2(G41), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n996), .A2(G125), .B1(new_n784), .B2(G150), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT116), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n773), .A2(new_n1126), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1119), .A2(G128), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(G132), .A2(new_n997), .B1(new_n843), .B2(G137), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n1181), .A2(KEYINPUT59), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1181), .A2(KEYINPUT59), .ZN(new_n1183));
  AOI211_X1 g0983(.A(G33), .B(G41), .C1(new_n1038), .C2(G124), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n385), .B2(new_n786), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(new_n1182), .A2(new_n1183), .A3(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n757), .B1(new_n1175), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n824), .A2(new_n201), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(new_n744), .A3(new_n1188), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1162), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1161), .A2(new_n1191), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1159), .A2(new_n1153), .B1(new_n1112), .B2(new_n1075), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n694), .B1(new_n1193), .B2(KEYINPUT57), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1112), .A2(new_n1075), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1160), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT57), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1192), .B1(new_n1194), .B2(new_n1198), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT117), .ZN(G375));
  NAND2_X1  g1000(.A1(new_n1111), .A2(new_n743), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n996), .A2(G132), .B1(new_n1038), .B2(G128), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n997), .A2(new_n1126), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n784), .A2(G50), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n399), .B1(new_n843), .B2(G150), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1169), .B1(new_n385), .B2(new_n772), .C1(new_n827), .C2(new_n768), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n779), .A2(new_n461), .B1(new_n780), .B2(new_n358), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT118), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1209), .B(new_n1027), .C1(new_n283), .C2(new_n772), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n279), .B1(new_n1038), .B2(G303), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(G294), .A2(new_n996), .B1(new_n1119), .B2(G283), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1007), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n1206), .A2(new_n1207), .B1(new_n1210), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n757), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n823), .B1(new_n824), .B2(new_n203), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(new_n924), .C2(new_n759), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1201), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n968), .B1(new_n1111), .B2(new_n1075), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1085), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n929), .A2(new_n1074), .A3(new_n646), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1221), .A2(new_n1222), .A3(new_n1109), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1220), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1219), .A2(new_n1224), .ZN(G381));
  INV_X1    g1025(.A(G375), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT119), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n1113), .A2(new_n1227), .A3(new_n1136), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1227), .B1(new_n1113), .B2(new_n1136), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n985), .A2(new_n1072), .A3(new_n1011), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NOR4_X1   g1032(.A1(G381), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1226), .A2(new_n1230), .A3(new_n1232), .A4(new_n1233), .ZN(G407));
  INV_X1    g1034(.A(G343), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(G213), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1226), .A2(new_n1230), .A3(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(G407), .A2(new_n1238), .A3(G213), .ZN(G409));
  AOI21_X1  g1039(.A(new_n1072), .B1(new_n985), .B2(new_n1011), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1241), .A2(KEYINPUT123), .A3(new_n1231), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT123), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n1232), .B2(new_n1240), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(G393), .B(new_n810), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1242), .A2(new_n1244), .A3(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT61), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1243), .B(new_n1245), .C1(new_n1232), .C2(new_n1240), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1247), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1190), .B1(new_n1160), .B2(new_n743), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n693), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1193), .A2(KEYINPUT57), .ZN(new_n1253));
  OAI211_X1 g1053(.A(G378), .B(new_n1251), .C1(new_n1252), .C2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1251), .B1(new_n968), .B2(new_n1196), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1229), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1113), .A2(new_n1136), .A3(new_n1227), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1255), .A2(new_n1256), .A3(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1254), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n1236), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1221), .A2(KEYINPUT60), .A3(new_n1222), .A4(new_n1109), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n693), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1086), .A2(KEYINPUT60), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1262), .B1(new_n1223), .B2(new_n1263), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n850), .B(new_n822), .C1(new_n1264), .C2(new_n1218), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1263), .A2(new_n1223), .ZN(new_n1266));
  OAI211_X1 g1066(.A(G384), .B(new_n1219), .C1(new_n1266), .C2(new_n1262), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(G2897), .ZN(new_n1269));
  NOR3_X1   g1069(.A1(new_n1268), .A2(new_n1269), .A3(new_n1236), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT121), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1236), .B1(new_n1271), .B2(new_n1269), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n1271), .B2(new_n1269), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1268), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT122), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1268), .A2(KEYINPUT122), .A3(new_n1273), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1270), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1250), .B1(new_n1260), .B2(new_n1278), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n1199), .A2(G378), .B1(new_n1230), .B2(new_n1255), .ZN(new_n1280));
  OAI21_X1  g1080(.A(KEYINPUT124), .B1(new_n1280), .B2(new_n1237), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT124), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1259), .A2(new_n1282), .A3(new_n1236), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1281), .A2(KEYINPUT63), .A3(new_n1268), .A4(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1285));
  AOI211_X1 g1085(.A(new_n1237), .B(new_n1285), .C1(new_n1254), .C2(new_n1258), .ZN(new_n1286));
  OR2_X1    g1086(.A1(new_n1286), .A2(KEYINPUT63), .ZN(new_n1287));
  AND2_X1   g1087(.A1(new_n1287), .A2(KEYINPUT120), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1287), .A2(KEYINPUT120), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1279), .B(new_n1284), .C1(new_n1288), .C2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT62), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1285), .A2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1281), .A2(new_n1283), .A3(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(KEYINPUT125), .B1(new_n1286), .B2(KEYINPUT62), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT125), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1295), .B(new_n1291), .C1(new_n1260), .C2(new_n1285), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1293), .A2(new_n1294), .A3(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1298));
  AOI21_X1  g1098(.A(KEYINPUT61), .B1(new_n1298), .B2(new_n1278), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1297), .A2(new_n1299), .A3(KEYINPUT126), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1247), .A2(new_n1249), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(KEYINPUT126), .B1(new_n1297), .B2(new_n1299), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1290), .B1(new_n1302), .B2(new_n1303), .ZN(G405));
  NAND2_X1  g1104(.A1(G375), .A2(new_n1230), .ZN(new_n1305));
  AND3_X1   g1105(.A1(new_n1301), .A2(new_n1254), .A3(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1301), .B1(new_n1254), .B2(new_n1305), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1285), .A2(KEYINPUT127), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  OAI22_X1  g1110(.A1(new_n1306), .A2(new_n1307), .B1(KEYINPUT127), .B2(new_n1285), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(G402));
endmodule


