//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 1 1 0 0 0 0 1 1 1 0 0 0 1 0 1 1 0 0 1 1 0 1 1 0 1 1 0 0 1 0 1 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1233, new_n1234, new_n1235, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT0), .Z(new_n206));
  INV_X1    g0006(.A(G87), .ZN(new_n207));
  INV_X1    g0007(.A(G250), .ZN(new_n208));
  INV_X1    g0008(.A(G97), .ZN(new_n209));
  INV_X1    g0009(.A(G257), .ZN(new_n210));
  OAI22_X1  g0010(.A1(new_n207), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g0011(.A(new_n211), .B1(G68), .B2(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G107), .ZN(new_n213));
  INV_X1    g0013(.A(G264), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G50), .ZN(new_n217));
  INV_X1    g0017(.A(G226), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G58), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n203), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G20), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT64), .ZN(new_n230));
  INV_X1    g0030(.A(G68), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n222), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G50), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n206), .B(new_n226), .C1(new_n230), .C2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT65), .B(G264), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G270), .ZN(new_n241));
  XOR2_X1   g0041(.A(G250), .B(G257), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n239), .B(new_n243), .Z(G358));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT66), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT67), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(new_n213), .ZN(new_n251));
  INV_X1    g0051(.A(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n249), .B(new_n254), .ZN(G351));
  XNOR2_X1  g0055(.A(KEYINPUT3), .B(G33), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G222), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G223), .A2(G1698), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n256), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  AND2_X1   g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(new_n227), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n260), .B(new_n262), .C1(G77), .C2(new_n256), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n264), .B1(G41), .B2(G45), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT68), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT68), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n267), .B(new_n264), .C1(G41), .C2(G45), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n262), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G226), .ZN(new_n270));
  INV_X1    g0070(.A(G274), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n265), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  AND3_X1   g0073(.A1(new_n263), .A2(new_n270), .A3(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G169), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n217), .A2(new_n222), .A3(new_n231), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G20), .A2(G33), .ZN(new_n279));
  AOI22_X1  g0079(.A1(new_n278), .A2(G20), .B1(G150), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT70), .ZN(new_n281));
  INV_X1    g0081(.A(G33), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n281), .B1(new_n282), .B2(G20), .ZN(new_n283));
  INV_X1    g0083(.A(G20), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n284), .A2(KEYINPUT70), .A3(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT8), .B(G58), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n280), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT69), .B1(new_n203), .B2(new_n282), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT69), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n290), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n289), .A2(new_n227), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n264), .A2(G20), .ZN(new_n293));
  INV_X1    g0093(.A(G13), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n288), .A2(new_n292), .B1(new_n217), .B2(new_n295), .ZN(new_n296));
  AND3_X1   g0096(.A1(new_n289), .A2(new_n227), .A3(new_n291), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n293), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n296), .B1(new_n217), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G179), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n274), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n277), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT9), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n299), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n274), .A2(G190), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n275), .A2(G200), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n299), .A2(new_n304), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NOR3_X1   g0110(.A1(new_n308), .A2(KEYINPUT10), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT10), .B1(new_n308), .B2(new_n310), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n303), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT3), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G33), .ZN(new_n316));
  AND3_X1   g0116(.A1(new_n282), .A2(KEYINPUT78), .A3(KEYINPUT3), .ZN(new_n317));
  AOI21_X1  g0117(.A(KEYINPUT78), .B1(new_n282), .B2(KEYINPUT3), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT7), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(new_n320), .A3(new_n284), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n282), .A2(KEYINPUT3), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT78), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(new_n315), .B2(G33), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n282), .A2(KEYINPUT78), .A3(KEYINPUT3), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n322), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(KEYINPUT7), .B1(new_n326), .B2(G20), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n321), .A2(new_n327), .A3(G68), .ZN(new_n328));
  NAND2_X1  g0128(.A1(G58), .A2(G68), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT79), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT79), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(G58), .A3(G68), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n330), .A2(new_n332), .A3(new_n232), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n333), .A2(G20), .B1(G159), .B2(new_n279), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n328), .A2(KEYINPUT16), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT16), .ZN(new_n336));
  INV_X1    g0136(.A(new_n334), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n320), .B1(new_n256), .B2(G20), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n282), .A2(KEYINPUT3), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n316), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n340), .A2(KEYINPUT7), .A3(new_n284), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n231), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n336), .B1(new_n337), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n335), .A2(new_n292), .A3(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n287), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n298), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(new_n295), .B2(new_n345), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n272), .B1(new_n269), .B2(G232), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n324), .A2(new_n325), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n351), .A2(G223), .A3(new_n257), .A4(new_n316), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT80), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(G33), .A2(G87), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n326), .A2(KEYINPUT80), .A3(G223), .A4(new_n257), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n326), .A2(G226), .A3(G1698), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n354), .A2(new_n355), .A3(new_n356), .A4(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n350), .B1(new_n358), .B2(new_n262), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n359), .A2(new_n276), .ZN(new_n360));
  AOI211_X1 g0160(.A(new_n300), .B(new_n350), .C1(new_n358), .C2(new_n262), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n348), .B(KEYINPUT18), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n358), .A2(new_n262), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n364), .A2(G179), .A3(new_n349), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(new_n276), .B2(new_n359), .ZN(new_n366));
  AOI21_X1  g0166(.A(KEYINPUT18), .B1(new_n366), .B2(new_n348), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT17), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n359), .A2(G190), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n371), .A2(new_n344), .A3(new_n347), .ZN(new_n372));
  INV_X1    g0172(.A(G200), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n359), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n370), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n348), .ZN(new_n376));
  INV_X1    g0176(.A(new_n374), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT17), .A4(new_n371), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n314), .A2(new_n369), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT73), .ZN(new_n382));
  INV_X1    g0182(.A(new_n295), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n382), .B1(new_n297), .B2(new_n383), .ZN(new_n384));
  NOR3_X1   g0184(.A1(new_n292), .A2(KEYINPUT73), .A3(new_n295), .ZN(new_n385));
  OAI211_X1 g0185(.A(G68), .B(new_n293), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT12), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n387), .B1(new_n383), .B2(G68), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n295), .A2(KEYINPUT12), .A3(new_n231), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n386), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT77), .ZN(new_n391));
  XNOR2_X1  g0191(.A(new_n390), .B(new_n391), .ZN(new_n392));
  OAI22_X1  g0192(.A1(new_n286), .A2(new_n219), .B1(new_n284), .B2(G68), .ZN(new_n393));
  INV_X1    g0193(.A(new_n279), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n394), .A2(new_n217), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n292), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  XNOR2_X1  g0196(.A(new_n396), .B(KEYINPUT11), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n272), .B1(new_n269), .B2(G238), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G33), .A2(G97), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n223), .A2(G1698), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n400), .B1(G226), .B2(G1698), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n399), .B1(new_n401), .B2(new_n340), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n262), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  XOR2_X1   g0204(.A(KEYINPUT76), .B(KEYINPUT13), .Z(new_n405));
  NOR2_X1   g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n404), .A2(KEYINPUT13), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n407), .A2(G190), .A3(new_n408), .ZN(new_n409));
  AND3_X1   g0209(.A1(new_n392), .A2(new_n397), .A3(new_n409), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n404), .A2(new_n405), .ZN(new_n411));
  OAI21_X1  g0211(.A(G200), .B1(new_n411), .B2(new_n406), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n392), .A2(new_n397), .ZN(new_n413));
  OAI21_X1  g0213(.A(G169), .B1(new_n411), .B2(new_n406), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT14), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n407), .A2(G179), .A3(new_n408), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT14), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n417), .B(G169), .C1(new_n411), .C2(new_n406), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n415), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n410), .A2(new_n412), .B1(new_n413), .B2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT75), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT74), .ZN(new_n422));
  AOI211_X1 g0222(.A(KEYINPUT71), .B(new_n272), .C1(new_n269), .C2(G244), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT71), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n266), .A2(new_n268), .ZN(new_n425));
  INV_X1    g0225(.A(new_n262), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n425), .A2(G244), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n424), .B1(new_n427), .B2(new_n273), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n423), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G238), .A2(G1698), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n256), .B(new_n430), .C1(new_n223), .C2(G1698), .ZN(new_n431));
  AND2_X1   g0231(.A1(KEYINPUT72), .A2(G107), .ZN(new_n432));
  NOR2_X1   g0232(.A1(KEYINPUT72), .A2(G107), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n431), .B(new_n262), .C1(new_n256), .C2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n373), .B1(new_n429), .B2(new_n435), .ZN(new_n436));
  OAI211_X1 g0236(.A(G77), .B(new_n293), .C1(new_n384), .C2(new_n385), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n295), .A2(new_n219), .ZN(new_n438));
  XNOR2_X1  g0238(.A(KEYINPUT15), .B(G87), .ZN(new_n439));
  OAI22_X1  g0239(.A1(new_n286), .A2(new_n439), .B1(new_n287), .B2(new_n394), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n284), .A2(new_n219), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n292), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n437), .A2(new_n438), .A3(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n422), .B1(new_n436), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n427), .A2(new_n273), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT71), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n427), .A2(new_n424), .A3(new_n273), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n446), .A2(new_n447), .A3(new_n435), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(G190), .ZN(new_n450));
  INV_X1    g0250(.A(new_n443), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n448), .A2(G200), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n451), .A2(new_n452), .A3(KEYINPUT74), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n444), .A2(new_n450), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n449), .A2(new_n300), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n448), .A2(new_n276), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n455), .A2(new_n443), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n421), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  AND3_X1   g0258(.A1(new_n454), .A2(new_n421), .A3(new_n457), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n420), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OR2_X1    g0260(.A1(new_n381), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT22), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n284), .A2(G87), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n462), .B1(new_n340), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G116), .ZN(new_n465));
  OAI21_X1  g0265(.A(KEYINPUT86), .B1(new_n465), .B2(G20), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT86), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n467), .A2(new_n284), .A3(G33), .A4(G116), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(G20), .B1(new_n432), .B2(new_n433), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT23), .ZN(new_n471));
  AND3_X1   g0271(.A1(new_n464), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT24), .ZN(new_n473));
  OR3_X1    g0273(.A1(new_n284), .A2(KEYINPUT23), .A3(G107), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n326), .A2(KEYINPUT22), .A3(new_n284), .A4(G87), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n472), .A2(new_n473), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n464), .A2(new_n471), .A3(new_n474), .A4(new_n469), .ZN(new_n477));
  NOR3_X1   g0277(.A1(new_n319), .A2(new_n462), .A3(new_n463), .ZN(new_n478));
  OAI21_X1  g0278(.A(KEYINPUT24), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n292), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n295), .A2(new_n213), .ZN(new_n482));
  XOR2_X1   g0282(.A(new_n482), .B(KEYINPUT25), .Z(new_n483));
  NOR2_X1   g0283(.A1(new_n282), .A2(G1), .ZN(new_n484));
  NOR3_X1   g0284(.A1(new_n292), .A2(new_n295), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G107), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G41), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n264), .B(G45), .C1(new_n489), .C2(KEYINPUT5), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(KEYINPUT5), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n426), .B(G264), .C1(new_n490), .C2(new_n492), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n491), .B(G274), .C1(new_n261), .C2(new_n227), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT5), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G41), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT83), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n496), .A2(new_n497), .A3(new_n264), .A4(G45), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n490), .A2(KEYINPUT83), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n494), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n208), .A2(new_n257), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n210), .A2(G1698), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n326), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G294), .ZN(new_n505));
  AND2_X1   g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n493), .B(new_n501), .C1(new_n506), .C2(new_n426), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G200), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n426), .B1(new_n504), .B2(new_n505), .ZN(new_n509));
  INV_X1    g0309(.A(new_n493), .ZN(new_n510));
  NOR3_X1   g0310(.A1(new_n509), .A2(new_n510), .A3(new_n500), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G190), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n481), .A2(new_n488), .A3(new_n508), .A4(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n507), .A2(new_n276), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n511), .A2(new_n300), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n297), .B1(new_n476), .B2(new_n479), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n514), .B(new_n515), .C1(new_n516), .C2(new_n487), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT85), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n326), .A2(new_n284), .A3(G68), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT19), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n284), .B1(new_n399), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n207), .A2(new_n209), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n523), .B1(new_n434), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n522), .B1(new_n286), .B2(new_n209), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n521), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n292), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n295), .A2(new_n439), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n485), .A2(G87), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(G238), .A2(G1698), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n532), .B1(new_n220), .B2(G1698), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n326), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n465), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n262), .ZN(new_n536));
  INV_X1    g0336(.A(G45), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n208), .B1(new_n537), .B2(G1), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n264), .A2(new_n271), .A3(G45), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n426), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n373), .B1(new_n536), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n520), .B1(new_n531), .B2(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n426), .B1(new_n534), .B2(new_n465), .ZN(new_n543));
  INV_X1    g0343(.A(new_n540), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G190), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n527), .A2(new_n292), .B1(new_n295), .B2(new_n439), .ZN(new_n547));
  OAI21_X1  g0347(.A(G200), .B1(new_n543), .B2(new_n544), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n547), .A2(new_n548), .A3(KEYINPUT85), .A4(new_n530), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n542), .A2(new_n546), .A3(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n485), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n547), .B1(new_n439), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n545), .A2(new_n300), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n552), .B(new_n553), .C1(G169), .C2(new_n545), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n252), .A2(G20), .ZN(new_n556));
  NAND2_X1  g0356(.A1(G33), .A2(G283), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n557), .B(new_n284), .C1(G33), .C2(new_n209), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n292), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT20), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n292), .A2(KEYINPUT20), .A3(new_n556), .A4(new_n558), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n561), .A2(new_n562), .B1(new_n252), .B2(new_n295), .ZN(new_n563));
  INV_X1    g0363(.A(new_n484), .ZN(new_n564));
  OAI211_X1 g0364(.A(G116), .B(new_n564), .C1(new_n384), .C2(new_n385), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n210), .A2(new_n257), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n214), .A2(G1698), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n326), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n340), .A2(G303), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n262), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n492), .A2(new_n490), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n573), .A2(new_n262), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n500), .B1(G270), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(G200), .ZN(new_n577));
  INV_X1    g0377(.A(G190), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n566), .B(new_n577), .C1(new_n578), .C2(new_n576), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT21), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n576), .A2(G169), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n580), .B1(new_n566), .B2(new_n581), .ZN(new_n582));
  AND2_X1   g0382(.A1(new_n499), .A2(new_n498), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n426), .B1(new_n490), .B2(new_n492), .ZN(new_n584));
  INV_X1    g0384(.A(G270), .ZN(new_n585));
  OAI22_X1  g0385(.A1(new_n583), .A2(new_n494), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n426), .B1(new_n569), .B2(new_n570), .ZN(new_n587));
  OAI211_X1 g0387(.A(KEYINPUT21), .B(G169), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n572), .A2(new_n575), .A3(G179), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n563), .A2(new_n565), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n579), .A2(new_n582), .A3(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n555), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT82), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT4), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n596), .A2(G1698), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n597), .A2(new_n339), .A3(new_n316), .A4(G244), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n596), .B1(new_n256), .B2(G250), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n557), .B(new_n598), .C1(new_n599), .C2(new_n257), .ZN(new_n600));
  AOI21_X1  g0400(.A(KEYINPUT4), .B1(new_n326), .B2(G244), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n595), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n596), .B1(new_n319), .B2(new_n220), .ZN(new_n603));
  OAI21_X1  g0403(.A(KEYINPUT4), .B1(new_n340), .B2(new_n208), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(G1698), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n598), .A2(new_n557), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n603), .A2(new_n605), .A3(KEYINPUT82), .A4(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n602), .A2(new_n262), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n500), .B1(G257), .B2(new_n574), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n276), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n383), .A2(G97), .ZN(new_n612));
  NOR4_X1   g0412(.A1(new_n292), .A2(new_n209), .A3(new_n295), .A4(new_n484), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT81), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT6), .ZN(new_n615));
  AND2_X1   g0415(.A1(G97), .A2(G107), .ZN(new_n616));
  NOR2_X1   g0416(.A1(G97), .A2(G107), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n213), .A2(KEYINPUT6), .A3(G97), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n284), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n394), .A2(new_n219), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n614), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n621), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n213), .A2(KEYINPUT6), .A3(G97), .ZN(new_n624));
  XNOR2_X1  g0424(.A(G97), .B(G107), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n624), .B1(new_n625), .B2(new_n615), .ZN(new_n626));
  OAI211_X1 g0426(.A(KEYINPUT81), .B(new_n623), .C1(new_n626), .C2(new_n284), .ZN(new_n627));
  AOI21_X1  g0427(.A(KEYINPUT7), .B1(new_n340), .B2(new_n284), .ZN(new_n628));
  AOI211_X1 g0428(.A(new_n320), .B(G20), .C1(new_n339), .C2(new_n316), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n434), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n622), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  AOI211_X1 g0431(.A(new_n612), .B(new_n613), .C1(new_n631), .C2(new_n292), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n608), .A2(new_n300), .A3(new_n609), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n611), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n610), .A2(G200), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n608), .A2(G190), .A3(new_n609), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(new_n632), .A3(new_n637), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n635), .A2(new_n638), .A3(KEYINPUT84), .ZN(new_n639));
  AOI21_X1  g0439(.A(KEYINPUT84), .B1(new_n635), .B2(new_n638), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n519), .B(new_n594), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n461), .A2(new_n641), .ZN(G372));
  NAND2_X1  g0442(.A1(new_n413), .A2(new_n419), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n643), .A2(new_n457), .B1(new_n410), .B2(new_n412), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n368), .B1(new_n644), .B2(new_n380), .ZN(new_n645));
  INV_X1    g0445(.A(new_n313), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n646), .A2(new_n311), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n302), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n381), .A2(new_n460), .ZN(new_n650));
  INV_X1    g0450(.A(new_n531), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n536), .A2(KEYINPUT87), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT87), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n543), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n544), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n651), .B(new_n546), .C1(new_n655), .C2(new_n373), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n517), .A2(new_n582), .A3(new_n592), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n659), .A2(new_n638), .A3(new_n513), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n658), .B1(new_n660), .B2(new_n635), .ZN(new_n661));
  OAI21_X1  g0461(.A(KEYINPUT26), .B1(new_n555), .B2(new_n635), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n655), .A2(G169), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n552), .A2(new_n553), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n650), .B1(new_n661), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n649), .A2(new_n668), .ZN(G369));
  XNOR2_X1  g0469(.A(new_n593), .B(KEYINPUT89), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n294), .A2(G20), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n264), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n673), .A2(G213), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G343), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT88), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n591), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n670), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n582), .A2(new_n592), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n680), .B1(new_n681), .B2(new_n679), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT90), .ZN(new_n683));
  XOR2_X1   g0483(.A(KEYINPUT91), .B(G330), .Z(new_n684));
  OAI21_X1  g0484(.A(new_n678), .B1(new_n516), .B2(new_n487), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n518), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n514), .A2(new_n515), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n678), .B(new_n687), .C1(new_n516), .C2(new_n487), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n683), .A2(new_n684), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n681), .A2(new_n677), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(new_n518), .ZN(new_n693));
  INV_X1    g0493(.A(new_n517), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n693), .B1(new_n694), .B2(new_n677), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n691), .A2(new_n695), .ZN(G399));
  OR3_X1    g0496(.A1(new_n434), .A2(G116), .A3(new_n524), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n204), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(G41), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n698), .A2(G1), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n233), .B2(new_n701), .ZN(new_n703));
  XOR2_X1   g0503(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n704));
  XNOR2_X1  g0504(.A(new_n703), .B(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n677), .B1(new_n661), .B2(new_n667), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT93), .ZN(new_n707));
  AOI21_X1  g0507(.A(KEYINPUT29), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n637), .A2(new_n632), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n373), .B1(new_n608), .B2(new_n609), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n513), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n712), .A2(new_n635), .A3(new_n659), .A4(new_n656), .ZN(new_n713));
  AND3_X1   g0513(.A1(new_n608), .A2(new_n300), .A3(new_n609), .ZN(new_n714));
  AOI21_X1  g0514(.A(G169), .B1(new_n608), .B2(new_n609), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n714), .A2(new_n715), .A3(new_n632), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n657), .B1(new_n716), .B2(new_n656), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n716), .A2(new_n657), .A3(new_n554), .A4(new_n550), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n713), .A2(new_n718), .A3(new_n666), .A4(new_n719), .ZN(new_n720));
  AOI22_X1  g0520(.A1(new_n706), .A2(KEYINPUT93), .B1(new_n720), .B2(new_n677), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n708), .B1(new_n721), .B2(KEYINPUT29), .ZN(new_n722));
  INV_X1    g0522(.A(new_n610), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n509), .A2(new_n510), .ZN(new_n724));
  INV_X1    g0524(.A(new_n545), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n589), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n723), .A2(KEYINPUT30), .A3(new_n724), .A4(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n655), .A2(G179), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n728), .A2(new_n507), .A3(new_n610), .A4(new_n576), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT30), .ZN(new_n730));
  INV_X1    g0530(.A(new_n726), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n608), .A2(new_n724), .A3(new_n609), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n727), .A2(new_n729), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n678), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT31), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n734), .A2(KEYINPUT31), .A3(new_n678), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n737), .B(new_n738), .C1(new_n641), .C2(new_n678), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n684), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n722), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n705), .B1(new_n742), .B2(G1), .ZN(G364));
  NAND2_X1  g0543(.A1(new_n671), .A2(G45), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n701), .A2(G1), .A3(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G13), .A2(G33), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G20), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n745), .B1(new_n682), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n256), .A2(G355), .A3(new_n204), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n249), .A2(new_n537), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n326), .A2(new_n699), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(G45), .B2(new_n233), .ZN(new_n753));
  OAI221_X1 g0553(.A(new_n750), .B1(G116), .B2(new_n204), .C1(new_n751), .C2(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n227), .B1(G20), .B2(new_n276), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n748), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n755), .ZN(new_n758));
  XNOR2_X1  g0558(.A(KEYINPUT95), .B(G159), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n284), .A2(G190), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G179), .A2(G200), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT32), .ZN(new_n765));
  OR3_X1    g0565(.A1(new_n373), .A2(KEYINPUT96), .A3(G179), .ZN(new_n766));
  OAI21_X1  g0566(.A(KEYINPUT96), .B1(new_n373), .B2(G179), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n284), .A2(new_n578), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n340), .B1(new_n770), .B2(G87), .ZN(new_n771));
  OR2_X1    g0571(.A1(new_n771), .A2(KEYINPUT97), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n766), .A2(new_n767), .A3(new_n761), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G107), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n771), .A2(KEYINPUT97), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n772), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT98), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n762), .A2(G190), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G20), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n209), .ZN(new_n782));
  NAND2_X1  g0582(.A1(G20), .A2(G179), .ZN(new_n783));
  XOR2_X1   g0583(.A(new_n783), .B(KEYINPUT94), .Z(new_n784));
  NOR2_X1   g0584(.A1(new_n578), .A2(G200), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n782), .B1(new_n787), .B2(G58), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n784), .A2(new_n578), .A3(G200), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G68), .ZN(new_n791));
  AND4_X1   g0591(.A1(new_n765), .A2(new_n778), .A3(new_n788), .A4(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n784), .A2(G190), .A3(G200), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n784), .A2(new_n578), .A3(new_n373), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n792), .B1(new_n217), .B2(new_n793), .C1(new_n219), .C2(new_n794), .ZN(new_n795));
  XOR2_X1   g0595(.A(KEYINPUT33), .B(G317), .Z(new_n796));
  INV_X1    g0596(.A(G322), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n789), .A2(new_n796), .B1(new_n786), .B2(new_n797), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n798), .B(KEYINPUT99), .Z(new_n799));
  INV_X1    g0599(.A(new_n793), .ZN(new_n800));
  INV_X1    g0600(.A(new_n763), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n800), .A2(G326), .B1(G329), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G303), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n802), .B(new_n340), .C1(new_n803), .C2(new_n769), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n799), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n780), .A2(G294), .ZN(new_n806));
  INV_X1    g0606(.A(new_n794), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G311), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n774), .A2(G283), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n805), .A2(new_n806), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  AND2_X1   g0610(.A1(new_n795), .A2(new_n810), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n749), .B(new_n757), .C1(new_n758), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n683), .A2(new_n684), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(new_n745), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n683), .A2(new_n684), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n812), .B1(new_n814), .B2(new_n815), .ZN(G396));
  NAND2_X1  g0616(.A1(new_n678), .A2(new_n443), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n454), .A2(new_n457), .A3(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n677), .A2(new_n451), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n819), .A2(KEYINPUT102), .A3(new_n456), .A4(new_n455), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT102), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n455), .A2(new_n456), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n821), .B1(new_n817), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n818), .A2(new_n820), .A3(new_n823), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n706), .B(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(new_n740), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n745), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n793), .A2(new_n803), .B1(new_n213), .B2(new_n769), .ZN(new_n828));
  INV_X1    g0628(.A(G311), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n340), .B1(new_n763), .B2(new_n829), .C1(new_n773), .C2(new_n207), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n794), .A2(new_n252), .ZN(new_n831));
  NOR4_X1   g0631(.A1(new_n828), .A2(new_n830), .A3(new_n831), .A4(new_n782), .ZN(new_n832));
  INV_X1    g0632(.A(G283), .ZN(new_n833));
  INV_X1    g0633(.A(G294), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n832), .B1(new_n833), .B2(new_n789), .C1(new_n834), .C2(new_n786), .ZN(new_n835));
  INV_X1    g0635(.A(G150), .ZN(new_n836));
  INV_X1    g0636(.A(G143), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n789), .A2(new_n836), .B1(new_n786), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(G137), .B2(new_n800), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n794), .B2(new_n760), .ZN(new_n840));
  XOR2_X1   g0640(.A(new_n840), .B(KEYINPUT34), .Z(new_n841));
  AOI22_X1  g0641(.A1(new_n770), .A2(G50), .B1(G132), .B2(new_n801), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n774), .A2(G68), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n842), .A2(new_n326), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(G58), .B2(new_n780), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT101), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n835), .B1(new_n841), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n755), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n755), .A2(new_n746), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n745), .B1(new_n219), .B2(new_n849), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(KEYINPUT100), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n848), .B(new_n851), .C1(new_n747), .C2(new_n824), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n827), .A2(new_n852), .ZN(G384));
  INV_X1    g0653(.A(new_n626), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n252), .B1(new_n854), .B2(KEYINPUT35), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n855), .B(new_n230), .C1(KEYINPUT35), .C2(new_n854), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT36), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n234), .A2(G77), .A3(new_n332), .A4(new_n330), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(KEYINPUT103), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(G50), .B2(new_n231), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n860), .A2(G1), .A3(new_n294), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT104), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT40), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n335), .A2(new_n292), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT16), .B1(new_n328), .B2(new_n334), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n347), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n675), .B(new_n867), .C1(new_n368), .C2(new_n379), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n376), .A2(new_n377), .A3(new_n371), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n366), .A2(new_n675), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n869), .B(new_n870), .C1(new_n871), .C2(new_n376), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n372), .A2(new_n374), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n360), .A2(new_n361), .ZN(new_n874));
  INV_X1    g0674(.A(new_n675), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n873), .B1(new_n876), .B2(new_n867), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n872), .B1(new_n877), .B2(new_n870), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n868), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT38), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n868), .A2(new_n878), .A3(KEYINPUT38), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n677), .B1(new_n392), .B2(new_n397), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n885), .A2(new_n419), .ZN(new_n886));
  INV_X1    g0686(.A(new_n885), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n886), .B1(new_n420), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n739), .A2(new_n889), .A3(new_n824), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n864), .B1(new_n884), .B2(new_n890), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n868), .A2(new_n878), .A3(KEYINPUT38), .ZN(new_n892));
  XOR2_X1   g0692(.A(KEYINPUT106), .B(KEYINPUT38), .Z(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n348), .B(new_n675), .C1(new_n368), .C2(new_n379), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n376), .B1(new_n874), .B2(new_n875), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT37), .B1(new_n896), .B2(new_n873), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n872), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n894), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(KEYINPUT40), .B1(new_n892), .B2(new_n899), .ZN(new_n900));
  OR2_X1    g0700(.A1(new_n900), .A2(new_n890), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n891), .A2(new_n901), .ZN(new_n902));
  XOR2_X1   g0702(.A(new_n902), .B(KEYINPUT107), .Z(new_n903));
  NAND2_X1  g0703(.A1(new_n650), .A2(new_n739), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n903), .B(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n684), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n677), .B(new_n824), .C1(new_n661), .C2(new_n667), .ZN(new_n907));
  OR2_X1    g0707(.A1(new_n457), .A2(new_n678), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT105), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n907), .A2(KEYINPUT105), .A3(new_n908), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n888), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n883), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT39), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n892), .B2(new_n899), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n881), .A2(KEYINPUT39), .A3(new_n882), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n413), .A2(new_n419), .A3(new_n677), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n916), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n368), .A2(new_n875), .ZN(new_n921));
  AND3_X1   g0721(.A1(new_n914), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n635), .A2(new_n656), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n719), .B(new_n666), .C1(new_n660), .C2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n677), .B1(new_n924), .B2(new_n717), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n517), .A2(new_n582), .A3(new_n592), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n635), .B1(new_n926), .B2(new_n711), .ZN(new_n927));
  INV_X1    g0727(.A(new_n658), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n716), .A2(new_n554), .A3(new_n550), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n665), .B1(new_n930), .B2(KEYINPUT26), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n678), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n925), .B(KEYINPUT29), .C1(new_n932), .C2(new_n707), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT29), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n932), .B2(KEYINPUT93), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n461), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n936), .A2(new_n648), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n922), .B(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n906), .B(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n671), .A2(new_n264), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n863), .B1(new_n939), .B2(new_n940), .ZN(G367));
  INV_X1    g0741(.A(G137), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n763), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n780), .A2(G68), .ZN(new_n944));
  OAI221_X1 g0744(.A(new_n944), .B1(new_n786), .B2(new_n836), .C1(new_n837), .C2(new_n793), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT113), .Z(new_n946));
  NAND2_X1  g0746(.A1(new_n807), .A2(G50), .ZN(new_n947));
  AOI22_X1  g0747(.A1(G58), .A2(new_n770), .B1(new_n774), .B2(G77), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n946), .A2(new_n256), .A3(new_n947), .A4(new_n948), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n943), .B(new_n949), .C1(new_n790), .C2(new_n759), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n780), .A2(new_n434), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n793), .A2(new_n829), .B1(new_n786), .B2(new_n803), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n952), .B(KEYINPUT112), .Z(new_n953));
  NAND2_X1  g0753(.A1(new_n774), .A2(G97), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n794), .B2(new_n833), .ZN(new_n955));
  AOI211_X1 g0755(.A(new_n326), .B(new_n955), .C1(G294), .C2(new_n790), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n770), .A2(KEYINPUT46), .A3(G116), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT46), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n769), .B2(new_n252), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n953), .A2(new_n956), .A3(new_n957), .A4(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(G317), .B2(new_n801), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n950), .B1(new_n951), .B2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT47), .Z(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n755), .ZN(new_n964));
  INV_X1    g0764(.A(new_n745), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n666), .A2(new_n656), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n678), .A2(new_n531), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT108), .ZN(new_n968));
  MUX2_X1   g0768(.A(new_n966), .B(new_n666), .S(new_n968), .Z(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT109), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n748), .ZN(new_n971));
  INV_X1    g0771(.A(new_n752), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n756), .B1(new_n204), .B2(new_n439), .C1(new_n243), .C2(new_n972), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n964), .A2(new_n965), .A3(new_n971), .A4(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n744), .A2(G1), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n709), .A2(new_n710), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n716), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n678), .A2(new_n633), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n716), .A2(new_n678), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n695), .A2(new_n981), .ZN(new_n982));
  XOR2_X1   g0782(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n983));
  XNOR2_X1  g0783(.A(new_n982), .B(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n695), .A2(new_n981), .ZN(new_n985));
  NOR2_X1   g0785(.A1(KEYINPUT111), .A2(KEYINPUT44), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n985), .B(new_n986), .Z(new_n987));
  AND2_X1   g0787(.A1(KEYINPUT111), .A2(KEYINPUT44), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n984), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(new_n691), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n693), .B1(new_n689), .B2(new_n692), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n683), .A2(new_n684), .A3(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n992), .B1(new_n683), .B2(new_n684), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n996), .A2(new_n741), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n990), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n742), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n700), .B(KEYINPUT41), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n975), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT43), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n970), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n693), .A2(new_n977), .A3(new_n978), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT42), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n977), .A2(new_n694), .A3(new_n978), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n678), .B1(new_n1006), .B2(new_n635), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1003), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n691), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1009), .A2(new_n1010), .A3(new_n981), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n981), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1003), .B(new_n1008), .C1(new_n691), .C2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n970), .A2(new_n1002), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n974), .B1(new_n1001), .B2(new_n1016), .ZN(G387));
  INV_X1    g0817(.A(G317), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n789), .A2(new_n829), .B1(new_n786), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(G322), .B2(new_n800), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n803), .B2(new_n794), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT48), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1022), .B1(new_n833), .B2(new_n781), .C1(new_n834), .C2(new_n769), .ZN(new_n1023));
  XOR2_X1   g0823(.A(KEYINPUT115), .B(KEYINPUT49), .Z(new_n1024));
  XNOR2_X1  g0824(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n773), .A2(new_n252), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n326), .B(new_n1026), .C1(G326), .C2(new_n801), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n787), .A2(G50), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n801), .A2(G150), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n770), .A2(G77), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(G159), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n954), .B1(new_n793), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n326), .B1(new_n789), .B2(new_n287), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n781), .A2(new_n439), .ZN(new_n1036));
  NOR4_X1   g0836(.A1(new_n1032), .A2(new_n1034), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n231), .B2(new_n794), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n758), .B1(new_n1028), .B2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n697), .A2(new_n204), .A3(new_n256), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n239), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n752), .B1(new_n1041), .B2(new_n537), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n345), .A2(new_n217), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n698), .B1(KEYINPUT50), .B2(new_n1043), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n1043), .A2(KEYINPUT50), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n231), .A2(new_n219), .ZN(new_n1046));
  NOR4_X1   g0846(.A1(new_n1044), .A2(new_n1045), .A3(G45), .A4(new_n1046), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1040), .B1(G107), .B2(new_n204), .C1(new_n1042), .C2(new_n1047), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT114), .Z(new_n1049));
  AOI211_X1 g0849(.A(new_n745), .B(new_n1039), .C1(new_n756), .C2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT116), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n689), .A2(new_n748), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n996), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n1051), .A2(new_n1052), .B1(new_n975), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n700), .B1(new_n1053), .B2(new_n742), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1054), .B1(new_n997), .B2(new_n1055), .ZN(G393));
  NOR2_X1   g0856(.A1(new_n990), .A2(new_n997), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1057), .A2(new_n701), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n998), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n990), .A2(new_n975), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n793), .A2(new_n1018), .B1(new_n786), .B2(new_n829), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT52), .Z(new_n1062));
  AOI211_X1 g0862(.A(new_n256), .B(new_n1062), .C1(G294), .C2(new_n807), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n833), .B2(new_n769), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n781), .A2(new_n252), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n763), .A2(new_n797), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n775), .B1(new_n789), .B2(new_n803), .ZN(new_n1067));
  NOR4_X1   g0867(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n789), .A2(new_n217), .B1(new_n207), .B2(new_n773), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n794), .A2(new_n287), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n326), .B1(new_n763), .B2(new_n837), .C1(new_n781), .C2(new_n219), .ZN(new_n1071));
  OR3_X1    g0871(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n793), .A2(new_n836), .B1(new_n786), .B2(new_n1033), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT51), .Z(new_n1074));
  AOI211_X1 g0874(.A(new_n1072), .B(new_n1074), .C1(G68), .C2(new_n770), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n755), .B1(new_n1068), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1012), .A2(new_n748), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n756), .B1(new_n209), .B2(new_n204), .C1(new_n254), .C2(new_n972), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1076), .A2(new_n965), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1059), .A2(new_n1060), .A3(new_n1079), .ZN(G390));
  NAND2_X1  g0880(.A1(new_n916), .A2(new_n917), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n913), .B2(new_n919), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n677), .B(new_n824), .C1(new_n924), .C2(new_n717), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n908), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n889), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n895), .A2(new_n898), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n893), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n919), .B1(new_n1087), .B2(new_n882), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1085), .A2(new_n1088), .A3(KEYINPUT117), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT117), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n918), .B1(new_n892), .B2(new_n899), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n888), .B1(new_n1083), .B2(new_n908), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1090), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1089), .A2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n739), .A2(new_n889), .A3(new_n684), .A4(new_n824), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n1082), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n739), .A2(new_n889), .A3(G330), .A4(new_n824), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(new_n1082), .B2(new_n1094), .ZN(new_n1098));
  AND3_X1   g0898(.A1(new_n650), .A2(new_n739), .A3(G330), .ZN(new_n1099));
  NOR3_X1   g0899(.A1(new_n936), .A2(new_n648), .A3(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n739), .A2(G330), .A3(new_n824), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n888), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1084), .ZN(new_n1103));
  AND3_X1   g0903(.A1(new_n1102), .A2(new_n1103), .A3(new_n1095), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n739), .A2(new_n684), .A3(new_n824), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n888), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1106), .A2(new_n1097), .B1(new_n911), .B2(new_n912), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1100), .B1(new_n1104), .B2(new_n1107), .ZN(new_n1108));
  NOR3_X1   g0908(.A1(new_n1096), .A2(new_n1098), .A3(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1109), .A2(new_n701), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n650), .A2(new_n739), .A3(G330), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n649), .B(new_n1112), .C1(new_n722), .C2(new_n461), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n1105), .A2(new_n888), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1097), .ZN(new_n1115));
  AOI21_X1  g0915(.A(KEYINPUT105), .B1(new_n907), .B2(new_n908), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n907), .A2(KEYINPUT105), .A3(new_n908), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n1114), .A2(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1102), .A2(new_n1103), .A3(new_n1095), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1113), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1110), .B1(new_n1111), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1111), .A2(new_n975), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n340), .B1(new_n787), .B2(G132), .ZN(new_n1123));
  AND3_X1   g0923(.A1(new_n770), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1124));
  AOI21_X1  g0924(.A(KEYINPUT53), .B1(new_n770), .B2(G150), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n1123), .B1(new_n942), .B2(new_n789), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n800), .A2(G128), .B1(G125), .B2(new_n801), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n1033), .B2(new_n781), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT54), .B(G143), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n794), .A2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n773), .A2(new_n217), .ZN(new_n1131));
  NOR4_X1   g0931(.A1(new_n1126), .A2(new_n1128), .A3(new_n1130), .A4(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n256), .B1(new_n800), .B2(G283), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n807), .A2(G97), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n770), .A2(G87), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .A4(new_n843), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n434), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n789), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n763), .A2(new_n834), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n786), .A2(new_n252), .B1(new_n781), .B2(new_n219), .ZN(new_n1140));
  NOR4_X1   g0940(.A1(new_n1136), .A2(new_n1138), .A3(new_n1139), .A4(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n755), .B1(new_n1132), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n849), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1142), .B(new_n965), .C1(new_n345), .C2(new_n1143), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1081), .A2(new_n746), .B1(KEYINPUT118), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(KEYINPUT118), .B2(new_n1144), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1121), .A2(new_n1122), .A3(new_n1146), .ZN(G378));
  INV_X1    g0947(.A(KEYINPUT121), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1148), .B1(new_n1109), .B2(new_n1113), .ZN(new_n1149));
  XOR2_X1   g0949(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1150));
  XNOR2_X1  g0950(.A(new_n314), .B(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n299), .A2(new_n675), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1151), .B(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(G330), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1153), .B1(new_n902), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1153), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1156), .A2(new_n891), .A3(new_n901), .A4(G330), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n1155), .A2(new_n922), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n922), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  AND2_X1   g0960(.A1(new_n1089), .A2(new_n1093), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n889), .B1(new_n1117), .B2(new_n1116), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n1162), .A2(new_n918), .B1(new_n916), .B2(new_n917), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1115), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1082), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1164), .A2(new_n1120), .A3(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1166), .A2(KEYINPUT121), .A3(new_n1100), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1149), .A2(new_n1160), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT57), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n701), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  AND3_X1   g0970(.A1(new_n1166), .A2(KEYINPUT121), .A3(new_n1100), .ZN(new_n1171));
  AOI21_X1  g0971(.A(KEYINPUT121), .B1(new_n1166), .B2(new_n1100), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT122), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1173), .A2(new_n1174), .A3(KEYINPUT57), .A4(new_n1160), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1149), .A2(KEYINPUT57), .A3(new_n1160), .A4(new_n1167), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(KEYINPUT122), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1170), .A2(new_n1175), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(G124), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n282), .B1(new_n763), .B2(new_n1179), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n790), .A2(G132), .B1(new_n800), .B2(G125), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n787), .A2(G128), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n807), .A2(G137), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1184), .B1(new_n836), .B2(new_n781), .C1(new_n769), .C2(new_n1129), .ZN(new_n1185));
  AOI211_X1 g0985(.A(G41), .B(new_n1180), .C1(new_n1185), .C2(KEYINPUT59), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1186), .B1(KEYINPUT59), .B2(new_n1185), .C1(new_n773), .C2(new_n760), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n774), .A2(G58), .ZN(new_n1188));
  AOI21_X1  g0988(.A(G41), .B1(new_n801), .B2(G283), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1188), .B(new_n1189), .C1(new_n439), .C2(new_n794), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n326), .B(new_n1190), .C1(G97), .C2(new_n790), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n787), .A2(G107), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n944), .B1(new_n793), .B2(new_n252), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n1193), .B(KEYINPUT119), .Z(new_n1194));
  NAND4_X1  g0994(.A1(new_n1191), .A2(new_n1031), .A3(new_n1192), .A4(new_n1194), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT58), .ZN(new_n1196));
  AOI21_X1  g0996(.A(G41), .B1(new_n326), .B2(G33), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1187), .B(new_n1196), .C1(G50), .C2(new_n1197), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT120), .Z(new_n1199));
  NOR2_X1   g0999(.A1(new_n1199), .A2(new_n758), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1143), .A2(G50), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1153), .A2(new_n747), .ZN(new_n1202));
  NOR4_X1   g1002(.A1(new_n1200), .A2(new_n745), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n1160), .B2(new_n975), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1178), .A2(new_n1204), .ZN(G375));
  NOR2_X1   g1005(.A1(new_n1104), .A2(new_n1107), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(new_n1113), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1207), .A2(new_n1000), .A3(new_n1108), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n889), .A2(new_n747), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1143), .A2(G68), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n340), .B1(new_n793), .B2(new_n834), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n786), .A2(new_n833), .B1(new_n773), .B2(new_n219), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n252), .B2(new_n789), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1036), .B(new_n1214), .C1(G97), .C2(new_n770), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n1215), .B1(new_n803), .B2(new_n763), .C1(new_n1137), .C2(new_n794), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1188), .B1(new_n786), .B2(new_n942), .C1(new_n789), .C2(new_n1129), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n319), .B(new_n1217), .C1(G132), .C2(new_n800), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n801), .A2(G128), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n770), .A2(G159), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n807), .A2(G150), .B1(G50), .B2(new_n780), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n758), .B1(new_n1216), .B2(new_n1222), .ZN(new_n1223));
  NOR4_X1   g1023(.A1(new_n1209), .A2(new_n745), .A3(new_n1210), .A4(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1206), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1224), .B1(new_n1225), .B2(new_n975), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1208), .A2(new_n1226), .ZN(G381));
  NOR2_X1   g1027(.A1(G375), .A2(G378), .ZN(new_n1228));
  INV_X1    g1028(.A(G381), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(G387), .A2(G390), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .A4(new_n1231), .ZN(G407));
  INV_X1    g1032(.A(G213), .ZN(new_n1233));
  INV_X1    g1033(.A(G343), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1233), .B1(new_n1228), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(G407), .ZN(G409));
  NAND3_X1  g1036(.A1(new_n1178), .A2(G378), .A3(new_n1204), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT123), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1178), .A2(KEYINPUT123), .A3(G378), .A4(new_n1204), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1173), .A2(new_n1000), .A3(new_n1160), .ZN(new_n1242));
  AOI21_X1  g1042(.A(G378), .B1(new_n1204), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1241), .A2(new_n1244), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1233), .A2(G343), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT60), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n701), .B1(new_n1207), .B2(new_n1248), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1249), .B(new_n1108), .C1(new_n1248), .C2(new_n1207), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n1226), .ZN(new_n1251));
  INV_X1    g1051(.A(G384), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1250), .A2(G384), .A3(new_n1226), .ZN(new_n1254));
  AND2_X1   g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1245), .A2(new_n1247), .A3(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT124), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT125), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1255), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1260));
  OAI21_X1  g1060(.A(KEYINPUT125), .B1(new_n1260), .B2(KEYINPUT124), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1259), .A2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1260), .A2(KEYINPUT124), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1246), .A2(G2897), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1262), .A2(new_n1265), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1259), .A2(new_n1264), .A3(new_n1261), .A4(new_n1263), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1268), .B1(new_n1245), .B2(new_n1247), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT63), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1256), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT61), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(G393), .B(G396), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  AND2_X1   g1074(.A1(G387), .A2(G390), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1274), .B1(new_n1230), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1230), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(G387), .A2(G390), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1277), .A2(new_n1273), .A3(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1276), .A2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1243), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1281));
  NOR3_X1   g1081(.A1(new_n1281), .A2(new_n1246), .A3(new_n1260), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1280), .B1(new_n1282), .B2(KEYINPUT63), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1271), .A2(new_n1272), .A3(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT126), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1277), .A2(new_n1273), .A3(new_n1278), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1273), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1285), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1276), .A2(KEYINPUT126), .A3(new_n1279), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1267), .B(new_n1266), .C1(new_n1281), .C2(new_n1246), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT62), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1291), .B1(new_n1282), .B2(new_n1292), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1245), .A2(new_n1292), .A3(new_n1247), .A4(new_n1255), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1272), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1290), .B1(new_n1293), .B2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1284), .A2(new_n1296), .ZN(G405));
  INV_X1    g1097(.A(KEYINPUT127), .ZN(new_n1298));
  AND3_X1   g1098(.A1(new_n1288), .A2(new_n1298), .A3(new_n1289), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1298), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(G378), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(G375), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1241), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1255), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1241), .A2(new_n1260), .A3(new_n1303), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  MUX2_X1   g1107(.A(new_n1301), .B(new_n1299), .S(new_n1307), .Z(G402));
endmodule


