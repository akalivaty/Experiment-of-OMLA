//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 1 0 0 1 0 0 1 1 1 0 0 0 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n548, new_n550, new_n551,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n568,
    new_n569, new_n570, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1160,
    new_n1161, new_n1162, new_n1164;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT65), .Z(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT66), .Z(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n454), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2106), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT67), .Z(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n460), .B1(new_n461), .B2(new_n455), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT68), .Z(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  XNOR2_X1  g042(.A(new_n467), .B(KEYINPUT69), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n464), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n465), .A2(G137), .ZN(new_n470));
  NAND2_X1  g045(.A1(G101), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(G2105), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n469), .A2(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n465), .A2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  NOR2_X1   g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  OAI21_X1  g052(.A(G2104), .B1(new_n464), .B2(G112), .ZN(new_n478));
  INV_X1    g053(.A(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(KEYINPUT3), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g058(.A(KEYINPUT70), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n465), .A2(new_n485), .A3(new_n464), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G136), .ZN(new_n488));
  OAI221_X1 g063(.A(new_n476), .B1(new_n477), .B2(new_n478), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  NAND3_X1  g065(.A1(new_n480), .A2(new_n482), .A3(G126), .ZN(new_n491));
  NAND2_X1  g066(.A1(G114), .A2(G2104), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n464), .A2(G102), .A3(G2104), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n480), .A2(new_n482), .A3(G138), .A4(new_n464), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n465), .A2(KEYINPUT4), .A3(G138), .A4(new_n464), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n494), .A2(new_n495), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(G62), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(KEYINPUT72), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT72), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT5), .A3(G543), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n502), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  AND2_X1   g083(.A1(G75), .A2(G543), .ZN(new_n509));
  OAI21_X1  g084(.A(G651), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n512), .B2(G651), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(KEYINPUT71), .A3(KEYINPUT6), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n513), .A2(new_n515), .B1(new_n512), .B2(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n505), .A2(new_n507), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n516), .A2(G88), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n516), .A2(G50), .A3(G543), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n510), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(G166));
  NAND3_X1  g096(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n513), .A2(new_n515), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n512), .A2(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(G543), .A3(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G51), .ZN(new_n526));
  INV_X1    g101(.A(G89), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n517), .A2(new_n523), .A3(new_n524), .ZN(new_n528));
  OAI221_X1 g103(.A(new_n522), .B1(new_n525), .B2(new_n526), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT73), .ZN(new_n531));
  XOR2_X1   g106(.A(new_n531), .B(KEYINPUT7), .Z(new_n532));
  NOR2_X1   g107(.A1(new_n529), .A2(new_n532), .ZN(G168));
  AOI22_X1  g108(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(new_n514), .ZN(new_n535));
  INV_X1    g110(.A(new_n528), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G90), .ZN(new_n537));
  INV_X1    g112(.A(new_n525), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G52), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n535), .A2(new_n537), .A3(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  AOI22_X1  g116(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(new_n514), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n536), .A2(G81), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n538), .A2(G43), .ZN(new_n545));
  AND3_X1   g120(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(new_n551), .ZN(G188));
  INV_X1    g127(.A(KEYINPUT74), .ZN(new_n553));
  AND3_X1   g128(.A1(new_n516), .A2(new_n553), .A3(new_n517), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n553), .B1(new_n516), .B2(new_n517), .ZN(new_n555));
  OAI21_X1  g130(.A(G91), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(G53), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT9), .B1(new_n525), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  NAND4_X1  g134(.A1(new_n516), .A2(new_n559), .A3(G53), .A4(G543), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  AND2_X1   g136(.A1(new_n517), .A2(G65), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT75), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n556), .A2(new_n561), .A3(new_n565), .ZN(G299));
  INV_X1    g141(.A(G168), .ZN(G286));
  NAND2_X1  g142(.A1(new_n520), .A2(KEYINPUT76), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT76), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n510), .A2(new_n518), .A3(new_n519), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(G303));
  NAND2_X1  g146(.A1(new_n528), .A2(KEYINPUT74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n516), .A2(new_n553), .A3(new_n517), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G87), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n538), .A2(G49), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(G288));
  NAND2_X1  g153(.A1(new_n538), .A2(G48), .ZN(new_n579));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n580), .B1(new_n505), .B2(new_n507), .ZN(new_n581));
  AND2_X1   g156(.A1(G73), .A2(G543), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(KEYINPUT77), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT77), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n585), .B(G651), .C1(new_n581), .C2(new_n582), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n579), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(G86), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n588), .B1(new_n572), .B2(new_n573), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n592), .A2(new_n514), .ZN(new_n593));
  XNOR2_X1  g168(.A(KEYINPUT78), .B(G85), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n536), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n538), .A2(G47), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n593), .A2(new_n595), .A3(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n574), .A2(G92), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(KEYINPUT10), .ZN(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(new_n517), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(G651), .A2(new_n604), .B1(new_n538), .B2(G54), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n574), .A2(new_n606), .A3(G92), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n600), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n598), .B1(new_n609), .B2(G868), .ZN(G284));
  OAI21_X1  g185(.A(new_n598), .B1(new_n609), .B2(G868), .ZN(G321));
  INV_X1    g186(.A(KEYINPUT79), .ZN(new_n612));
  INV_X1    g187(.A(G868), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(G168), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g189(.A1(G168), .A2(new_n613), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n615), .B1(new_n613), .B2(G299), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n614), .B1(new_n616), .B2(new_n612), .ZN(G297));
  OAI21_X1  g192(.A(new_n614), .B1(new_n616), .B2(new_n612), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n609), .B1(new_n619), .B2(G860), .ZN(G148));
  NAND3_X1  g195(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(new_n613), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n608), .A2(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(new_n613), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g200(.A(new_n487), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n626), .A2(G135), .B1(G123), .B2(new_n475), .ZN(new_n627));
  NOR2_X1   g202(.A1(G99), .A2(G2105), .ZN(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(new_n464), .B2(G111), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT80), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2096), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT12), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT13), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2100), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n632), .A2(new_n636), .ZN(G156));
  XNOR2_X1  g212(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(KEYINPUT15), .B(G2435), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2438), .ZN(new_n641));
  XOR2_X1   g216(.A(G2427), .B(G2430), .Z(new_n642));
  OAI21_X1  g217(.A(KEYINPUT14), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT82), .Z(new_n644));
  NAND2_X1  g219(.A1(new_n641), .A2(new_n642), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT83), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2451), .B(G2454), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2443), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2446), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n647), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n651), .A2(new_n653), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n639), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n658), .A2(new_n638), .A3(new_n654), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n657), .A2(new_n659), .A3(G14), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(G401));
  XOR2_X1   g236(.A(G2072), .B(G2078), .Z(new_n662));
  XOR2_X1   g237(.A(G2067), .B(G2678), .Z(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n662), .B1(new_n666), .B2(KEYINPUT18), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G2096), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2100), .ZN(new_n669));
  AND2_X1   g244(.A1(new_n666), .A2(KEYINPUT17), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n664), .A2(new_n665), .ZN(new_n671));
  AOI21_X1  g246(.A(KEYINPUT18), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n669), .B(new_n672), .Z(G227));
  XNOR2_X1  g248(.A(KEYINPUT22), .B(G1981), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1971), .B(G1976), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT84), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT19), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1956), .B(G2474), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1961), .B(G1966), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n680), .B(new_n681), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n680), .A2(new_n681), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n679), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT85), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n686), .A2(KEYINPUT20), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(KEYINPUT20), .ZN(new_n688));
  OAI221_X1 g263(.A(new_n682), .B1(new_n679), .B2(new_n683), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(G1986), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n691), .A2(new_n693), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n675), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n696), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n698), .A2(new_n674), .A3(new_n694), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n697), .A2(new_n699), .ZN(G229));
  INV_X1    g275(.A(KEYINPUT88), .ZN(new_n701));
  NAND2_X1  g276(.A1(G288), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g277(.A1(new_n575), .A2(KEYINPUT88), .A3(new_n576), .A4(new_n577), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G16), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G16), .B2(G23), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT33), .B(G1976), .Z(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G22), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G166), .B2(new_n710), .ZN(new_n712));
  INV_X1    g287(.A(G1971), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n706), .A2(new_n708), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n710), .A2(G6), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(new_n590), .B2(new_n710), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT32), .B(G1981), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND4_X1  g294(.A1(new_n709), .A2(new_n714), .A3(new_n715), .A4(new_n719), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n720), .A2(KEYINPUT34), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n720), .A2(KEYINPUT34), .B1(KEYINPUT89), .B2(KEYINPUT36), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n710), .A2(G24), .ZN(new_n723));
  INV_X1    g298(.A(G290), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(new_n710), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(G1986), .Z(new_n726));
  AOI22_X1  g301(.A1(new_n626), .A2(G131), .B1(G119), .B2(new_n475), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT86), .ZN(new_n728));
  OR3_X1    g303(.A1(new_n728), .A2(G95), .A3(G2105), .ZN(new_n729));
  INV_X1    g304(.A(G107), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n479), .B1(new_n730), .B2(G2105), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n728), .B1(G95), .B2(G2105), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n729), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT87), .Z(new_n734));
  NAND2_X1  g309(.A1(new_n727), .A2(new_n734), .ZN(new_n735));
  MUX2_X1   g310(.A(G25), .B(new_n735), .S(G29), .Z(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT35), .B(G1991), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n736), .B(new_n738), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n721), .A2(new_n722), .A3(new_n726), .A4(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(KEYINPUT89), .A2(KEYINPUT36), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(G16), .A2(G19), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n546), .B2(G16), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT90), .B(G1341), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(G5), .A2(G16), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G171), .B2(G16), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT31), .ZN(new_n749));
  OAI22_X1  g324(.A1(new_n748), .A2(G1961), .B1(new_n749), .B2(G11), .ZN(new_n750));
  AOI211_X1 g325(.A(new_n746), .B(new_n750), .C1(new_n749), .C2(G11), .ZN(new_n751));
  OR2_X1    g326(.A1(KEYINPUT24), .A2(G34), .ZN(new_n752));
  INV_X1    g327(.A(G29), .ZN(new_n753));
  NAND2_X1  g328(.A1(KEYINPUT24), .A2(G34), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G160), .B2(new_n753), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT94), .B(G2084), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n753), .A2(G27), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G164), .B2(new_n753), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G2078), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT98), .B(G28), .Z(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT30), .ZN(new_n763));
  AOI211_X1 g338(.A(new_n758), .B(new_n761), .C1(new_n753), .C2(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(G29), .A2(G32), .ZN(new_n765));
  NAND3_X1  g340(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT26), .Z(new_n767));
  NAND3_X1  g342(.A1(new_n464), .A2(G105), .A3(G2104), .ZN(new_n768));
  INV_X1    g343(.A(G129), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n767), .B(new_n768), .C1(new_n769), .C2(new_n474), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n626), .A2(G141), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n771), .A2(KEYINPUT95), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(KEYINPUT95), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n770), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n765), .B1(new_n774), .B2(G29), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT27), .B(G1996), .Z(new_n776));
  AOI22_X1  g351(.A1(new_n775), .A2(new_n776), .B1(new_n748), .B2(G1961), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n751), .A2(new_n764), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n753), .A2(G35), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G162), .B2(new_n753), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT29), .B(G2090), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n630), .A2(new_n753), .ZN(new_n783));
  NOR3_X1   g358(.A1(new_n778), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n710), .A2(G20), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT100), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT23), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G299), .B2(G16), .ZN(new_n788));
  INV_X1    g363(.A(G1956), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n744), .B2(new_n745), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n753), .A2(G26), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n626), .A2(G140), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n475), .A2(G128), .ZN(new_n794));
  OR2_X1    g369(.A1(G104), .A2(G2105), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n795), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n793), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n792), .B1(new_n798), .B2(new_n753), .ZN(new_n799));
  MUX2_X1   g374(.A(new_n792), .B(new_n799), .S(KEYINPUT28), .Z(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(G2067), .ZN(new_n801));
  NAND2_X1  g376(.A1(G168), .A2(G16), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G16), .B2(G21), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT97), .B(G1966), .Z(new_n804));
  OAI21_X1  g379(.A(new_n801), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n803), .A2(new_n804), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT99), .Z(new_n807));
  NAND2_X1  g382(.A1(new_n710), .A2(G4), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(new_n609), .B2(new_n710), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(G1348), .ZN(new_n810));
  NOR3_X1   g385(.A1(new_n805), .A2(new_n807), .A3(new_n810), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n784), .A2(new_n791), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n740), .B2(new_n741), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n775), .A2(new_n776), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT96), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n816), .A2(new_n464), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT91), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n626), .A2(G139), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT25), .Z(new_n821));
  NAND3_X1  g396(.A1(new_n818), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT92), .Z(new_n823));
  MUX2_X1   g398(.A(G33), .B(new_n823), .S(G29), .Z(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT93), .B(G2072), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n742), .A2(new_n813), .A3(new_n815), .A4(new_n826), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n800), .A2(G2067), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n827), .A2(new_n829), .ZN(G311));
  INV_X1    g405(.A(G311), .ZN(G150));
  NAND2_X1  g406(.A1(new_n536), .A2(G93), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n538), .A2(G55), .ZN(new_n833));
  AOI22_X1  g408(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n832), .B(new_n833), .C1(new_n514), .C2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(G860), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT37), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n609), .A2(G559), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT38), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT39), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT101), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n835), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n835), .A2(new_n841), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n842), .A2(new_n621), .A3(new_n843), .ZN(new_n844));
  OR3_X1    g419(.A1(new_n835), .A2(new_n621), .A3(new_n841), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n840), .B(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n837), .B1(new_n848), .B2(G860), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT102), .Z(G145));
  INV_X1    g425(.A(G37), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n735), .B(new_n634), .Z(new_n852));
  NAND2_X1  g427(.A1(new_n475), .A2(G130), .ZN(new_n853));
  INV_X1    g428(.A(G142), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n464), .A2(G118), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT104), .ZN(new_n856));
  OAI21_X1  g431(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n857));
  OAI221_X1 g432(.A(new_n853), .B1(new_n487), .B2(new_n854), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n852), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n852), .A2(new_n858), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT105), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT105), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n859), .B2(new_n860), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n797), .B(new_n500), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n774), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n822), .A2(KEYINPUT103), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n867), .B(new_n823), .C1(KEYINPUT92), .C2(KEYINPUT103), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n865), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n630), .B(G160), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(G162), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n861), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n872), .B(new_n875), .C1(new_n871), .C2(new_n876), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n862), .A2(new_n869), .A3(new_n870), .A4(new_n864), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n872), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(KEYINPUT106), .B1(new_n879), .B2(new_n874), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT106), .ZN(new_n881));
  AOI211_X1 g456(.A(new_n881), .B(new_n875), .C1(new_n872), .C2(new_n878), .ZN(new_n882));
  OAI211_X1 g457(.A(new_n851), .B(new_n877), .C1(new_n880), .C2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g459(.A1(new_n835), .A2(new_n613), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n702), .A2(new_n703), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(new_n724), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n704), .A2(G290), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(KEYINPUT108), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT108), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n887), .A2(new_n891), .A3(new_n888), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n590), .B(new_n520), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n890), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n893), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n889), .A2(KEYINPUT108), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT42), .ZN(new_n898));
  XOR2_X1   g473(.A(KEYINPUT107), .B(KEYINPUT41), .Z(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n608), .A2(G299), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n608), .A2(G299), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n902), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n903), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n846), .B(new_n623), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(new_n905), .B2(new_n908), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n898), .B(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n885), .B1(new_n911), .B2(new_n613), .ZN(G295));
  OAI21_X1  g487(.A(new_n885), .B1(new_n911), .B2(new_n613), .ZN(G331));
  INV_X1    g488(.A(KEYINPUT109), .ZN(new_n914));
  NAND2_X1  g489(.A1(G171), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(G301), .A2(KEYINPUT109), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(G286), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(G168), .A2(G171), .A3(new_n914), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n846), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT110), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n844), .A2(new_n917), .A3(new_n845), .A4(new_n918), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n847), .A2(KEYINPUT110), .A3(new_n918), .A4(new_n917), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n920), .A2(new_n922), .ZN(new_n926));
  OAI22_X1  g501(.A1(new_n925), .A2(new_n907), .B1(new_n904), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT111), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI221_X1 g504(.A(KEYINPUT111), .B1(new_n904), .B2(new_n926), .C1(new_n925), .C2(new_n907), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(new_n930), .A3(new_n897), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n926), .A2(new_n904), .ZN(new_n932));
  INV_X1    g507(.A(new_n925), .ZN(new_n933));
  INV_X1    g508(.A(new_n907), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n894), .A2(new_n896), .ZN(new_n936));
  AOI21_X1  g511(.A(G37), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n931), .A2(new_n937), .A3(KEYINPUT43), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT43), .ZN(new_n939));
  AOI22_X1  g514(.A1(new_n905), .A2(new_n899), .B1(new_n920), .B2(new_n922), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n905), .B1(new_n925), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(KEYINPUT41), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n936), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n851), .B1(new_n927), .B2(new_n897), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n939), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n938), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n931), .A2(new_n937), .A3(new_n939), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT43), .B1(new_n943), .B2(new_n944), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(new_n950), .A3(KEYINPUT44), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT112), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n951), .A2(new_n952), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n948), .B1(new_n953), .B2(new_n954), .ZN(G397));
  INV_X1    g530(.A(G1384), .ZN(new_n956));
  INV_X1    g531(.A(new_n492), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n957), .B1(new_n465), .B2(G126), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n495), .B1(new_n958), .B2(new_n464), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n498), .A2(new_n499), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n956), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT45), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n466), .A2(new_n468), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(G2105), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n470), .A2(new_n471), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(new_n464), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n965), .A2(new_n967), .A3(G40), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n963), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n969), .B(KEYINPUT113), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G2067), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n797), .B(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G1996), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n973), .B1(new_n974), .B2(new_n774), .ZN(new_n975));
  INV_X1    g550(.A(new_n969), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n976), .A2(G1996), .ZN(new_n977));
  AOI22_X1  g552(.A1(new_n971), .A2(new_n975), .B1(new_n774), .B2(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n978), .A2(new_n738), .A3(new_n734), .A4(new_n727), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n798), .A2(new_n972), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n970), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n977), .B(KEYINPUT46), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n970), .B1(new_n774), .B2(new_n973), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n984), .B(KEYINPUT47), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n735), .B(new_n737), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n986), .B(KEYINPUT114), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n971), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n988), .A2(new_n978), .ZN(new_n989));
  NOR3_X1   g564(.A1(new_n976), .A2(G1986), .A3(G290), .ZN(new_n990));
  XOR2_X1   g565(.A(new_n990), .B(KEYINPUT48), .Z(new_n991));
  AOI211_X1 g566(.A(new_n981), .B(new_n985), .C1(new_n989), .C2(new_n991), .ZN(new_n992));
  XOR2_X1   g567(.A(KEYINPUT58), .B(G1341), .Z(new_n993));
  OAI21_X1  g568(.A(new_n993), .B1(new_n961), .B2(new_n968), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT120), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G40), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n469), .A2(new_n472), .A3(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n500), .A2(KEYINPUT45), .A3(new_n956), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n963), .A2(new_n974), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  OAI211_X1 g575(.A(KEYINPUT120), .B(new_n993), .C1(new_n961), .C2(new_n968), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n996), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n546), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT59), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT59), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1002), .A2(new_n1005), .A3(new_n546), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT50), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1008), .B(new_n956), .C1(new_n959), .C2(new_n960), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n998), .ZN(new_n1010));
  XNOR2_X1  g585(.A(KEYINPUT115), .B(KEYINPUT50), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1012), .B1(new_n500), .B2(new_n956), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n789), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g589(.A(KEYINPUT56), .B(G2072), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n963), .A2(new_n998), .A3(new_n999), .A4(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT57), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n556), .A2(new_n561), .A3(new_n1018), .A4(new_n565), .ZN(new_n1019));
  AOI22_X1  g594(.A1(new_n1014), .A2(new_n1016), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT121), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT61), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1014), .A2(new_n1016), .A3(new_n1017), .A4(new_n1019), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1022), .A2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1025), .A2(new_n1021), .A3(KEYINPUT61), .A4(new_n1026), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1007), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT122), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1007), .A2(new_n1028), .A3(KEYINPUT122), .A4(new_n1029), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT116), .B1(new_n961), .B2(new_n1011), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT116), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n500), .A2(new_n1035), .A3(new_n956), .A4(new_n1012), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n968), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n961), .A2(KEYINPUT50), .ZN(new_n1038));
  AOI21_X1  g613(.A(G1348), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n961), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n998), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1041), .A2(G2067), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1039), .A2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n608), .B1(new_n1043), .B2(KEYINPUT60), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT60), .ZN(new_n1045));
  NOR4_X1   g620(.A1(new_n1039), .A2(new_n609), .A3(new_n1045), .A4(new_n1042), .ZN(new_n1046));
  OAI22_X1  g621(.A1(new_n1044), .A2(new_n1046), .B1(KEYINPUT60), .B2(new_n1043), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1032), .A2(new_n1033), .A3(new_n1047), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n609), .B(new_n1026), .C1(new_n1039), .C2(new_n1042), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n1049), .A2(new_n1025), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  XOR2_X1   g626(.A(KEYINPUT117), .B(G8), .Z(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1054));
  INV_X1    g629(.A(G2084), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1054), .A2(new_n1055), .A3(new_n998), .A4(new_n1038), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n963), .A2(new_n998), .A3(new_n999), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(new_n804), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1053), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(G168), .A2(new_n1053), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1059), .A2(KEYINPUT51), .A3(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g636(.A(new_n1061), .B(KEYINPUT124), .ZN(new_n1062));
  INV_X1    g637(.A(G8), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1063), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT123), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1060), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1067), .B1(new_n1064), .B2(KEYINPUT123), .ZN(new_n1068));
  OAI21_X1  g643(.A(KEYINPUT51), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(new_n1052), .ZN(new_n1072));
  OAI22_X1  g647(.A1(new_n1062), .A2(new_n1070), .B1(G168), .B2(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g648(.A(G301), .B(KEYINPUT54), .ZN(new_n1074));
  AOI21_X1  g649(.A(G1961), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT53), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n963), .A2(new_n999), .ZN(new_n1077));
  INV_X1    g652(.A(G2078), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(new_n1078), .A3(new_n998), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1075), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT53), .B1(new_n968), .B2(KEYINPUT125), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1081), .B1(KEYINPUT125), .B2(new_n968), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1082), .A2(new_n1078), .A3(new_n1077), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1074), .B1(new_n1080), .B2(new_n1083), .ZN(new_n1084));
  OR2_X1    g659(.A1(new_n1079), .A2(new_n1076), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1080), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1084), .B1(new_n1086), .B2(new_n1074), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT118), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n536), .A2(G86), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1089), .A2(new_n579), .A3(new_n584), .A4(new_n586), .ZN(new_n1090));
  AND2_X1   g665(.A1(new_n1090), .A2(G1981), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n587), .A2(G1981), .A3(new_n589), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1088), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT49), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1041), .A2(new_n1052), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT49), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1088), .B(new_n1097), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1094), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G1976), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT52), .B1(G288), .B2(new_n1100), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1096), .B(new_n1101), .C1(new_n886), .C2(new_n1100), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1100), .B1(new_n702), .B2(new_n703), .ZN(new_n1103));
  OAI21_X1  g678(.A(KEYINPUT52), .B1(new_n1103), .B2(new_n1095), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1099), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(G2090), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1054), .A2(new_n1107), .A3(new_n998), .A4(new_n1038), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1057), .A2(new_n713), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT55), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1111), .B1(G303), .B2(G8), .ZN(new_n1112));
  AOI211_X1 g687(.A(KEYINPUT55), .B(new_n1063), .C1(new_n568), .C2(new_n570), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1110), .A2(G8), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1114), .ZN(new_n1116));
  NOR3_X1   g691(.A1(new_n1010), .A2(new_n1013), .A3(G2090), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1117), .B1(new_n713), .B2(new_n1057), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1116), .B1(new_n1118), .B2(new_n1053), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1106), .A2(KEYINPUT126), .A3(new_n1115), .A4(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT126), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1121), .B1(new_n1105), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1087), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1051), .A2(new_n1073), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT127), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1072), .A2(G286), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1063), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1106), .B(new_n1127), .C1(new_n1114), .C2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT63), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT63), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1127), .A2(new_n1131), .A3(new_n1119), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(new_n1115), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n1106), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1095), .B(KEYINPUT119), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1136), .A2(G288), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1135), .B1(new_n1137), .B2(new_n1092), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1130), .A2(new_n1134), .A3(new_n1138), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1125), .A2(new_n1126), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1126), .B1(new_n1125), .B2(new_n1139), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(new_n1073), .B2(KEYINPUT62), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1086), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1072), .A2(G168), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1059), .A2(KEYINPUT51), .ZN(new_n1146));
  AOI21_X1  g721(.A(KEYINPUT124), .B1(new_n1146), .B2(new_n1067), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT124), .ZN(new_n1148));
  NOR4_X1   g723(.A1(new_n1059), .A2(new_n1148), .A3(KEYINPUT51), .A4(new_n1060), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1145), .B1(new_n1150), .B2(new_n1069), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT62), .ZN(new_n1152));
  OAI211_X1 g727(.A(G171), .B(new_n1144), .C1(new_n1151), .C2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1143), .A2(new_n1153), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1140), .A2(new_n1141), .A3(new_n1154), .ZN(new_n1155));
  XOR2_X1   g730(.A(G290), .B(G1986), .Z(new_n1156));
  OAI21_X1  g731(.A(new_n989), .B1(new_n976), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n992), .B1(new_n1155), .B2(new_n1157), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g733(.A1(new_n946), .A2(new_n883), .A3(G319), .ZN(new_n1160));
  INV_X1    g734(.A(G227), .ZN(new_n1161));
  NAND4_X1  g735(.A1(new_n660), .A2(new_n697), .A3(new_n699), .A4(new_n1161), .ZN(new_n1162));
  NOR2_X1   g736(.A1(new_n1160), .A2(new_n1162), .ZN(G308));
  AND4_X1   g737(.A1(new_n660), .A2(new_n697), .A3(new_n699), .A4(new_n1161), .ZN(new_n1164));
  NAND4_X1  g738(.A1(new_n1164), .A2(G319), .A3(new_n883), .A4(new_n946), .ZN(G225));
endmodule


