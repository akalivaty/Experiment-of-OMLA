//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 0 1 0 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1283, new_n1284, new_n1285,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT64), .Z(new_n208));
  AOI22_X1  g0008(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n211));
  NAND3_X1  g0011(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n206), .B1(new_n208), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT65), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT1), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n215), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n206), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT0), .Z(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n221), .A2(new_n204), .ZN(new_n222));
  OAI21_X1  g0022(.A(G50), .B1(G58), .B2(G68), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n220), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n216), .A2(new_n217), .A3(new_n225), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT66), .Z(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n230), .B(new_n231), .Z(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G107), .B(G116), .Z(new_n237));
  XNOR2_X1  g0037(.A(G87), .B(G97), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  INV_X1    g0039(.A(G50), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(G68), .ZN(new_n241));
  INV_X1    g0041(.A(G68), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n239), .B(new_n246), .ZN(G351));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n221), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT8), .B(G58), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(G20), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G150), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n204), .A2(new_n251), .ZN(new_n255));
  OAI22_X1  g0055(.A1(new_n250), .A2(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G58), .A2(G68), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n204), .B1(new_n257), .B2(new_n240), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n249), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(new_n249), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n204), .A2(G1), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(new_n240), .ZN(new_n264));
  AOI22_X1  g0064(.A1(new_n262), .A2(new_n264), .B1(new_n240), .B2(new_n261), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n259), .A2(new_n265), .ZN(new_n266));
  XOR2_X1   g0066(.A(new_n266), .B(KEYINPUT70), .Z(new_n267));
  INV_X1    g0067(.A(KEYINPUT9), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n267), .B(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G41), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT68), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n221), .ZN(new_n273));
  NAND3_X1  g0073(.A1(KEYINPUT68), .A2(G33), .A3(G41), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G41), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT67), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT67), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G41), .ZN(new_n279));
  INV_X1    g0079(.A(G45), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n277), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n275), .A2(new_n281), .A3(new_n203), .A4(G274), .ZN(new_n282));
  INV_X1    g0082(.A(G226), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n275), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT3), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G1698), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n291), .A2(G223), .B1(G77), .B2(new_n289), .ZN(new_n292));
  AND2_X1   g0092(.A1(new_n287), .A2(new_n288), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n293), .A2(G222), .A3(new_n290), .ZN(new_n294));
  AND2_X1   g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n273), .A2(new_n270), .ZN(new_n296));
  OAI221_X1 g0096(.A(new_n282), .B1(new_n283), .B2(new_n285), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G190), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n299), .B1(G200), .B2(new_n297), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n269), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n301), .B(KEYINPUT10), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n297), .A2(G179), .ZN(new_n303));
  INV_X1    g0103(.A(G169), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n297), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n303), .A2(new_n266), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G244), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n291), .A2(G238), .B1(G107), .B2(new_n289), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n293), .A2(G232), .A3(new_n290), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI221_X1 g0110(.A(new_n282), .B1(new_n307), .B2(new_n285), .C1(new_n310), .C2(new_n296), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G200), .ZN(new_n312));
  INV_X1    g0112(.A(new_n262), .ZN(new_n313));
  OAI21_X1  g0113(.A(G77), .B1(new_n204), .B2(G1), .ZN(new_n314));
  OAI22_X1  g0114(.A1(new_n313), .A2(new_n314), .B1(G77), .B2(new_n260), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT69), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n250), .B1(new_n316), .B2(new_n255), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(new_n316), .B2(new_n255), .ZN(new_n318));
  INV_X1    g0118(.A(G77), .ZN(new_n319));
  XNOR2_X1  g0119(.A(KEYINPUT15), .B(G87), .ZN(new_n320));
  OAI221_X1 g0120(.A(new_n318), .B1(new_n204), .B2(new_n319), .C1(new_n253), .C2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n315), .B1(new_n321), .B2(new_n249), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n312), .B(new_n322), .C1(new_n298), .C2(new_n311), .ZN(new_n323));
  OR2_X1    g0123(.A1(new_n311), .A2(G179), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n322), .B1(new_n304), .B2(new_n311), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n302), .A2(new_n306), .A3(new_n323), .A4(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n282), .B1(new_n229), .B2(new_n285), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT76), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n251), .A2(KEYINPUT72), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT72), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(G33), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n331), .A2(new_n333), .A3(KEYINPUT3), .ZN(new_n334));
  OAI21_X1  g0134(.A(KEYINPUT73), .B1(new_n251), .B2(KEYINPUT3), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT73), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(new_n286), .A3(G33), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n334), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n283), .A2(G1698), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n339), .B1(G223), .B2(G1698), .ZN(new_n340));
  INV_X1    g0140(.A(G87), .ZN(new_n341));
  OAI22_X1  g0141(.A1(new_n338), .A2(new_n340), .B1(new_n251), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n296), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n282), .B(KEYINPUT76), .C1(new_n229), .C2(new_n285), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n330), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G169), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n328), .A2(new_n329), .B1(new_n342), .B2(new_n343), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n348), .A2(G179), .A3(new_n345), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  AND2_X1   g0150(.A1(G58), .A2(G68), .ZN(new_n351));
  OAI21_X1  g0151(.A(G20), .B1(new_n351), .B2(new_n257), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT74), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n204), .A2(new_n251), .A3(G159), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n353), .B1(new_n352), .B2(new_n354), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT7), .ZN(new_n359));
  AND3_X1   g0159(.A1(new_n331), .A2(new_n333), .A3(KEYINPUT3), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n335), .A2(new_n337), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n359), .B(new_n204), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G68), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n359), .B1(new_n338), .B2(new_n204), .ZN(new_n364));
  OAI211_X1 g0164(.A(KEYINPUT16), .B(new_n358), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT16), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n359), .A2(G20), .ZN(new_n367));
  AOI21_X1  g0167(.A(KEYINPUT3), .B1(new_n331), .B2(new_n333), .ZN(new_n368));
  INV_X1    g0168(.A(new_n288), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n359), .B1(new_n293), .B2(G20), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n242), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n352), .A2(new_n354), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT74), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n355), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n366), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n365), .A2(new_n376), .A3(new_n249), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n250), .A2(new_n263), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n313), .B1(KEYINPUT75), .B2(new_n378), .ZN(new_n379));
  OR2_X1    g0179(.A1(new_n378), .A2(KEYINPUT75), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n379), .A2(new_n380), .B1(new_n261), .B2(new_n250), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n350), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT18), .ZN(new_n384));
  INV_X1    g0184(.A(new_n382), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n346), .A2(G200), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n298), .A2(KEYINPUT77), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n298), .A2(KEYINPUT77), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n348), .A2(new_n345), .A3(new_n390), .ZN(new_n391));
  AND2_X1   g0191(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n385), .A2(new_n392), .A3(KEYINPUT17), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT18), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n350), .A2(new_n382), .A3(new_n394), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n386), .A2(new_n377), .A3(new_n391), .A4(new_n381), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT17), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n384), .A2(new_n393), .A3(new_n395), .A4(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT71), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n291), .A2(G232), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G33), .A2(G97), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n293), .A2(G226), .A3(new_n290), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n343), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT13), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n275), .A2(new_n284), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G238), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n405), .A2(new_n406), .A3(new_n282), .A4(new_n408), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n291), .A2(G232), .B1(G33), .B2(G97), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n296), .B1(new_n410), .B2(new_n403), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n408), .A2(new_n282), .ZN(new_n412));
  OAI21_X1  g0212(.A(KEYINPUT13), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n409), .A2(new_n413), .A3(G190), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n261), .A2(new_n242), .ZN(new_n415));
  XNOR2_X1  g0215(.A(new_n415), .B(KEYINPUT12), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n242), .A2(G20), .ZN(new_n417));
  OAI221_X1 g0217(.A(new_n417), .B1(new_n240), .B2(new_n255), .C1(new_n253), .C2(new_n319), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n418), .A2(KEYINPUT11), .A3(new_n249), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n262), .B(G68), .C1(G1), .C2(new_n204), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n416), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT11), .B1(new_n418), .B2(new_n249), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n414), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(G200), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(new_n409), .B2(new_n413), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n400), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n426), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n428), .A2(KEYINPUT71), .A3(new_n414), .A4(new_n423), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n423), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n409), .A2(new_n413), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT14), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n432), .A2(new_n433), .A3(G169), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n409), .A2(new_n413), .A3(G179), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n304), .B1(new_n409), .B2(new_n413), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n437), .A2(new_n433), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n431), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n430), .A2(new_n439), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n327), .A2(new_n399), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT4), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(new_n307), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n444), .A2(new_n290), .A3(new_n287), .A4(new_n288), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n287), .A2(new_n288), .A3(G250), .A4(G1698), .ZN(new_n446));
  NAND2_X1  g0246(.A1(G33), .A2(G283), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n307), .A2(G1698), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n334), .A2(new_n335), .A3(new_n337), .A4(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n443), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT79), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n448), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n450), .A2(KEYINPUT79), .A3(new_n443), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n296), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT5), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n278), .A2(G41), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n276), .A2(KEYINPUT67), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n456), .A2(G41), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n203), .A2(G45), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n459), .A2(G274), .A3(new_n275), .A4(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(KEYINPUT5), .B1(new_n277), .B2(new_n279), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n203), .B(G45), .C1(new_n456), .C2(G41), .ZN(new_n465));
  OAI211_X1 g0265(.A(G257), .B(new_n275), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n304), .B1(new_n455), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT80), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n463), .A2(new_n466), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n469), .B1(new_n463), .B2(new_n466), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(G179), .ZN(new_n473));
  AND3_X1   g0273(.A1(new_n450), .A2(KEYINPUT79), .A3(new_n443), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT79), .B1(new_n450), .B2(new_n443), .ZN(new_n475));
  NOR3_X1   g0275(.A1(new_n474), .A2(new_n475), .A3(new_n448), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n472), .B(new_n473), .C1(new_n476), .C2(new_n296), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT6), .ZN(new_n478));
  AND2_X1   g0278(.A1(G97), .A2(G107), .ZN(new_n479));
  NOR2_X1   g0279(.A1(G97), .A2(G107), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(KEYINPUT6), .A2(G97), .ZN(new_n482));
  OAI21_X1  g0282(.A(KEYINPUT78), .B1(new_n482), .B2(G107), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT78), .ZN(new_n484));
  INV_X1    g0284(.A(G107), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n484), .A2(new_n485), .A3(KEYINPUT6), .A4(G97), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n481), .A2(new_n483), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G20), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(new_n319), .B2(new_n255), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n485), .B1(new_n370), .B2(new_n371), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n249), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n260), .A2(G97), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n203), .A2(G33), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n260), .A2(new_n493), .A3(new_n221), .A4(new_n248), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n492), .B1(new_n495), .B2(G97), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n468), .A2(new_n477), .A3(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n280), .A2(G1), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n275), .A2(G274), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n331), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n251), .A2(KEYINPUT72), .ZN(new_n503));
  OAI21_X1  g0303(.A(G116), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(G238), .A2(G1698), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n505), .B1(new_n307), .B2(G1698), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n504), .B1(new_n338), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n501), .B1(new_n508), .B2(new_n343), .ZN(new_n509));
  INV_X1    g0309(.A(G250), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n499), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n275), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT82), .ZN(new_n513));
  XNOR2_X1  g0313(.A(new_n512), .B(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n509), .A2(G190), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n425), .B1(new_n509), .B2(new_n514), .ZN(new_n516));
  AOI21_X1  g0316(.A(KEYINPUT19), .B1(new_n252), .B2(G97), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n341), .A2(KEYINPUT83), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT83), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(G87), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n518), .A2(new_n520), .A3(new_n480), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT19), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n522), .B1(new_n402), .B2(new_n204), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n517), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n334), .A2(new_n204), .A3(new_n335), .A4(new_n337), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n524), .B1(new_n525), .B2(new_n242), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n249), .ZN(new_n527));
  INV_X1    g0327(.A(new_n320), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n528), .A2(new_n260), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n494), .A2(new_n341), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n527), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n516), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n509), .A2(G179), .A3(new_n514), .ZN(new_n535));
  XNOR2_X1  g0335(.A(new_n512), .B(KEYINPUT82), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n335), .A2(new_n337), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n537), .A2(new_n334), .A3(new_n506), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n296), .B1(new_n538), .B2(new_n504), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n536), .A2(new_n539), .A3(new_n501), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n535), .B1(new_n540), .B2(new_n304), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n494), .A2(new_n320), .ZN(new_n542));
  XNOR2_X1  g0342(.A(new_n542), .B(KEYINPUT84), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n527), .A2(new_n530), .A3(new_n543), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n515), .A2(new_n534), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n451), .A2(new_n452), .ZN(new_n546));
  INV_X1    g0346(.A(new_n448), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n546), .A2(new_n454), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n467), .B1(new_n548), .B2(new_n343), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n497), .B1(new_n549), .B2(G190), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n467), .A2(KEYINPUT80), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n463), .A2(new_n466), .A3(new_n469), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(G200), .B1(new_n455), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(KEYINPUT81), .B1(new_n550), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n497), .ZN(new_n556));
  INV_X1    g0356(.A(new_n467), .ZN(new_n557));
  OAI211_X1 g0357(.A(G190), .B(new_n557), .C1(new_n476), .C2(new_n296), .ZN(new_n558));
  AND4_X1   g0358(.A1(KEYINPUT81), .A2(new_n554), .A3(new_n556), .A4(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n498), .B(new_n545), .C1(new_n555), .C2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n261), .A2(KEYINPUT25), .A3(new_n485), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(KEYINPUT25), .B1(new_n261), .B2(new_n485), .ZN(new_n563));
  OAI22_X1  g0363(.A1(new_n562), .A2(new_n563), .B1(new_n485), .B2(new_n494), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT22), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n566), .A2(new_n341), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n537), .A2(new_n204), .A3(new_n334), .A4(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n204), .A2(G87), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n566), .B1(new_n289), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n485), .A2(G20), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT23), .ZN(new_n573));
  XNOR2_X1  g0373(.A(new_n572), .B(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n204), .B(G116), .C1(new_n502), .C2(new_n503), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n571), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(KEYINPUT87), .B1(new_n569), .B2(new_n576), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n574), .A2(new_n575), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT87), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n578), .A2(new_n568), .A3(new_n579), .A4(new_n571), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n577), .A2(new_n580), .A3(KEYINPUT24), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n249), .B1(new_n577), .B2(KEYINPUT24), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n565), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(G294), .B1(new_n502), .B2(new_n503), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n510), .A2(new_n290), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(G257), .B2(new_n290), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n584), .B1(new_n338), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n343), .ZN(new_n588));
  OAI211_X1 g0388(.A(G264), .B(new_n275), .C1(new_n464), .C2(new_n465), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n588), .A2(new_n463), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(KEYINPUT88), .ZN(new_n591));
  XNOR2_X1  g0391(.A(KEYINPUT67), .B(G41), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n462), .B1(KEYINPUT5), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT88), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n593), .A2(new_n594), .A3(G264), .A4(new_n275), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n596), .A2(new_n588), .A3(new_n463), .ZN(new_n597));
  OAI22_X1  g0397(.A1(new_n590), .A2(new_n304), .B1(new_n597), .B2(new_n473), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n583), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n425), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n588), .A2(new_n298), .A3(new_n463), .A4(new_n589), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n577), .A2(new_n580), .A3(KEYINPUT24), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n571), .A2(new_n574), .A3(new_n575), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n579), .B1(new_n604), .B2(new_n568), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT24), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n603), .A2(new_n607), .A3(new_n249), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n602), .A2(new_n608), .A3(new_n565), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n599), .A2(new_n609), .ZN(new_n610));
  OR2_X1    g0410(.A1(G257), .A2(G1698), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(G264), .B2(new_n290), .ZN(new_n612));
  INV_X1    g0412(.A(G303), .ZN(new_n613));
  OAI22_X1  g0413(.A1(new_n338), .A2(new_n612), .B1(new_n613), .B2(new_n293), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n343), .ZN(new_n615));
  OAI211_X1 g0415(.A(G270), .B(new_n275), .C1(new_n464), .C2(new_n465), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n463), .A2(new_n616), .A3(KEYINPUT85), .ZN(new_n617));
  AOI21_X1  g0417(.A(KEYINPUT85), .B1(new_n463), .B2(new_n616), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n615), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(G97), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n447), .B(new_n204), .C1(G33), .C2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(G116), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(G20), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n621), .A2(new_n249), .A3(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT20), .ZN(new_n625));
  OR2_X1    g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(KEYINPUT86), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n260), .A2(new_n622), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(new_n495), .B2(new_n622), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT86), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n624), .A2(new_n631), .A3(new_n625), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n628), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n619), .A2(G169), .A3(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT21), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n633), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n390), .B(new_n615), .C1(new_n617), .C2(new_n618), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n463), .A2(new_n616), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT85), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n463), .A2(new_n616), .A3(KEYINPUT85), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n641), .A2(new_n642), .B1(new_n343), .B2(new_n614), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n637), .B(new_n638), .C1(new_n643), .C2(new_n425), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(G179), .A3(new_n633), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n619), .A2(new_n633), .A3(KEYINPUT21), .A4(G169), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n636), .A2(new_n644), .A3(new_n645), .A4(new_n646), .ZN(new_n647));
  NOR4_X1   g0447(.A1(new_n442), .A2(new_n560), .A3(new_n610), .A4(new_n647), .ZN(G372));
  INV_X1    g0448(.A(new_n306), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n393), .A2(new_n398), .ZN(new_n650));
  INV_X1    g0450(.A(new_n439), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n326), .B1(new_n427), .B2(new_n429), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n395), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n394), .B1(new_n350), .B2(new_n382), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n649), .B1(new_n657), .B2(new_n302), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n509), .A2(G179), .A3(new_n514), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n304), .B1(new_n509), .B2(new_n514), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n544), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AOI211_X1 g0461(.A(new_n529), .B(new_n531), .C1(new_n526), .C2(new_n249), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n662), .B(new_n515), .C1(new_n540), .C2(new_n425), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n468), .A2(new_n477), .A3(new_n497), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n554), .A2(new_n556), .A3(new_n558), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT81), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n550), .A2(KEYINPUT81), .A3(new_n554), .ZN(new_n669));
  AOI211_X1 g0469(.A(new_n664), .B(new_n665), .C1(new_n668), .C2(new_n669), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n645), .A2(new_n646), .ZN(new_n671));
  AOI21_X1  g0471(.A(KEYINPUT89), .B1(new_n671), .B2(new_n636), .ZN(new_n672));
  AND4_X1   g0472(.A1(KEYINPUT89), .A2(new_n636), .A3(new_n645), .A4(new_n646), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n599), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n670), .A2(new_n674), .A3(new_n609), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT90), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n545), .A2(new_n665), .A3(KEYINPUT26), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT26), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n664), .B2(new_n498), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n676), .B1(new_n680), .B2(new_n661), .ZN(new_n681));
  INV_X1    g0481(.A(new_n661), .ZN(new_n682));
  AOI211_X1 g0482(.A(KEYINPUT90), .B(new_n682), .C1(new_n677), .C2(new_n679), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n675), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n658), .B1(new_n442), .B2(new_n685), .ZN(G369));
  NAND3_X1  g0486(.A1(new_n203), .A2(new_n204), .A3(G13), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n687), .A2(KEYINPUT27), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(KEYINPUT27), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n688), .A2(G213), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G343), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n691), .B(KEYINPUT91), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n633), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n647), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n672), .A2(new_n673), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n695), .B1(new_n696), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT92), .ZN(new_n698));
  XNOR2_X1  g0498(.A(KEYINPUT93), .B(G330), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n599), .A2(new_n609), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n583), .A2(new_n693), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n583), .A2(new_n598), .A3(new_n693), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n701), .A2(new_n707), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n671), .A2(new_n636), .ZN(new_n709));
  OR2_X1    g0509(.A1(new_n709), .A2(new_n693), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n710), .A2(new_n610), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n599), .B2(new_n693), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  XOR2_X1   g0513(.A(new_n713), .B(KEYINPUT94), .Z(G399));
  NAND2_X1  g0514(.A1(new_n218), .A2(new_n592), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n521), .A2(G116), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n715), .A2(G1), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(new_n223), .B2(new_n715), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT28), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n684), .A2(new_n692), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n720), .A2(KEYINPUT29), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n709), .A2(new_n599), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n670), .A2(new_n609), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n682), .B1(new_n677), .B2(new_n679), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n693), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(KEYINPUT29), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n721), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT97), .ZN(new_n728));
  INV_X1    g0528(.A(new_n647), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n702), .A2(new_n729), .A3(new_n692), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n728), .B1(new_n730), .B2(new_n560), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n610), .A2(new_n647), .A3(new_n693), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n665), .B1(new_n668), .B2(new_n669), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n732), .A2(KEYINPUT97), .A3(new_n733), .A4(new_n545), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  OAI211_X1 g0535(.A(G179), .B(new_n615), .C1(new_n617), .C2(new_n618), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n508), .A2(new_n343), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n514), .A2(new_n738), .A3(new_n500), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n596), .A2(new_n588), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n737), .A2(new_n741), .A3(KEYINPUT30), .A4(new_n549), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(KEYINPUT96), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n509), .A2(new_n596), .A3(new_n514), .A4(new_n588), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n744), .A2(new_n455), .A3(new_n467), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT96), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n745), .A2(new_n746), .A3(KEYINPUT30), .A4(new_n737), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n743), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n737), .A2(new_n741), .A3(new_n549), .ZN(new_n749));
  XOR2_X1   g0549(.A(KEYINPUT95), .B(KEYINPUT30), .Z(new_n750));
  AND4_X1   g0550(.A1(new_n473), .A2(new_n619), .A3(new_n597), .A4(new_n739), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n472), .B1(new_n476), .B2(new_n296), .ZN(new_n752));
  AOI22_X1  g0552(.A1(new_n749), .A2(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n748), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(KEYINPUT31), .B1(new_n754), .B2(new_n693), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT31), .ZN(new_n756));
  AOI211_X1 g0556(.A(new_n756), .B(new_n692), .C1(new_n748), .C2(new_n753), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n699), .B1(new_n735), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n727), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n719), .B1(new_n760), .B2(G1), .ZN(G364));
  INV_X1    g0561(.A(new_n701), .ZN(new_n762));
  INV_X1    g0562(.A(new_n715), .ZN(new_n763));
  INV_X1    g0563(.A(G13), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(G20), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n203), .B1(new_n765), .B2(G45), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n762), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n769), .B1(new_n700), .B2(new_n698), .ZN(new_n770));
  INV_X1    g0570(.A(new_n338), .ZN(new_n771));
  INV_X1    g0571(.A(new_n218), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n224), .A2(new_n280), .ZN(new_n774));
  OAI211_X1 g0574(.A(new_n773), .B(new_n774), .C1(new_n280), .C2(new_n246), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n772), .A2(new_n289), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n776), .A2(G355), .B1(new_n622), .B2(new_n772), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n778), .A2(KEYINPUT98), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G13), .A2(G33), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(G20), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n221), .B1(G20), .B2(new_n304), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n784), .B1(new_n778), .B2(KEYINPUT98), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n768), .B1(new_n779), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n204), .A2(G179), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n787), .A2(new_n298), .A3(G200), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n789), .A2(KEYINPUT100), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(KEYINPUT100), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n485), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n204), .A2(new_n473), .A3(G200), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n390), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR3_X1   g0596(.A1(new_n204), .A2(new_n473), .A3(new_n425), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(G190), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n796), .A2(G58), .B1(G68), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(G179), .A2(G200), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n204), .B1(new_n801), .B2(G190), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n620), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n518), .A2(new_n520), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n787), .A2(G190), .A3(G200), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n803), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n801), .A2(G20), .A3(new_n298), .ZN(new_n808));
  INV_X1    g0608(.A(G159), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT32), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n798), .A2(new_n389), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n289), .B1(new_n812), .B2(G50), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n800), .A2(new_n807), .A3(new_n811), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n794), .A2(new_n298), .ZN(new_n815));
  AND2_X1   g0615(.A1(new_n815), .A2(KEYINPUT99), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n815), .A2(KEYINPUT99), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n793), .B(new_n814), .C1(G77), .C2(new_n819), .ZN(new_n820));
  OR2_X1    g0620(.A1(new_n820), .A2(KEYINPUT101), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(KEYINPUT101), .ZN(new_n822));
  INV_X1    g0622(.A(G283), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n792), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n812), .A2(G326), .ZN(new_n825));
  INV_X1    g0625(.A(G294), .ZN(new_n826));
  INV_X1    g0626(.A(G322), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n825), .B1(new_n826), .B2(new_n802), .C1(new_n827), .C2(new_n795), .ZN(new_n828));
  INV_X1    g0628(.A(new_n808), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n293), .B1(G329), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n613), .B2(new_n805), .ZN(new_n831));
  INV_X1    g0631(.A(new_n799), .ZN(new_n832));
  XOR2_X1   g0632(.A(KEYINPUT33), .B(G317), .Z(new_n833));
  INV_X1    g0633(.A(G311), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n832), .A2(new_n833), .B1(new_n815), .B2(new_n834), .ZN(new_n835));
  OR4_X1    g0635(.A1(new_n824), .A2(new_n828), .A3(new_n831), .A4(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n821), .A2(new_n822), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n786), .B1(new_n837), .B2(new_n783), .ZN(new_n838));
  INV_X1    g0638(.A(new_n782), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n838), .B1(new_n698), .B2(new_n839), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n770), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(G396));
  INV_X1    g0642(.A(new_n759), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n326), .A2(new_n693), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n323), .B1(new_n322), .B2(new_n692), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n844), .B1(new_n326), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n684), .A2(new_n692), .A3(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n846), .B1(new_n684), .B2(new_n692), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n843), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n849), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n851), .A2(new_n759), .A3(new_n847), .ZN(new_n852));
  INV_X1    g0652(.A(new_n768), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n850), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n846), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n780), .ZN(new_n856));
  AOI22_X1  g0656(.A1(G137), .A2(new_n812), .B1(new_n799), .B2(G150), .ZN(new_n857));
  INV_X1    g0657(.A(G143), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n857), .B1(new_n858), .B2(new_n795), .C1(new_n818), .C2(new_n809), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT34), .ZN(new_n860));
  INV_X1    g0660(.A(new_n792), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(G68), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n338), .B1(G132), .B2(new_n829), .ZN(new_n863));
  INV_X1    g0663(.A(new_n802), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n806), .A2(G50), .B1(new_n864), .B2(G58), .ZN(new_n865));
  AND4_X1   g0665(.A1(new_n860), .A2(new_n862), .A3(new_n863), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n861), .A2(G87), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n799), .A2(KEYINPUT102), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n799), .A2(KEYINPUT102), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI221_X1 g0671(.A(new_n867), .B1(new_n818), .B2(new_n622), .C1(new_n823), .C2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n289), .B1(new_n808), .B2(new_n834), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n796), .A2(G294), .B1(G107), .B2(new_n806), .ZN(new_n874));
  INV_X1    g0674(.A(new_n812), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n874), .B1(new_n613), .B2(new_n875), .ZN(new_n876));
  NOR4_X1   g0676(.A1(new_n872), .A2(new_n803), .A3(new_n873), .A4(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n783), .B1(new_n866), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n783), .A2(new_n780), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n319), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n856), .A2(new_n768), .A3(new_n878), .A4(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n854), .A2(new_n881), .ZN(G384));
  NOR2_X1   g0682(.A1(new_n765), .A2(new_n203), .ZN(new_n883));
  INV_X1    g0683(.A(new_n690), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n654), .B2(new_n655), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT38), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n365), .A2(new_n249), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n204), .B1(new_n360), .B2(new_n361), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(KEYINPUT7), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n889), .A2(G68), .A3(new_n362), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT16), .B1(new_n890), .B2(new_n358), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n381), .B1(new_n887), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n350), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n690), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n893), .A2(new_n894), .A3(new_n396), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT37), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n382), .A2(new_n690), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT37), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n383), .A2(new_n897), .A3(new_n898), .A4(new_n396), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n896), .A2(KEYINPUT104), .A3(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n894), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n399), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT104), .B1(new_n896), .B2(new_n899), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n886), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT104), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n385), .A2(new_n392), .B1(new_n892), .B2(new_n690), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n898), .B1(new_n907), .B2(new_n893), .ZN(new_n908));
  INV_X1    g0708(.A(new_n899), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n910), .A2(KEYINPUT38), .A3(new_n902), .A4(new_n900), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n905), .A2(KEYINPUT39), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n897), .B1(new_n650), .B2(new_n656), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n383), .A2(new_n897), .A3(new_n396), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(new_n898), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n886), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n911), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n912), .B1(new_n917), .B2(KEYINPUT39), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n651), .A2(new_n692), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n885), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n905), .A2(new_n911), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(KEYINPUT105), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT105), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n905), .A2(new_n923), .A3(new_n911), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n693), .A2(new_n431), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT103), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n926), .B1(new_n440), .B2(new_n927), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n436), .A2(new_n438), .A3(new_n926), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n430), .B(new_n929), .C1(new_n651), .C2(KEYINPUT103), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n844), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n931), .B1(new_n847), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n920), .B1(new_n925), .B2(new_n933), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n441), .B(new_n726), .C1(new_n720), .C2(KEYINPUT29), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n658), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n934), .B(new_n936), .Z(new_n937));
  NAND2_X1  g0737(.A1(new_n735), .A2(new_n758), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n928), .A2(new_n930), .A3(new_n846), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT40), .ZN(new_n941));
  NOR3_X1   g0741(.A1(new_n940), .A2(new_n917), .A3(new_n941), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n938), .A2(new_n939), .ZN(new_n943));
  AND3_X1   g0743(.A1(new_n905), .A2(new_n923), .A3(new_n911), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n923), .B1(new_n905), .B2(new_n911), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n942), .B1(new_n946), .B2(new_n941), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n441), .A2(new_n938), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n699), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n949), .B2(new_n948), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n883), .B1(new_n937), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n937), .B2(new_n951), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n487), .A2(KEYINPUT35), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n487), .A2(KEYINPUT35), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n954), .A2(G116), .A3(new_n222), .A4(new_n955), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT36), .ZN(new_n957));
  INV_X1    g0757(.A(G58), .ZN(new_n958));
  OAI21_X1  g0758(.A(G77), .B1(new_n958), .B2(new_n242), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n241), .B1(new_n959), .B2(new_n223), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n960), .A2(G1), .A3(new_n764), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n953), .A2(new_n957), .A3(new_n961), .ZN(G367));
  INV_X1    g0762(.A(new_n773), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n784), .B1(new_n218), .B2(new_n320), .C1(new_n963), .C2(new_n235), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n853), .B1(new_n964), .B2(KEYINPUT109), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(KEYINPUT109), .B2(new_n964), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n771), .B1(G317), .B2(new_n829), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT46), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n806), .A2(G116), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(new_n968), .B2(new_n969), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n819), .A2(G283), .ZN(new_n972));
  INV_X1    g0772(.A(new_n871), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(G294), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n875), .A2(new_n834), .B1(new_n795), .B2(new_n613), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n788), .A2(new_n620), .B1(new_n802), .B2(new_n485), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n971), .A2(new_n972), .A3(new_n974), .A4(new_n977), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n973), .A2(G159), .B1(G50), .B2(new_n819), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n806), .A2(G58), .B1(new_n829), .B2(G137), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n875), .A2(new_n858), .B1(new_n795), .B2(new_n254), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(G68), .B2(new_n864), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n979), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n293), .B1(new_n788), .B2(new_n319), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT110), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n978), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  XOR2_X1   g0786(.A(KEYINPUT111), .B(KEYINPUT47), .Z(new_n987));
  XNOR2_X1  g0787(.A(new_n986), .B(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n966), .B1(new_n988), .B2(new_n783), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n693), .A2(new_n533), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n664), .B(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n989), .B1(new_n839), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n693), .A2(new_n497), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n733), .A2(new_n995), .B1(new_n665), .B2(new_n693), .ZN(new_n996));
  OAI21_X1  g0796(.A(KEYINPUT42), .B1(new_n711), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n599), .B1(new_n668), .B2(new_n669), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n692), .B1(new_n998), .B2(new_n665), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  NOR3_X1   g0800(.A1(new_n711), .A2(KEYINPUT42), .A3(new_n996), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT106), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1002), .B(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n992), .A2(KEYINPUT43), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n992), .A2(KEYINPUT43), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1004), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n708), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1011), .A2(new_n996), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(KEYINPUT107), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT107), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1010), .A2(new_n1016), .A3(new_n1012), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1013), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n715), .B(KEYINPUT41), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n712), .A2(new_n996), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT44), .Z(new_n1022));
  NOR2_X1   g0822(.A1(new_n712), .A2(new_n996), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT45), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n708), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1022), .A2(new_n1011), .A3(new_n1024), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n707), .A2(new_n710), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n711), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT108), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1030), .B1(new_n701), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n1031), .B2(new_n701), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n762), .A2(KEYINPUT108), .A3(new_n1030), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n760), .A2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1028), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n760), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1020), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n766), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n994), .B1(new_n1018), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(G387));
  INV_X1    g0842(.A(new_n776), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n1043), .A2(new_n716), .B1(G107), .B2(new_n218), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n232), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT113), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n250), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n240), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT50), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n716), .B(new_n280), .C1(new_n242), .C2(new_n319), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n773), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n1045), .A2(G45), .B1(new_n1046), .B2(new_n1051), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1051), .A2(new_n1046), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1044), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n784), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n768), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n875), .A2(new_n809), .B1(new_n319), .B2(new_n805), .ZN(new_n1057));
  XOR2_X1   g0857(.A(KEYINPUT114), .B(G150), .Z(new_n1058));
  INV_X1    g0858(.A(new_n1058), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n338), .B(new_n1057), .C1(new_n829), .C2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n861), .A2(G97), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n796), .A2(G50), .B1(new_n528), .B2(new_n864), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n815), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n799), .A2(new_n1047), .B1(new_n1063), .B2(G68), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .A4(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n771), .B1(G326), .B2(new_n829), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n805), .A2(new_n826), .B1(new_n802), .B2(new_n823), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n796), .A2(G317), .B1(G322), .B2(new_n812), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1068), .B1(new_n613), .B2(new_n818), .C1(new_n871), .C2(new_n834), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT48), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1067), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n1070), .B2(new_n1069), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT49), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1066), .B1(new_n622), .B2(new_n788), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1065), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1056), .B1(new_n1076), .B2(new_n783), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n706), .B2(new_n839), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT115), .ZN(new_n1079));
  OR2_X1    g0879(.A1(new_n760), .A2(new_n1035), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n715), .B1(new_n760), .B2(new_n1035), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1079), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n766), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT112), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1082), .A2(new_n1084), .ZN(G393));
  NAND3_X1  g0885(.A1(new_n1026), .A2(new_n767), .A3(new_n1027), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n996), .A2(new_n782), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n973), .A2(G50), .B1(new_n1047), .B2(new_n819), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n802), .A2(new_n319), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n771), .B1(new_n858), .B2(new_n808), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n1089), .B(new_n1090), .C1(G68), .C2(new_n806), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1088), .A2(new_n867), .A3(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n796), .A2(G159), .B1(G150), .B2(new_n812), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT51), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n796), .A2(G311), .B1(G317), .B2(new_n812), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT52), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n289), .B1(new_n827), .B2(new_n808), .C1(new_n815), .C2(new_n826), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n805), .A2(new_n823), .B1(new_n802), .B2(new_n622), .ZN(new_n1098));
  NOR3_X1   g0898(.A1(new_n793), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n613), .B2(new_n871), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n1092), .A2(new_n1094), .B1(new_n1096), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n783), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n784), .B1(new_n620), .B2(new_n218), .C1(new_n963), .C2(new_n239), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1087), .A2(new_n768), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1086), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT116), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1105), .B(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1037), .A2(new_n715), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1028), .A2(new_n1036), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1107), .A2(new_n1110), .ZN(G390));
  INV_X1    g0911(.A(new_n919), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n918), .B1(new_n933), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n911), .A2(new_n916), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n845), .A2(new_n326), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n844), .B1(new_n725), .B2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n919), .B(new_n1114), .C1(new_n1116), .C2(new_n931), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT117), .ZN(new_n1119));
  AND4_X1   g0919(.A1(new_n1119), .A2(new_n938), .A3(new_n939), .A4(G330), .ZN(new_n1120));
  INV_X1    g0920(.A(G330), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n735), .B2(new_n758), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1119), .B1(new_n1122), .B2(new_n939), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1118), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n931), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n759), .A2(new_n846), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1113), .A2(new_n1117), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n441), .A2(new_n1122), .ZN(new_n1131));
  AND3_X1   g0931(.A1(new_n935), .A2(new_n658), .A3(new_n1131), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n848), .A2(new_n844), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n938), .A2(new_n700), .A3(new_n846), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n931), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1133), .B1(new_n1124), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1122), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n931), .B1(new_n1137), .B2(new_n855), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n1138), .A2(new_n1116), .A3(new_n1128), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1132), .B1(new_n1136), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n715), .B1(new_n1130), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT118), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n935), .A2(new_n658), .A3(new_n1131), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n938), .A2(new_n939), .A3(G330), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(KEYINPUT117), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1122), .A2(new_n1119), .A3(new_n939), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1145), .A2(new_n1135), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1133), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n1128), .A2(new_n1116), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n1138), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1143), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  AND4_X1   g0952(.A1(new_n1142), .A2(new_n1152), .A3(new_n1129), .A4(new_n1126), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n1113), .A2(new_n1117), .A3(new_n1128), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1124), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1142), .B1(new_n1156), .B2(new_n1152), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1141), .B1(new_n1153), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n918), .A2(new_n780), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n879), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n768), .B1(new_n1047), .B2(new_n1160), .ZN(new_n1161));
  XOR2_X1   g0961(.A(new_n1161), .B(KEYINPUT119), .Z(new_n1162));
  NAND2_X1  g0962(.A1(new_n973), .A2(G137), .ZN(new_n1163));
  XOR2_X1   g0963(.A(KEYINPUT54), .B(G143), .Z(new_n1164));
  NAND2_X1  g0964(.A1(new_n819), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n812), .A2(G128), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n796), .A2(G132), .B1(G50), .B2(new_n789), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1163), .A2(new_n1165), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT53), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1059), .A2(new_n806), .A3(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(KEYINPUT53), .B1(new_n1058), .B2(new_n805), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n864), .A2(G159), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n289), .B1(new_n829), .B2(G125), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .A4(new_n1173), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n862), .B1(new_n818), .B2(new_n620), .C1(new_n485), .C2(new_n871), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n796), .A2(G116), .B1(G87), .B2(new_n806), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n293), .B(new_n1089), .C1(G294), .C2(new_n829), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1176), .B(new_n1177), .C1(new_n823), .C2(new_n875), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n1168), .A2(new_n1174), .B1(new_n1175), .B2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1162), .B1(new_n1179), .B2(new_n783), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1159), .A2(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT120), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n767), .B2(new_n1156), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1158), .A2(new_n1183), .ZN(G378));
  INV_X1    g0984(.A(KEYINPUT123), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n934), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n943), .A2(KEYINPUT40), .A3(new_n1114), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n940), .B1(new_n922), .B2(new_n924), .ZN(new_n1188));
  OAI211_X1 g0988(.A(G330), .B(new_n1187), .C1(new_n1188), .C2(KEYINPUT40), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n302), .A2(new_n306), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n267), .A2(new_n884), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n302), .B(new_n306), .C1(new_n267), .C2(new_n884), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1194), .B(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1189), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1197), .B1(new_n947), .B2(G330), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1186), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1189), .A2(new_n1198), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n947), .A2(G330), .A3(new_n1197), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1202), .A2(new_n1203), .A3(new_n934), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n766), .B1(new_n1201), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1198), .A2(new_n780), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n768), .B1(G50), .B2(new_n1160), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n799), .A2(G132), .B1(new_n1063), .B2(G137), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT122), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n796), .A2(G128), .B1(G150), .B2(new_n864), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n812), .A2(G125), .B1(new_n806), .B2(new_n1164), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1209), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n1214), .A2(KEYINPUT59), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(KEYINPUT59), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n789), .A2(G159), .ZN(new_n1217));
  AOI211_X1 g1017(.A(G33), .B(G41), .C1(new_n829), .C2(G124), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n796), .A2(G107), .B1(G116), .B2(new_n812), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n958), .B2(new_n788), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n802), .A2(new_n242), .B1(new_n808), .B2(new_n823), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n832), .A2(new_n620), .B1(new_n815), .B2(new_n320), .ZN(new_n1223));
  NOR3_X1   g1023(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n338), .B(new_n592), .C1(new_n319), .C2(new_n805), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT121), .ZN(new_n1226));
  OR2_X1    g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1224), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT58), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n338), .A2(new_n592), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1233), .B(new_n240), .C1(G33), .C2(G41), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1219), .A2(new_n1231), .A3(new_n1232), .A4(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1207), .B1(new_n1235), .B2(new_n783), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1206), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1185), .B1(new_n1205), .B2(new_n1238), .ZN(new_n1239));
  AND3_X1   g1039(.A1(new_n1202), .A2(new_n1203), .A3(new_n934), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n934), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n767), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1242), .A2(KEYINPUT123), .A3(new_n1237), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1239), .A2(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1132), .B1(new_n1153), .B2(new_n1157), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(KEYINPUT57), .B1(new_n1245), .B2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(KEYINPUT118), .B1(new_n1130), .B2(new_n1140), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1156), .A2(new_n1142), .A3(new_n1152), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1143), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(KEYINPUT57), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n763), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1244), .B1(new_n1248), .B2(new_n1253), .ZN(G375));
  NOR3_X1   g1054(.A1(new_n1136), .A2(new_n1132), .A3(new_n1139), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(new_n1255), .A2(new_n1152), .A3(new_n1019), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n1256), .B(KEYINPUT124), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n853), .B1(new_n242), .B2(new_n879), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n783), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n871), .A2(new_n622), .B1(new_n485), .B2(new_n818), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(G77), .B2(new_n861), .ZN(new_n1261));
  OAI221_X1 g1061(.A(new_n289), .B1(new_n808), .B2(new_n613), .C1(new_n320), .C2(new_n802), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n795), .A2(new_n823), .B1(new_n620), .B2(new_n805), .ZN(new_n1263));
  AOI211_X1 g1063(.A(new_n1262), .B(new_n1263), .C1(G294), .C2(new_n812), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n973), .A2(new_n1164), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n812), .A2(G132), .B1(G50), .B2(new_n864), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n796), .A2(G137), .B1(G159), .B2(new_n806), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n338), .B1(G128), .B2(new_n829), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1063), .A2(G150), .B1(new_n789), .B2(G58), .ZN(new_n1269));
  AND4_X1   g1069(.A1(new_n1266), .A2(new_n1267), .A3(new_n1268), .A4(new_n1269), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n1261), .A2(new_n1264), .B1(new_n1265), .B2(new_n1270), .ZN(new_n1271));
  OAI221_X1 g1071(.A(new_n1258), .B1(new_n1259), .B2(new_n1271), .C1(new_n1127), .C2(new_n781), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n1147), .A2(new_n1148), .B1(new_n1150), .B2(new_n1138), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1272), .B1(new_n1273), .B2(new_n766), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1257), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(G381));
  XNOR2_X1  g1076(.A(G375), .B(KEYINPUT125), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1082), .A2(new_n841), .A3(new_n1084), .ZN(new_n1278));
  NOR3_X1   g1078(.A1(G390), .A2(G384), .A3(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(G378), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n1279), .A2(new_n1041), .A3(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1277), .A2(new_n1281), .A3(new_n1275), .ZN(G407));
  INV_X1    g1082(.A(G213), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1283), .A2(G343), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1277), .A2(new_n1280), .A3(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(G407), .A2(new_n1285), .A3(G213), .ZN(G409));
  NAND2_X1  g1086(.A1(G393), .A2(G396), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(G390), .A2(new_n1278), .A3(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1278), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1289), .A2(new_n1107), .A3(new_n1110), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n1041), .A2(new_n1288), .A3(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1041), .B1(new_n1290), .B2(new_n1288), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  AND2_X1   g1094(.A1(new_n1284), .A2(G2897), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT127), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n854), .A2(KEYINPUT126), .A3(new_n881), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1298), .B(new_n1272), .C1(new_n1273), .C2(new_n766), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1255), .A2(KEYINPUT60), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1273), .A2(KEYINPUT60), .A3(new_n1143), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1302), .A2(new_n1140), .A3(new_n763), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1300), .B1(new_n1301), .B2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT126), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(G384), .A2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1304), .A2(new_n1307), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1300), .B(new_n1306), .C1(new_n1301), .C2(new_n1303), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1297), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  AOI211_X1 g1112(.A(new_n1296), .B(new_n1295), .C1(new_n1308), .C2(new_n1309), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1245), .A2(new_n1247), .A3(new_n1020), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1205), .A2(new_n1238), .ZN(new_n1316));
  AOI21_X1  g1116(.A(G378), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT57), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1318), .B1(new_n1201), .B2(new_n1204), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n715), .B1(new_n1245), .B2(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1318), .B1(new_n1251), .B2(new_n1246), .ZN(new_n1321));
  AOI22_X1  g1121(.A1(new_n1320), .A2(new_n1321), .B1(new_n1239), .B2(new_n1243), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1317), .B1(new_n1322), .B2(G378), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1314), .B1(new_n1323), .B2(new_n1284), .ZN(new_n1324));
  OAI211_X1 g1124(.A(new_n1244), .B(G378), .C1(new_n1248), .C2(new_n1253), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(new_n1280), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1325), .A2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT62), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1284), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1328), .A2(new_n1329), .A3(new_n1330), .A4(new_n1310), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT61), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1324), .A2(new_n1331), .A3(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1284), .B1(new_n1325), .B2(new_n1327), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1329), .B1(new_n1334), .B2(new_n1310), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1294), .B1(new_n1333), .B2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT63), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1328), .A2(new_n1330), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1310), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1337), .B1(new_n1338), .B2(new_n1339), .ZN(new_n1340));
  AOI21_X1  g1140(.A(KEYINPUT61), .B1(new_n1338), .B2(new_n1314), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1334), .A2(KEYINPUT63), .A3(new_n1310), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1340), .A2(new_n1341), .A3(new_n1293), .A4(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1336), .A2(new_n1343), .ZN(G405));
  NAND2_X1  g1144(.A1(G375), .A2(new_n1280), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1345), .A2(new_n1325), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1346), .A2(new_n1339), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1345), .A2(new_n1325), .A3(new_n1310), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1349));
  XNOR2_X1  g1149(.A(new_n1349), .B(new_n1293), .ZN(G402));
endmodule


