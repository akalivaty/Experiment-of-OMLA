//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 1 1 1 1 0 1 1 0 1 0 0 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n449, new_n450, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n571, new_n572, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n623,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1200, new_n1201, new_n1202;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT66), .B(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT67), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  INV_X1    g023(.A(G567), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT68), .Z(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g027(.A1(G219), .A2(G218), .A3(G220), .A4(G221), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n454), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2106), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n455), .A2(new_n449), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND3_X1   g038(.A1(KEYINPUT69), .A2(G113), .A3(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(KEYINPUT69), .B1(G113), .B2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(G125), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n463), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  OAI211_X1 g045(.A(G137), .B(new_n463), .C1(new_n467), .C2(new_n468), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n463), .A2(G101), .A3(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n470), .A2(new_n473), .ZN(G160));
  OAI21_X1  g049(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(G112), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n475), .B1(new_n476), .B2(G2105), .ZN(new_n477));
  OR2_X1    g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n463), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT70), .ZN(new_n482));
  AOI21_X1  g057(.A(G2105), .B1(new_n478), .B2(new_n479), .ZN(new_n483));
  AOI211_X1 g058(.A(new_n477), .B(new_n482), .C1(G136), .C2(new_n483), .ZN(G162));
  OAI211_X1 g059(.A(G126), .B(G2105), .C1(new_n467), .C2(new_n468), .ZN(new_n485));
  OR2_X1    g060(.A1(G102), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G114), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n486), .A2(new_n488), .A3(G2104), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n492), .B1(new_n467), .B2(new_n468), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n492), .B(new_n495), .C1(new_n468), .C2(new_n467), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n490), .B1(new_n494), .B2(new_n496), .ZN(G164));
  INV_X1    g072(.A(G50), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT6), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n499), .B1(new_n500), .B2(G651), .ZN(new_n501));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(KEYINPUT71), .A3(KEYINPUT6), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n500), .A2(G651), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n504), .A2(G543), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n504), .A2(new_n511), .A3(new_n505), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n498), .A2(new_n506), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT72), .ZN(new_n516));
  OR3_X1    g091(.A1(new_n515), .A2(new_n516), .A3(new_n502), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n515), .B2(new_n502), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n514), .B1(new_n517), .B2(new_n518), .ZN(G166));
  AND2_X1   g094(.A1(G63), .A2(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT7), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT7), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n523), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n511), .A2(new_n520), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G51), .ZN(new_n526));
  INV_X1    g101(.A(G89), .ZN(new_n527));
  OAI221_X1 g102(.A(new_n525), .B1(new_n506), .B2(new_n526), .C1(new_n527), .C2(new_n512), .ZN(G286));
  INV_X1    g103(.A(G286), .ZN(G168));
  AOI22_X1  g104(.A1(new_n501), .A2(new_n503), .B1(new_n500), .B2(G651), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n530), .A2(G52), .A3(G543), .ZN(new_n531));
  INV_X1    g106(.A(G64), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n532), .B1(new_n509), .B2(new_n510), .ZN(new_n533));
  AND2_X1   g108(.A1(G77), .A2(G543), .ZN(new_n534));
  OAI21_X1  g109(.A(G651), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(G90), .ZN(new_n536));
  OAI211_X1 g111(.A(new_n531), .B(new_n535), .C1(new_n536), .C2(new_n512), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT73), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n537), .B(new_n538), .ZN(G171));
  INV_X1    g114(.A(G43), .ZN(new_n540));
  INV_X1    g115(.A(G81), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n540), .A2(new_n506), .B1(new_n512), .B2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n544), .B1(new_n509), .B2(new_n510), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT74), .ZN(new_n546));
  AND2_X1   g121(.A1(G68), .A2(G543), .ZN(new_n547));
  OR3_X1    g122(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n546), .B1(new_n545), .B2(new_n547), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n548), .A2(G651), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n543), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  INV_X1    g132(.A(G53), .ZN(new_n558));
  OAI21_X1  g133(.A(KEYINPUT9), .B1(new_n506), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n530), .A2(new_n560), .A3(G53), .A4(G543), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n530), .A2(G91), .A3(new_n511), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n564), .B1(new_n509), .B2(new_n510), .ZN(new_n565));
  AND2_X1   g140(.A1(G78), .A2(G543), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AND2_X1   g142(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n562), .A2(new_n568), .ZN(G299));
  XNOR2_X1  g144(.A(new_n537), .B(KEYINPUT73), .ZN(G301));
  NAND2_X1  g145(.A1(new_n517), .A2(new_n518), .ZN(new_n571));
  INV_X1    g146(.A(new_n514), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(G303));
  INV_X1    g148(.A(G87), .ZN(new_n574));
  OAI21_X1  g149(.A(KEYINPUT75), .B1(new_n512), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT75), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n530), .A2(new_n576), .A3(G87), .A4(new_n511), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n510), .ZN(new_n579));
  NOR2_X1   g154(.A1(KEYINPUT5), .A2(G543), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(G74), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n502), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n506), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n583), .B1(new_n584), .B2(G49), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n578), .A2(new_n585), .ZN(G288));
  INV_X1    g161(.A(G48), .ZN(new_n587));
  INV_X1    g162(.A(G86), .ZN(new_n588));
  OAI22_X1  g163(.A1(new_n587), .A2(new_n506), .B1(new_n512), .B2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(G61), .ZN(new_n591));
  OAI21_X1  g166(.A(KEYINPUT76), .B1(new_n581), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT76), .ZN(new_n593));
  OAI211_X1 g168(.A(new_n593), .B(G61), .C1(new_n579), .C2(new_n580), .ZN(new_n594));
  NAND2_X1  g169(.A1(G73), .A2(G543), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT77), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n592), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(KEYINPUT78), .B1(new_n597), .B2(G651), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n596), .A2(new_n594), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n593), .B1(new_n511), .B2(G61), .ZN(new_n600));
  OAI211_X1 g175(.A(KEYINPUT78), .B(G651), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n590), .B1(new_n598), .B2(new_n602), .ZN(G305));
  NAND2_X1  g178(.A1(new_n584), .A2(G47), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n605));
  XNOR2_X1  g180(.A(KEYINPUT79), .B(G85), .ZN(new_n606));
  OAI221_X1 g181(.A(new_n604), .B1(new_n502), .B2(new_n605), .C1(new_n512), .C2(new_n606), .ZN(G290));
  NAND2_X1  g182(.A1(new_n584), .A2(KEYINPUT80), .ZN(new_n608));
  INV_X1    g183(.A(G54), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT80), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n609), .B1(new_n506), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n581), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n608), .A2(new_n611), .B1(G651), .B2(new_n614), .ZN(new_n615));
  NAND4_X1  g190(.A1(new_n504), .A2(G92), .A3(new_n511), .A4(new_n505), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT10), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  MUX2_X1   g194(.A(new_n619), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g195(.A(new_n619), .B(G301), .S(G868), .Z(G321));
  NAND2_X1  g196(.A1(G286), .A2(G868), .ZN(new_n622));
  INV_X1    g197(.A(G299), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G868), .ZN(G297));
  OAI21_X1  g199(.A(new_n622), .B1(new_n623), .B2(G868), .ZN(G280));
  INV_X1    g200(.A(new_n619), .ZN(new_n626));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(G860), .ZN(G148));
  INV_X1    g203(.A(G868), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n551), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n619), .A2(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(new_n629), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g208(.A1(new_n483), .A2(G135), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n480), .A2(G123), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n463), .A2(G111), .ZN(new_n636));
  OAI21_X1  g211(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n634), .B(new_n635), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(G2096), .Z(new_n639));
  NAND3_X1  g214(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT12), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT13), .ZN(new_n642));
  INV_X1    g217(.A(G2100), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n639), .A2(new_n644), .A3(new_n645), .ZN(G156));
  INV_X1    g221(.A(KEYINPUT14), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2427), .B(G2438), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2430), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT15), .B(G2435), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n647), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n651), .B1(new_n650), .B2(new_n649), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2451), .B(G2454), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1341), .B(G1348), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n652), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2443), .B(G2446), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n659), .A2(new_n660), .A3(G14), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT81), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(G401));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT82), .Z(new_n667));
  NOR2_X1   g242(.A1(G2072), .A2(G2078), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n442), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n665), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(KEYINPUT17), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n670), .B1(new_n667), .B2(new_n671), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n665), .B(new_n666), .C1(new_n442), .C2(new_n668), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT18), .Z(new_n674));
  NAND3_X1  g249(.A1(new_n667), .A2(new_n671), .A3(new_n665), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n672), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2096), .B(G2100), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G227));
  XNOR2_X1  g253(.A(G1956), .B(G2474), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1961), .B(G1966), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G1971), .B(G1976), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n679), .A2(new_n680), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n681), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n683), .A2(KEYINPUT83), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n683), .A2(new_n684), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT20), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1981), .B(G1986), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT84), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n693), .A2(new_n695), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1991), .B(G1996), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n696), .A2(new_n699), .A3(new_n697), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(G229));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n705), .A2(G23), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G288), .B2(G16), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT85), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT33), .B(G1976), .Z(new_n709));
  OR2_X1    g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n705), .A2(G22), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G166), .B2(new_n705), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(G1971), .Z(new_n713));
  NAND2_X1  g288(.A1(new_n708), .A2(new_n709), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n705), .A2(G6), .ZN(new_n715));
  OAI21_X1  g290(.A(G651), .B1(new_n599), .B2(new_n600), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT78), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n589), .B1(new_n718), .B2(new_n601), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n715), .B1(new_n719), .B2(new_n705), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT32), .B(G1981), .Z(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND4_X1  g297(.A1(new_n710), .A2(new_n713), .A3(new_n714), .A4(new_n722), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n723), .A2(KEYINPUT34), .ZN(new_n724));
  OR2_X1    g299(.A1(G16), .A2(G24), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G290), .B2(new_n705), .ZN(new_n726));
  INV_X1    g301(.A(G1986), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n726), .A2(new_n727), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n483), .A2(G131), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n480), .A2(G119), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n463), .A2(G107), .ZN(new_n732));
  OAI21_X1  g307(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n730), .B(new_n731), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  MUX2_X1   g309(.A(G25), .B(new_n734), .S(G29), .Z(new_n735));
  XOR2_X1   g310(.A(KEYINPUT35), .B(G1991), .Z(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n735), .B(new_n737), .ZN(new_n738));
  OR4_X1    g313(.A1(KEYINPUT86), .A2(new_n728), .A3(new_n729), .A4(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n723), .B2(KEYINPUT34), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n724), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT87), .B(KEYINPUT36), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n742), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n724), .A2(new_n740), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(G5), .A2(G16), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT101), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G171), .B2(G16), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT102), .ZN(new_n750));
  INV_X1    g325(.A(G1961), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(G29), .A2(G33), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT89), .Z(new_n754));
  NAND2_X1  g329(.A1(new_n483), .A2(G139), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT90), .Z(new_n756));
  NAND3_X1  g331(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT25), .Z(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT3), .B(G2104), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n759), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n756), .B(new_n758), .C1(new_n463), .C2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G29), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n754), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT91), .Z(new_n764));
  AND2_X1   g339(.A1(new_n764), .A2(G2072), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n764), .A2(G2072), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT97), .B(KEYINPUT26), .Z(new_n767));
  NAND3_X1  g342(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n463), .A2(G105), .A3(G2104), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT96), .Z(new_n771));
  NAND2_X1  g346(.A1(new_n480), .A2(G129), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n769), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n483), .A2(G141), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT95), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n776), .A2(new_n762), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n762), .B2(G32), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT27), .B(G1996), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT98), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n762), .A2(G26), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT28), .Z(new_n784));
  OAI21_X1  g359(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n785));
  INV_X1    g360(.A(G116), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n785), .B1(new_n786), .B2(G2105), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT88), .ZN(new_n788));
  AOI22_X1  g363(.A1(G128), .A2(new_n480), .B1(new_n483), .B2(G140), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n784), .B1(new_n790), .B2(G29), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G2067), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT92), .B(KEYINPUT24), .Z(new_n793));
  INV_X1    g368(.A(G34), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n762), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n794), .B2(new_n793), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT93), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G29), .B2(G160), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(G2084), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT94), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n792), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NOR4_X1   g376(.A1(new_n765), .A2(new_n766), .A3(new_n782), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(G162), .A2(G29), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G29), .B2(G35), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT29), .B(G2090), .Z(new_n805));
  OR2_X1    g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n778), .A2(new_n781), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n804), .A2(new_n805), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n799), .A2(new_n800), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n806), .A2(new_n807), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n705), .A2(G21), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G168), .B2(new_n705), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n812), .A2(G1966), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n552), .A2(G16), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(G16), .B2(G19), .ZN(new_n815));
  INV_X1    g390(.A(G1341), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n813), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(new_n816), .B2(new_n815), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n798), .A2(G2084), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n812), .A2(G1966), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT99), .B(KEYINPUT31), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(G11), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT30), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n762), .B1(new_n823), .B2(G28), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n824), .A2(KEYINPUT100), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(G28), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n824), .B2(KEYINPUT100), .ZN(new_n827));
  OAI221_X1 g402(.A(new_n822), .B1(new_n825), .B2(new_n827), .C1(new_n638), .C2(new_n762), .ZN(new_n828));
  NAND2_X1  g403(.A1(G164), .A2(G29), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(G27), .B2(G29), .ZN(new_n830));
  INV_X1    g405(.A(G2078), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n828), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n830), .A2(new_n831), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n819), .A2(new_n820), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  NOR3_X1   g409(.A1(new_n810), .A2(new_n818), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n626), .A2(G16), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(G4), .B2(G16), .ZN(new_n837));
  INV_X1    g412(.A(G1348), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n837), .A2(new_n838), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n705), .A2(G20), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT23), .Z(new_n842));
  AOI21_X1  g417(.A(new_n842), .B1(G299), .B2(G16), .ZN(new_n843));
  INV_X1    g418(.A(G1956), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NOR3_X1   g420(.A1(new_n839), .A2(new_n840), .A3(new_n845), .ZN(new_n846));
  AND3_X1   g421(.A1(new_n802), .A2(new_n835), .A3(new_n846), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n746), .A2(new_n752), .A3(new_n847), .ZN(G150));
  INV_X1    g423(.A(G150), .ZN(G311));
  NAND2_X1  g424(.A1(new_n626), .A2(G559), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT38), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n530), .A2(G93), .A3(new_n511), .ZN(new_n852));
  AOI22_X1  g427(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n853));
  INV_X1    g428(.A(G55), .ZN(new_n854));
  OAI221_X1 g429(.A(new_n852), .B1(new_n853), .B2(new_n502), .C1(new_n854), .C2(new_n506), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n551), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n506), .A2(new_n854), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n853), .A2(new_n502), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n543), .A2(new_n859), .A3(new_n550), .A4(new_n852), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n851), .B(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT39), .ZN(new_n863));
  AOI21_X1  g438(.A(G860), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(new_n863), .B2(new_n862), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n855), .A2(G860), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n866), .B(KEYINPUT37), .Z(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(G145));
  XNOR2_X1  g443(.A(new_n638), .B(G160), .ZN(new_n869));
  XNOR2_X1  g444(.A(G162), .B(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n496), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n495), .B1(new_n759), .B2(new_n492), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n485), .B(new_n489), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n790), .B(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n480), .A2(G130), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n463), .A2(G118), .ZN(new_n876));
  OAI21_X1  g451(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n877));
  AND3_X1   g452(.A1(new_n483), .A2(KEYINPUT104), .A3(G142), .ZN(new_n878));
  AOI21_X1  g453(.A(KEYINPUT104), .B1(new_n483), .B2(G142), .ZN(new_n879));
  OAI221_X1 g454(.A(new_n875), .B1(new_n876), .B2(new_n877), .C1(new_n878), .C2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n874), .B(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n761), .A2(KEYINPUT103), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n776), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n883), .A2(new_n776), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n734), .B(new_n641), .ZN(new_n887));
  NOR3_X1   g462(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n887), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n761), .A2(KEYINPUT103), .ZN(new_n890));
  INV_X1    g465(.A(new_n776), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n889), .B1(new_n892), .B2(new_n884), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n882), .B1(new_n888), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n887), .B1(new_n885), .B2(new_n886), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n892), .A2(new_n884), .A3(new_n889), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n895), .A2(new_n881), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n870), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n898), .A2(G37), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n894), .A2(new_n897), .A3(new_n870), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n900), .A2(KEYINPUT105), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n900), .A2(KEYINPUT105), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n899), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  XOR2_X1   g478(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n904));
  XNOR2_X1  g479(.A(new_n903), .B(new_n904), .ZN(G395));
  XNOR2_X1  g480(.A(new_n719), .B(G166), .ZN(new_n906));
  XNOR2_X1  g481(.A(G290), .B(G288), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n906), .B(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT42), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n861), .A2(new_n631), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n861), .A2(new_n631), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n619), .A2(G299), .ZN(new_n913));
  AOI22_X1  g488(.A1(new_n615), .A2(new_n618), .B1(new_n562), .B2(new_n568), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n912), .A2(KEYINPUT107), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n623), .A2(new_n618), .A3(new_n615), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n619), .A2(G299), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT41), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(KEYINPUT41), .B1(new_n913), .B2(new_n914), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n912), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n910), .A2(new_n911), .A3(new_n915), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT107), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n916), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT108), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n928), .B(new_n916), .C1(new_n922), .C2(new_n925), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n909), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n929), .A2(new_n909), .ZN(new_n931));
  OAI21_X1  g506(.A(G868), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n855), .A2(new_n629), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(G295));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n933), .ZN(G331));
  NAND2_X1  g510(.A1(new_n921), .A2(new_n920), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n551), .A2(new_n855), .ZN(new_n937));
  AOI22_X1  g512(.A1(new_n543), .A2(new_n550), .B1(new_n859), .B2(new_n852), .ZN(new_n938));
  OAI21_X1  g513(.A(G301), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(G171), .A2(new_n856), .A3(new_n860), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n939), .A2(new_n940), .A3(G168), .ZN(new_n941));
  AOI21_X1  g516(.A(G168), .B1(new_n939), .B2(new_n940), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n936), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n939), .A2(new_n940), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(G286), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n939), .A2(new_n940), .A3(G168), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n945), .A2(new_n915), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n943), .A2(new_n947), .A3(new_n908), .ZN(new_n948));
  INV_X1    g523(.A(G37), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n908), .B1(new_n943), .B2(new_n947), .ZN(new_n951));
  OAI21_X1  g526(.A(KEYINPUT43), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT109), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n921), .A2(new_n920), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n915), .A2(KEYINPUT109), .A3(new_n919), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n954), .B(new_n955), .C1(new_n941), .C2(new_n942), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n947), .ZN(new_n957));
  INV_X1    g532(.A(new_n908), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n959), .A2(new_n960), .A3(new_n949), .A4(new_n948), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n952), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  OR3_X1    g538(.A1(new_n950), .A2(KEYINPUT43), .A3(new_n951), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT110), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n908), .B1(new_n956), .B2(new_n947), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n965), .B1(new_n950), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n950), .A2(new_n965), .A3(new_n966), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n964), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n963), .B1(new_n970), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g546(.A(G1384), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n873), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT111), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT45), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT112), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n976), .B1(G160), .B2(G40), .ZN(new_n977));
  INV_X1    g552(.A(G125), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n978), .B1(new_n478), .B2(new_n479), .ZN(new_n979));
  NAND2_X1  g554(.A1(G113), .A2(G2104), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT69), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(KEYINPUT69), .A2(G113), .A3(G2104), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(G2105), .B1(new_n979), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n472), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n986), .B1(new_n483), .B2(G137), .ZN(new_n987));
  AND4_X1   g562(.A1(new_n976), .A2(new_n985), .A3(new_n987), .A4(G40), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n977), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(G164), .A2(G1384), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT111), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n975), .A2(new_n989), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n790), .A2(G2067), .ZN(new_n994));
  INV_X1    g569(.A(G2067), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n788), .A2(new_n995), .A3(new_n789), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1996), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n776), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n993), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n992), .A2(G1996), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n1002), .A2(KEYINPUT113), .A3(new_n891), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT113), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1004), .B1(new_n1001), .B2(new_n776), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1000), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT114), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  OAI211_X1 g583(.A(KEYINPUT114), .B(new_n1000), .C1(new_n1003), .C2(new_n1005), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n734), .B(new_n736), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1008), .B(new_n1009), .C1(new_n992), .C2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(G290), .B(G1986), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1011), .B1(new_n993), .B2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(KEYINPUT119), .B(KEYINPUT63), .ZN(new_n1014));
  XNOR2_X1  g589(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n1015));
  NAND3_X1  g590(.A1(G303), .A2(G8), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1015), .ZN(new_n1017));
  INV_X1    g592(.A(G8), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1017), .B1(G166), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n871), .A2(new_n872), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1023), .B(new_n972), .C1(new_n1024), .C2(new_n490), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n985), .A2(new_n987), .A3(G40), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT112), .ZN(new_n1027));
  NAND3_X1  g602(.A1(G160), .A2(new_n976), .A3(G40), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1022), .A2(new_n1025), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G2090), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT45), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1032), .B1(G164), .B2(G1384), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n873), .A2(KEYINPUT45), .A3(new_n972), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1033), .A2(new_n1034), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1035));
  XOR2_X1   g610(.A(KEYINPUT115), .B(G1971), .Z(new_n1036));
  AOI22_X1  g611(.A1(new_n1030), .A2(new_n1031), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1021), .B1(new_n1037), .B2(new_n1018), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n990), .A2(new_n1028), .A3(new_n1027), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n578), .A2(new_n585), .A3(G1976), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1039), .A2(G8), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT52), .ZN(new_n1042));
  XNOR2_X1  g617(.A(KEYINPUT117), .B(G1976), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT52), .B1(G288), .B2(new_n1043), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1044), .A2(G8), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1042), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1039), .A2(G8), .ZN(new_n1048));
  INV_X1    g623(.A(G1981), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1049), .B(new_n590), .C1(new_n598), .C2(new_n602), .ZN(new_n1050));
  INV_X1    g625(.A(new_n716), .ZN(new_n1051));
  OAI21_X1  g626(.A(G1981), .B1(new_n1051), .B2(new_n589), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT49), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1048), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1050), .A2(KEYINPUT49), .A3(new_n1052), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1029), .A2(G2090), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1020), .B(G8), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1038), .A2(new_n1047), .A3(new_n1057), .A4(new_n1060), .ZN(new_n1061));
  XOR2_X1   g636(.A(KEYINPUT118), .B(G2084), .Z(new_n1062));
  INV_X1    g637(.A(G1966), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1030), .A2(new_n1062), .B1(new_n1035), .B2(new_n1063), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n1064), .A2(new_n1018), .A3(G286), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1014), .B1(new_n1061), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT120), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT121), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1046), .B1(new_n1056), .B2(new_n1055), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1070), .A2(new_n1060), .A3(new_n1038), .A4(new_n1065), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT63), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1069), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1061), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1074), .A2(KEYINPUT121), .A3(KEYINPUT63), .A4(new_n1065), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1071), .A2(new_n1076), .A3(new_n1014), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1068), .A2(new_n1073), .A3(new_n1075), .A4(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1070), .ZN(new_n1079));
  NOR2_X1   g654(.A1(G288), .A2(G1976), .ZN(new_n1080));
  AOI22_X1  g655(.A1(new_n1057), .A2(new_n1080), .B1(new_n1049), .B2(new_n719), .ZN(new_n1081));
  OAI22_X1  g656(.A1(new_n1079), .A2(new_n1060), .B1(new_n1081), .B2(new_n1048), .ZN(new_n1082));
  NAND2_X1  g657(.A1(G286), .A2(G8), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT125), .ZN(new_n1084));
  XNOR2_X1  g659(.A(new_n1083), .B(new_n1084), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1086));
  AOI21_X1  g661(.A(G1966), .B1(new_n1086), .B2(new_n989), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1062), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1029), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1085), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n989), .A2(new_n1022), .A3(new_n1025), .A4(new_n1062), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1035), .A2(new_n1063), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1018), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1090), .B(KEYINPUT51), .C1(new_n1085), .C2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1085), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT51), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1095), .B(new_n1096), .C1(new_n1064), .C2(new_n1018), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1094), .A2(KEYINPUT62), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(KEYINPUT62), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1101), .B1(new_n1035), .B2(G2078), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1101), .A2(G2078), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1086), .A2(new_n989), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1029), .A2(new_n751), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1102), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(G171), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1061), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1082), .B1(new_n1100), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1078), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT127), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT126), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1029), .A2(new_n1112), .A3(new_n751), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1112), .B1(new_n1029), .B2(new_n751), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n989), .A2(new_n831), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n975), .A2(new_n991), .ZN(new_n1117));
  AND4_X1   g692(.A1(G40), .A2(new_n1034), .A3(G160), .A4(new_n1103), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1116), .A2(new_n1101), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(G301), .B1(new_n1115), .B2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1102), .A2(new_n1104), .A3(G301), .A4(new_n1105), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(KEYINPUT54), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1111), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1105), .A2(KEYINPUT126), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1029), .A2(new_n1112), .A3(new_n751), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1124), .A2(new_n1125), .A3(new_n1102), .A4(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(G171), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1128), .A2(KEYINPUT127), .A3(KEYINPUT54), .A4(new_n1121), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1123), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1115), .A2(G301), .A3(new_n1119), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT54), .B1(new_n1131), .B2(new_n1107), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1090), .A2(KEYINPUT51), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1085), .B1(new_n1134), .B2(G8), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1097), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1132), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1130), .A2(new_n1137), .A3(new_n1074), .ZN(new_n1138));
  XNOR2_X1  g713(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n1139));
  XNOR2_X1  g714(.A(KEYINPUT56), .B(G2072), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n989), .A2(new_n1033), .A3(new_n1034), .A4(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1029), .A2(new_n844), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT57), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n562), .A2(new_n1143), .A3(new_n568), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1143), .B1(new_n562), .B2(new_n568), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1141), .A2(new_n1142), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(KEYINPUT122), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT122), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1141), .A2(new_n1142), .A3(new_n1146), .A4(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1146), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1139), .B1(new_n1151), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1035), .ZN(new_n1156));
  AOI22_X1  g731(.A1(new_n1156), .A2(new_n1140), .B1(new_n844), .B2(new_n1029), .ZN(new_n1157));
  OAI21_X1  g732(.A(KEYINPUT61), .B1(new_n1157), .B2(new_n1146), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1147), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1039), .ZN(new_n1160));
  XNOR2_X1  g735(.A(KEYINPUT58), .B(G1341), .ZN(new_n1161));
  OAI22_X1  g736(.A1(new_n1160), .A2(new_n1161), .B1(new_n1035), .B2(G1996), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT59), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1162), .A2(new_n1163), .A3(new_n552), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1163), .B1(new_n1162), .B2(new_n552), .ZN(new_n1165));
  OAI22_X1  g740(.A1(new_n1158), .A2(new_n1159), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(KEYINPUT124), .B1(new_n1155), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1162), .A2(new_n552), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1162), .A2(new_n1163), .A3(new_n552), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1171), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1172));
  AOI22_X1  g747(.A1(new_n1169), .A2(new_n1170), .B1(new_n1172), .B2(new_n1147), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT124), .ZN(new_n1174));
  AOI22_X1  g749(.A1(new_n1148), .A2(new_n1150), .B1(new_n1153), .B2(new_n1152), .ZN(new_n1175));
  OAI211_X1 g750(.A(new_n1173), .B(new_n1174), .C1(new_n1175), .C2(new_n1139), .ZN(new_n1176));
  AOI22_X1  g751(.A1(new_n1160), .A2(new_n995), .B1(new_n1029), .B2(new_n838), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(KEYINPUT60), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1178), .B(new_n626), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1179), .B1(KEYINPUT60), .B2(new_n1177), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1167), .A2(new_n1176), .A3(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1154), .B1(new_n619), .B2(new_n1177), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(new_n1151), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1138), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1013), .B1(new_n1110), .B2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n993), .B1(new_n891), .B2(new_n997), .ZN(new_n1186));
  AND2_X1   g761(.A1(new_n1002), .A2(KEYINPUT46), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1002), .A2(KEYINPUT46), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1186), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n1189), .B(KEYINPUT47), .ZN(new_n1190));
  NOR3_X1   g765(.A1(new_n992), .A2(G1986), .A3(G290), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n1191), .B(KEYINPUT48), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1190), .B1(new_n1011), .B2(new_n1192), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n734), .A2(new_n737), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1008), .A2(new_n1009), .A3(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n992), .B1(new_n1195), .B2(new_n996), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1193), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1185), .A2(new_n1197), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g773(.A1(G227), .A2(new_n461), .ZN(new_n1200));
  AND4_X1   g774(.A1(new_n663), .A2(new_n701), .A3(new_n702), .A4(new_n1200), .ZN(new_n1201));
  NAND2_X1  g775(.A1(new_n952), .A2(new_n961), .ZN(new_n1202));
  NAND3_X1  g776(.A1(new_n1201), .A2(new_n903), .A3(new_n1202), .ZN(G225));
  INV_X1    g777(.A(G225), .ZN(G308));
endmodule


