//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 1 1 1 0 0 0 0 0 1 0 1 0 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1331, new_n1332, new_n1333;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n206));
  INV_X1    g0006(.A(G68), .ZN(new_n207));
  INV_X1    g0007(.A(G238), .ZN(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n206), .B1(new_n207), .B2(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(G58), .ZN(new_n213));
  INV_X1    g0013(.A(G232), .ZN(new_n214));
  INV_X1    g0014(.A(G97), .ZN(new_n215));
  INV_X1    g0015(.A(G257), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n205), .B1(new_n211), .B2(new_n217), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  OR2_X1    g0019(.A1(new_n202), .A2(KEYINPUT64), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n202), .A2(KEYINPUT64), .ZN(new_n221));
  AND3_X1   g0021(.A1(new_n220), .A2(G50), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n205), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT0), .ZN(new_n229));
  NAND3_X1  g0029(.A1(new_n219), .A2(new_n226), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n218), .ZN(G361));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT65), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT66), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n236), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n242), .B(new_n243), .Z(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  INV_X1    g0048(.A(G1), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G274), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT67), .B(G45), .ZN(new_n251));
  INV_X1    g0051(.A(G41), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G226), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G1698), .ZN(new_n255));
  AND2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  OAI221_X1 g0057(.A(new_n255), .B1(G223), .B2(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G87), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT73), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n259), .B(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n223), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G41), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n253), .B1(new_n262), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n264), .A2(KEYINPUT68), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT68), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(G33), .A3(G41), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n268), .A2(new_n270), .A3(new_n263), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n249), .B1(G41), .B2(G45), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G232), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n267), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G200), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n256), .A2(new_n257), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT72), .B(KEYINPUT7), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(new_n278), .A3(new_n224), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT3), .ZN(new_n280));
  INV_X1    g0080(.A(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(new_n224), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT7), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n279), .A2(new_n285), .A3(G68), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G159), .ZN(new_n288));
  AND2_X1   g0088(.A1(G58), .A2(G68), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(new_n201), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n288), .B1(new_n290), .B2(new_n224), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n286), .A2(KEYINPUT16), .A3(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n223), .B1(new_n205), .B2(new_n281), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n284), .A2(new_n278), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n282), .A2(KEYINPUT7), .A3(new_n224), .A4(new_n283), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n291), .B1(new_n297), .B2(G68), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n293), .B(new_n294), .C1(new_n298), .C2(KEYINPUT16), .ZN(new_n299));
  XOR2_X1   g0099(.A(KEYINPUT8), .B(G58), .Z(new_n300));
  INV_X1    g0100(.A(KEYINPUT69), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n301), .B1(new_n224), .B2(G1), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n249), .A2(KEYINPUT69), .A3(G20), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AND2_X1   g0104(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n249), .A2(G13), .A3(G20), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n306), .B(new_n223), .C1(new_n281), .C2(new_n205), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n306), .ZN(new_n309));
  INV_X1    g0109(.A(new_n300), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n305), .A2(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n267), .A2(G190), .A3(new_n274), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n276), .A2(new_n299), .A3(new_n311), .A4(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT17), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n299), .A2(new_n311), .ZN(new_n316));
  INV_X1    g0116(.A(G169), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n317), .B1(new_n267), .B2(new_n274), .ZN(new_n318));
  AND3_X1   g0118(.A1(new_n267), .A2(G179), .A3(new_n274), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n316), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(KEYINPUT18), .ZN(new_n321));
  INV_X1    g0121(.A(new_n318), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n267), .A2(G179), .A3(new_n274), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n322), .A2(new_n323), .B1(new_n299), .B2(new_n311), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT18), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT17), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n313), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n315), .A2(new_n321), .A3(new_n326), .A4(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(G1698), .B1(new_n282), .B2(new_n283), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G222), .ZN(new_n332));
  INV_X1    g0132(.A(G77), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n282), .A2(new_n283), .ZN(new_n334));
  INV_X1    g0134(.A(G223), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(G1698), .ZN(new_n336));
  OAI221_X1 g0136(.A(new_n332), .B1(new_n333), .B2(new_n334), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n266), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n253), .B1(new_n273), .B2(G226), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G200), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n338), .A2(G190), .A3(new_n339), .ZN(new_n342));
  INV_X1    g0142(.A(new_n294), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n224), .A2(G33), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n300), .A2(new_n345), .B1(G150), .B2(new_n287), .ZN(new_n346));
  OAI21_X1  g0146(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n343), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n304), .A2(G50), .ZN(new_n349));
  OAI22_X1  g0149(.A1(new_n349), .A2(new_n307), .B1(G50), .B2(new_n306), .ZN(new_n350));
  OR2_X1    g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT9), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n348), .A2(new_n350), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT9), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n341), .A2(new_n342), .A3(new_n353), .A4(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT10), .ZN(new_n357));
  XNOR2_X1  g0157(.A(new_n354), .B(new_n352), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT10), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n358), .A2(new_n359), .A3(new_n342), .A4(new_n341), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n354), .B1(new_n340), .B2(new_n317), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(G179), .B2(new_n340), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n308), .A2(G77), .A3(new_n304), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(G77), .B2(new_n306), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n300), .A2(new_n287), .B1(G20), .B2(G77), .ZN(new_n366));
  XNOR2_X1  g0166(.A(KEYINPUT15), .B(G87), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n345), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n343), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n365), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n331), .A2(G232), .ZN(new_n372));
  INV_X1    g0172(.A(G107), .ZN(new_n373));
  OAI221_X1 g0173(.A(new_n372), .B1(new_n373), .B2(new_n334), .C1(new_n208), .C2(new_n336), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n266), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n253), .B1(new_n273), .B2(G244), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n371), .B1(new_n377), .B2(new_n317), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(G179), .B2(new_n377), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(G200), .ZN(new_n380));
  INV_X1    g0180(.A(G190), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n380), .B(new_n371), .C1(new_n381), .C2(new_n377), .ZN(new_n382));
  AND2_X1   g0182(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n330), .A2(new_n361), .A3(new_n363), .A4(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n271), .A2(G238), .A3(new_n272), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n251), .A2(new_n252), .ZN(new_n386));
  INV_X1    g0186(.A(new_n250), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(G226), .A2(G1698), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n389), .B1(new_n214), .B2(G1698), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n390), .A2(new_n334), .B1(G33), .B2(G97), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n385), .B(new_n388), .C1(new_n391), .C2(new_n265), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n392), .A2(KEYINPUT13), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT13), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n214), .A2(G1698), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(G226), .B2(G1698), .ZN(new_n396));
  OAI22_X1  g0196(.A1(new_n396), .A2(new_n277), .B1(new_n281), .B2(new_n215), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n253), .B1(new_n397), .B2(new_n266), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n394), .B1(new_n398), .B2(new_n385), .ZN(new_n399));
  OAI21_X1  g0199(.A(G169), .B1(new_n393), .B2(new_n399), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n393), .A2(new_n399), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n400), .A2(KEYINPUT14), .B1(new_n401), .B2(G179), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n392), .A2(KEYINPUT13), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n398), .A2(new_n394), .A3(new_n385), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n317), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT71), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT14), .ZN(new_n407));
  AND3_X1   g0207(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n406), .B1(new_n405), .B2(new_n407), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n402), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n345), .A2(G77), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n287), .A2(G50), .B1(G20), .B2(new_n207), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n343), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  XNOR2_X1  g0213(.A(new_n413), .B(KEYINPUT11), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n308), .A2(G68), .A3(new_n304), .ZN(new_n415));
  INV_X1    g0215(.A(G13), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n416), .A2(G1), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n417), .A2(G20), .A3(new_n207), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT12), .ZN(new_n419));
  OR2_X1    g0219(.A1(new_n419), .A2(KEYINPUT70), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(KEYINPUT70), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n418), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n415), .B(new_n422), .C1(new_n420), .C2(new_n418), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n414), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n410), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(G200), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n401), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n403), .A2(new_n404), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n424), .B1(new_n429), .B2(new_n381), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n426), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n384), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(G45), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n436), .A2(G1), .ZN(new_n437));
  AND2_X1   g0237(.A1(KEYINPUT5), .A2(G41), .ZN(new_n438));
  NOR2_X1   g0238(.A1(KEYINPUT5), .A2(G41), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n271), .A2(new_n440), .A3(G270), .ZN(new_n441));
  XNOR2_X1  g0241(.A(KEYINPUT5), .B(G41), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n249), .A2(G45), .A3(G274), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n271), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  OAI211_X1 g0246(.A(G264), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n447));
  INV_X1    g0247(.A(G1698), .ZN(new_n448));
  OAI211_X1 g0248(.A(G257), .B(new_n448), .C1(new_n256), .C2(new_n257), .ZN(new_n449));
  INV_X1    g0249(.A(G303), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n447), .B(new_n449), .C1(new_n450), .C2(new_n334), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n266), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n446), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT80), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G283), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n455), .B(new_n224), .C1(G33), .C2(new_n215), .ZN(new_n456));
  INV_X1    g0256(.A(G116), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G20), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n456), .A2(new_n294), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT20), .ZN(new_n460));
  XNOR2_X1  g0260(.A(new_n459), .B(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n306), .A2(G116), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT74), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n463), .B1(new_n281), .B2(G1), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n249), .A2(KEYINPUT74), .A3(G33), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n307), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n462), .B1(new_n467), .B2(G116), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n317), .B1(new_n461), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT80), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n446), .A2(new_n452), .A3(new_n470), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n454), .A2(new_n469), .A3(KEYINPUT21), .A4(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(G179), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n453), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n461), .A2(new_n468), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AND2_X1   g0276(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n471), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n470), .B1(new_n446), .B2(new_n452), .ZN(new_n479));
  OAI21_X1  g0279(.A(G190), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n454), .A2(G200), .A3(new_n471), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n480), .A2(new_n481), .A3(new_n461), .A4(new_n468), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n454), .A2(new_n469), .A3(new_n471), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT21), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n477), .A2(new_n482), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT82), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n271), .A2(new_n440), .A3(G264), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n210), .A2(new_n448), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n216), .A2(G1698), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n489), .B(new_n490), .C1(new_n256), .C2(new_n257), .ZN(new_n491));
  AND2_X1   g0291(.A1(KEYINPUT81), .A2(G294), .ZN(new_n492));
  NOR2_X1   g0292(.A1(KEYINPUT81), .A2(G294), .ZN(new_n493));
  OAI21_X1  g0293(.A(G33), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n265), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n487), .B1(new_n488), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n271), .A2(new_n440), .A3(G264), .ZN(new_n497));
  NOR2_X1   g0297(.A1(G250), .A2(G1698), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n498), .B1(new_n216), .B2(G1698), .ZN(new_n499));
  XNOR2_X1  g0299(.A(KEYINPUT81), .B(G294), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n499), .A2(new_n334), .B1(new_n500), .B2(G33), .ZN(new_n501));
  OAI211_X1 g0301(.A(KEYINPUT82), .B(new_n497), .C1(new_n501), .C2(new_n265), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n496), .A2(new_n502), .A3(new_n445), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n427), .ZN(new_n504));
  INV_X1    g0304(.A(new_n445), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n488), .A2(new_n505), .A3(new_n495), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n381), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT25), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n306), .B2(G107), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n309), .A2(KEYINPUT25), .A3(new_n373), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n467), .A2(G107), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n224), .B(G87), .C1(new_n256), .C2(new_n257), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT22), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT22), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n334), .A2(new_n516), .A3(new_n224), .A4(G87), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G116), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(G20), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT23), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(new_n224), .B2(G107), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n373), .A2(KEYINPUT23), .A3(G20), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT24), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT24), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n518), .A2(new_n527), .A3(new_n524), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n513), .B1(new_n529), .B2(new_n294), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n508), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(G244), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n532));
  OAI211_X1 g0332(.A(G238), .B(new_n448), .C1(new_n256), .C2(new_n257), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n532), .A2(new_n533), .A3(new_n519), .ZN(new_n534));
  OAI21_X1  g0334(.A(G250), .B1(new_n436), .B2(G1), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n443), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n534), .A2(new_n266), .B1(new_n271), .B2(new_n536), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n537), .A2(new_n473), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n537), .A2(G169), .ZN(new_n539));
  OAI21_X1  g0339(.A(KEYINPUT78), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n537), .A2(new_n473), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT78), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n541), .B(new_n542), .C1(G169), .C2(new_n537), .ZN(new_n543));
  NAND3_X1  g0343(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT79), .ZN(new_n545));
  AND3_X1   g0345(.A1(new_n544), .A2(new_n545), .A3(new_n224), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n545), .B1(new_n544), .B2(new_n224), .ZN(new_n547));
  NOR3_X1   g0347(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n548));
  NOR3_X1   g0348(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n224), .B(G68), .C1(new_n256), .C2(new_n257), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n344), .A2(new_n215), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n550), .B1(KEYINPUT19), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n294), .B1(new_n549), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n367), .A2(new_n309), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n467), .A2(new_n368), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n540), .A2(new_n543), .A3(new_n556), .ZN(new_n557));
  AND3_X1   g0357(.A1(new_n518), .A2(new_n527), .A3(new_n524), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n527), .B1(new_n518), .B2(new_n524), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n294), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n512), .ZN(new_n561));
  OAI22_X1  g0361(.A1(new_n503), .A2(new_n473), .B1(new_n506), .B2(new_n317), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n467), .A2(G87), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n553), .A2(new_n554), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n534), .A2(new_n266), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n271), .A2(new_n536), .ZN(new_n567));
  AND3_X1   g0367(.A1(new_n566), .A2(G190), .A3(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(new_n427), .B2(new_n537), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n531), .A2(new_n557), .A3(new_n563), .A4(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n486), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n297), .A2(G107), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT6), .ZN(new_n574));
  AND2_X1   g0374(.A1(G97), .A2(G107), .ZN(new_n575));
  NOR2_X1   g0375(.A1(G97), .A2(G107), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n373), .A2(KEYINPUT6), .A3(G97), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n579), .A2(G20), .B1(G77), .B2(new_n287), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n343), .B1(new_n573), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n306), .A2(G97), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n582), .B1(new_n467), .B2(G97), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(KEYINPUT77), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n579), .A2(G20), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n287), .A2(G77), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n373), .B1(new_n295), .B2(new_n296), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n294), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT77), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n590), .A2(new_n591), .A3(new_n583), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n585), .A2(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(G250), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n594));
  OAI211_X1 g0394(.A(G244), .B(new_n448), .C1(new_n256), .C2(new_n257), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT4), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n455), .B(new_n594), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(KEYINPUT4), .B1(new_n331), .B2(G244), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n266), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n271), .A2(new_n440), .A3(G257), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n600), .A2(new_n445), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n599), .A2(KEYINPUT76), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(KEYINPUT76), .B1(new_n599), .B2(new_n601), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n317), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n600), .A2(new_n445), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n595), .A2(new_n596), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n334), .A2(KEYINPUT4), .A3(G244), .A4(new_n448), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n606), .A2(new_n607), .A3(new_n455), .A4(new_n594), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n605), .B1(new_n608), .B2(new_n266), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n473), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n593), .A2(new_n604), .A3(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(KEYINPUT75), .B1(new_n609), .B2(new_n427), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n599), .A2(new_n601), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT75), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(new_n614), .A3(G200), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT76), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n599), .A2(KEYINPUT76), .A3(new_n601), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n618), .A2(G190), .A3(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n581), .A2(new_n584), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n616), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n611), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n572), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n435), .A2(new_n625), .ZN(G372));
  NAND2_X1  g0426(.A1(new_n426), .A2(new_n379), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n315), .A2(new_n328), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n627), .A2(new_n432), .A3(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n321), .A2(new_n326), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n361), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n363), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n557), .A2(new_n570), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT85), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT26), .ZN(new_n637));
  NOR4_X1   g0437(.A1(new_n635), .A2(new_n611), .A3(new_n636), .A4(new_n637), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n635), .A2(new_n611), .A3(new_n637), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n621), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n604), .A2(new_n610), .A3(new_n641), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n532), .A2(new_n533), .A3(new_n519), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT83), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n271), .A2(new_n644), .A3(new_n536), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n644), .B1(new_n271), .B2(new_n536), .ZN(new_n646));
  OAI22_X1  g0446(.A1(new_n643), .A2(new_n265), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(G200), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n569), .A2(new_n648), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n647), .A2(new_n317), .B1(new_n473), .B2(new_n537), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n556), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n637), .B1(new_n642), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(KEYINPUT85), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n638), .B1(new_n640), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT84), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n561), .A2(new_n562), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n656), .B1(new_n561), .B2(new_n562), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n485), .B(new_n477), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n569), .A2(new_n648), .B1(new_n650), .B2(new_n556), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n611), .A2(new_n622), .A3(new_n531), .A4(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n651), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n434), .B1(new_n655), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n634), .A2(new_n664), .ZN(G369));
  NAND2_X1  g0465(.A1(new_n477), .A2(new_n485), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n417), .A2(new_n224), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(G213), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(G343), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n475), .A2(new_n673), .ZN(new_n674));
  MUX2_X1   g0474(.A(new_n486), .B(new_n667), .S(new_n674), .Z(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT86), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(G330), .ZN(new_n677));
  INV_X1    g0477(.A(new_n673), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n531), .B(new_n563), .C1(new_n530), .C2(new_n678), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n679), .B(KEYINPUT87), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n563), .A2(new_n678), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n667), .A2(new_n673), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  OR3_X1    g0485(.A1(new_n657), .A2(new_n658), .A3(new_n673), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n683), .A2(new_n687), .ZN(G399));
  INV_X1    g0488(.A(new_n227), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(G41), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n548), .A2(new_n457), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n690), .A2(new_n691), .A3(new_n249), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n692), .B1(new_n222), .B2(new_n690), .ZN(new_n693));
  XOR2_X1   g0493(.A(new_n693), .B(KEYINPUT28), .Z(new_n694));
  INV_X1    g0494(.A(G330), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n486), .A2(new_n571), .A3(new_n623), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n503), .A2(new_n473), .A3(new_n613), .A4(new_n647), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n454), .A2(new_n471), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n618), .A2(KEYINPUT30), .A3(new_n619), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n496), .A2(new_n502), .A3(new_n537), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT88), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n496), .A2(new_n502), .A3(new_n537), .A4(KEYINPUT88), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n704), .A2(new_n474), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n699), .B1(new_n701), .B2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT30), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n704), .A2(new_n474), .A3(new_n705), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n618), .A2(new_n619), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n678), .B1(new_n707), .B2(new_n711), .ZN(new_n712));
  AOI22_X1  g0512(.A1(new_n696), .A2(new_n678), .B1(KEYINPUT31), .B2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n710), .ZN(new_n714));
  AOI21_X1  g0514(.A(KEYINPUT30), .B1(new_n706), .B2(new_n714), .ZN(new_n715));
  OAI22_X1  g0515(.A1(new_n709), .A2(new_n700), .B1(new_n698), .B2(new_n697), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n673), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT31), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n695), .B1(new_n713), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n678), .B1(new_n655), .B2(new_n663), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT29), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n557), .A2(new_n570), .ZN(new_n724));
  INV_X1    g0524(.A(new_n611), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n724), .A2(new_n725), .A3(new_n637), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n661), .A2(new_n604), .A3(new_n610), .A4(new_n641), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(KEYINPUT26), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n726), .A2(new_n728), .A3(new_n651), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n662), .B1(new_n667), .B2(new_n563), .ZN(new_n730));
  OAI211_X1 g0530(.A(KEYINPUT29), .B(new_n678), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n720), .B1(new_n723), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n732), .B(KEYINPUT89), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n694), .B1(new_n734), .B2(G1), .ZN(G364));
  NOR2_X1   g0535(.A1(new_n416), .A2(G20), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n249), .B1(new_n736), .B2(G45), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n690), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n689), .A2(new_n277), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G355), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n741), .B1(G116), .B2(new_n227), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n244), .A2(new_n436), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n689), .A2(new_n334), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n745), .B1(new_n222), .B2(new_n251), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n742), .B1(new_n743), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n263), .B1(new_n224), .B2(G169), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n748), .A2(KEYINPUT90), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(KEYINPUT90), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G13), .A2(G33), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(G20), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n739), .B1(new_n747), .B2(new_n756), .ZN(new_n757));
  XOR2_X1   g0557(.A(new_n757), .B(KEYINPUT91), .Z(new_n758));
  INV_X1    g0558(.A(new_n751), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n381), .A2(G200), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(new_n473), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G20), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n215), .ZN(new_n764));
  NAND2_X1  g0564(.A1(G20), .A2(G179), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT92), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n427), .A2(G190), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n764), .B1(new_n769), .B2(G68), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT94), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n224), .A2(G179), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G190), .A2(G200), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G159), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g0576(.A(KEYINPUT93), .B(KEYINPUT32), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n381), .A2(new_n427), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(new_n772), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n277), .B1(new_n781), .B2(G87), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n767), .A2(new_n772), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n778), .B(new_n782), .C1(new_n373), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n766), .A2(new_n773), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n766), .A2(new_n760), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n786), .A2(G77), .B1(new_n788), .B2(G58), .ZN(new_n789));
  INV_X1    g0589(.A(G50), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n766), .A2(new_n779), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n771), .A2(new_n784), .A3(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n794), .A2(KEYINPUT95), .ZN(new_n795));
  INV_X1    g0595(.A(new_n500), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n277), .B1(new_n780), .B2(new_n450), .C1(new_n763), .C2(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(G311), .B2(new_n786), .ZN(new_n798));
  XNOR2_X1  g0598(.A(KEYINPUT33), .B(G317), .ZN(new_n799));
  INV_X1    g0599(.A(new_n791), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n769), .A2(new_n799), .B1(new_n800), .B2(G326), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n788), .A2(G322), .ZN(new_n802));
  INV_X1    g0602(.A(new_n783), .ZN(new_n803));
  INV_X1    g0603(.A(new_n774), .ZN(new_n804));
  AOI22_X1  g0604(.A1(G283), .A2(new_n803), .B1(new_n804), .B2(G329), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT96), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n798), .A2(new_n801), .A3(new_n802), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n794), .A2(KEYINPUT95), .ZN(new_n808));
  AND3_X1   g0608(.A1(new_n795), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n754), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n758), .B1(new_n759), .B2(new_n809), .C1(new_n676), .C2(new_n810), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n811), .A2(KEYINPUT97), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n811), .A2(KEYINPUT97), .ZN(new_n813));
  OR2_X1    g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n739), .B1(new_n676), .B2(G330), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(G330), .B2(new_n676), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n814), .A2(KEYINPUT98), .A3(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(KEYINPUT98), .B1(new_n814), .B2(new_n816), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(G396));
  OAI21_X1  g0621(.A(new_n382), .B1(new_n371), .B2(new_n678), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n379), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n379), .A2(new_n673), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n721), .A2(new_n825), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n823), .A2(new_n824), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n678), .B(new_n827), .C1(new_n655), .C2(new_n663), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n720), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n829), .A2(new_n739), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n826), .A2(new_n720), .A3(new_n828), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n739), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n751), .A2(new_n752), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n833), .B1(new_n834), .B2(new_n333), .ZN(new_n835));
  XNOR2_X1  g0635(.A(KEYINPUT99), .B(G283), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  AOI22_X1  g0637(.A1(G116), .A2(new_n786), .B1(new_n769), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(G294), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n838), .B1(new_n839), .B2(new_n787), .C1(new_n450), .C2(new_n791), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n277), .B1(new_n780), .B2(new_n373), .ZN(new_n841));
  INV_X1    g0641(.A(G311), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n783), .A2(new_n209), .B1(new_n774), .B2(new_n842), .ZN(new_n843));
  NOR4_X1   g0643(.A1(new_n840), .A2(new_n764), .A3(new_n841), .A4(new_n843), .ZN(new_n844));
  AOI22_X1  g0644(.A1(G137), .A2(new_n800), .B1(new_n788), .B2(G143), .ZN(new_n845));
  INV_X1    g0645(.A(G150), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n845), .B1(new_n846), .B2(new_n768), .C1(new_n775), .C2(new_n785), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT34), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n334), .B1(new_n780), .B2(new_n790), .ZN(new_n849));
  INV_X1    g0649(.A(G132), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n783), .A2(new_n207), .B1(new_n774), .B2(new_n850), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n849), .B(new_n851), .C1(G58), .C2(new_n762), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n844), .B1(new_n848), .B2(new_n852), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n835), .B1(new_n853), .B2(new_n759), .C1(new_n827), .C2(new_n753), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n832), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(G384));
  OR2_X1    g0656(.A1(new_n579), .A2(KEYINPUT35), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n579), .A2(KEYINPUT35), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n857), .A2(G116), .A3(new_n225), .A4(new_n858), .ZN(new_n859));
  XOR2_X1   g0659(.A(new_n859), .B(KEYINPUT36), .Z(new_n860));
  OAI211_X1 g0660(.A(new_n222), .B(G77), .C1(new_n213), .C2(new_n207), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n790), .A2(G68), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n249), .B(G13), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT39), .ZN(new_n865));
  INV_X1    g0665(.A(new_n671), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n316), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT37), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n320), .A2(new_n867), .A3(new_n868), .A4(new_n313), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n319), .A2(new_n318), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT16), .B1(new_n286), .B2(new_n292), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT100), .B1(new_n872), .B2(new_n343), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT100), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n207), .B1(new_n284), .B2(KEYINPUT7), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n291), .B1(new_n875), .B2(new_n279), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n874), .B(new_n294), .C1(new_n876), .C2(KEYINPUT16), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n873), .A2(new_n293), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n871), .B1(new_n878), .B2(new_n311), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT101), .B1(new_n879), .B2(new_n314), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT101), .ZN(new_n881));
  INV_X1    g0681(.A(new_n311), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n294), .B1(new_n876), .B2(KEYINPUT16), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n883), .A2(KEYINPUT100), .B1(KEYINPUT16), .B2(new_n876), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n882), .B1(new_n884), .B2(new_n877), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n881), .B(new_n313), .C1(new_n885), .C2(new_n871), .ZN(new_n886));
  OR2_X1    g0686(.A1(new_n885), .A2(new_n671), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n880), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n870), .B1(new_n888), .B2(KEYINPUT37), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT38), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n887), .B1(new_n628), .B2(new_n630), .ZN(new_n891));
  NOR3_X1   g0691(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n314), .A2(new_n324), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n893), .A2(KEYINPUT102), .A3(new_n868), .A4(new_n867), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT102), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n869), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n320), .A2(new_n867), .A3(new_n313), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(KEYINPUT37), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n894), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n329), .A2(new_n316), .A3(new_n866), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT38), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n865), .B1(new_n892), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n426), .A2(new_n673), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n890), .B1(new_n889), .B2(new_n891), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n885), .A2(new_n671), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n329), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n313), .B1(new_n885), .B2(new_n871), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n905), .B1(new_n907), .B2(KEYINPUT101), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n868), .B1(new_n908), .B2(new_n886), .ZN(new_n909));
  OAI211_X1 g0709(.A(KEYINPUT38), .B(new_n906), .C1(new_n909), .C2(new_n870), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n904), .A2(new_n910), .A3(KEYINPUT39), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n902), .A2(new_n903), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n828), .A2(new_n824), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n904), .A2(new_n910), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n425), .B(new_n673), .C1(new_n410), .C2(new_n431), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n425), .A2(new_n673), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n403), .A2(new_n404), .A3(G179), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n405), .B2(new_n407), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n429), .A2(new_n407), .A3(G169), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(KEYINPUT71), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n432), .B(new_n916), .C1(new_n922), .C2(new_n424), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n915), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n913), .A2(new_n914), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n631), .A2(new_n671), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n912), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT103), .ZN(new_n928));
  NAND4_X1  g0728(.A1(new_n723), .A2(new_n928), .A3(new_n434), .A4(new_n731), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n724), .A2(new_n725), .A3(KEYINPUT85), .A4(KEYINPUT26), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n636), .B1(new_n727), .B2(new_n637), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n930), .B1(new_n931), .B2(new_n639), .ZN(new_n932));
  INV_X1    g0732(.A(new_n651), .ZN(new_n933));
  AND4_X1   g0733(.A1(new_n611), .A2(new_n622), .A3(new_n531), .A4(new_n661), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n933), .B1(new_n934), .B2(new_n659), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n673), .B1(new_n932), .B2(new_n935), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n434), .B(new_n731), .C1(new_n936), .C2(KEYINPUT29), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(KEYINPUT103), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n633), .B1(new_n929), .B2(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n927), .B(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n924), .A2(new_n827), .ZN(new_n941));
  OAI21_X1  g0741(.A(KEYINPUT104), .B1(new_n712), .B2(KEYINPUT31), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT104), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n717), .A2(new_n943), .A3(new_n718), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n941), .B1(new_n945), .B2(new_n713), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n914), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT40), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n901), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n910), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n951), .A2(new_n946), .A3(KEYINPUT40), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  AND3_X1   g0753(.A1(new_n717), .A2(new_n943), .A3(new_n718), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n943), .B1(new_n717), .B2(new_n718), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n712), .A2(KEYINPUT31), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n625), .B2(new_n673), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n434), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n953), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n953), .A2(new_n959), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n960), .A2(G330), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n940), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n249), .B2(new_n736), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n940), .A2(new_n962), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n864), .B1(new_n964), .B2(new_n965), .ZN(G367));
  OAI221_X1 g0766(.A(new_n755), .B1(new_n227), .B2(new_n367), .C1(new_n236), .C2(new_n745), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n739), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n786), .A2(G50), .B1(new_n800), .B2(G143), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n969), .B1(new_n846), .B2(new_n787), .C1(new_n775), .C2(new_n768), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n763), .A2(new_n207), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n334), .B1(new_n780), .B2(new_n213), .ZN(new_n972));
  XNOR2_X1  g0772(.A(KEYINPUT107), .B(G137), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n783), .A2(new_n333), .B1(new_n774), .B2(new_n973), .ZN(new_n974));
  NOR4_X1   g0774(.A1(new_n970), .A2(new_n971), .A3(new_n972), .A4(new_n974), .ZN(new_n975));
  AOI22_X1  g0775(.A1(G303), .A2(new_n788), .B1(new_n800), .B2(G311), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n785), .B2(new_n836), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n781), .A2(KEYINPUT46), .A3(G116), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT46), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n780), .B2(new_n457), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n978), .B(new_n980), .C1(new_n373), .C2(new_n763), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n768), .A2(new_n796), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n803), .A2(G97), .ZN(new_n983));
  INV_X1    g0783(.A(G317), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n983), .B(new_n277), .C1(new_n984), .C2(new_n774), .ZN(new_n985));
  NOR4_X1   g0785(.A1(new_n977), .A2(new_n981), .A3(new_n982), .A4(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n975), .A2(new_n986), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n987), .A2(KEYINPUT47), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n759), .B1(new_n987), .B2(KEYINPUT47), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n968), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n565), .A2(new_n673), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT105), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n933), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n652), .B2(new_n992), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n990), .B1(new_n994), .B2(new_n810), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n682), .B1(new_n667), .B2(new_n673), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n685), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n677), .B(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n733), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n641), .A2(new_n673), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n623), .A2(new_n1000), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n604), .A2(new_n610), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1002), .A2(new_n1000), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n687), .A2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT45), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n683), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n687), .A2(new_n1004), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT44), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1006), .A2(new_n1007), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n683), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n999), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n734), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n690), .B(new_n1016), .Z(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n738), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n685), .A2(new_n1004), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n611), .B1(new_n1004), .B2(new_n563), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1020), .A2(KEYINPUT42), .B1(new_n678), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(KEYINPUT42), .B2(new_n1020), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n994), .A2(KEYINPUT43), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n994), .A2(KEYINPUT43), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NOR3_X1   g0827(.A1(new_n1023), .A2(KEYINPUT43), .A3(new_n994), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1007), .A2(new_n1004), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1029), .B(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n995), .B1(new_n1019), .B2(new_n1031), .ZN(G387));
  INV_X1    g0832(.A(new_n690), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n999), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n998), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1034), .B1(new_n734), .B2(new_n1035), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n240), .A2(new_n251), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n1037), .A2(new_n744), .B1(new_n691), .B2(new_n740), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n436), .B1(new_n207), .B2(new_n333), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT50), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n310), .B2(G50), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n300), .A2(KEYINPUT50), .A3(new_n790), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n691), .B(new_n1039), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n1038), .A2(new_n1043), .B1(G107), .B2(new_n227), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n833), .B1(new_n1044), .B2(new_n755), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n780), .A2(new_n333), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(G150), .B2(new_n804), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1047), .A2(new_n334), .A3(new_n983), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n790), .A2(new_n787), .B1(new_n768), .B2(new_n310), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n207), .A2(new_n785), .B1(new_n791), .B2(new_n775), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n763), .A2(new_n367), .ZN(new_n1051));
  NOR4_X1   g0851(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(G326), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n277), .B1(new_n774), .B2(new_n1053), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n450), .A2(new_n785), .B1(new_n787), .B2(new_n984), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT108), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n769), .A2(G311), .B1(new_n800), .B2(G322), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT48), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n762), .A2(new_n837), .B1(new_n781), .B2(new_n500), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT49), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n1054), .B(new_n1067), .C1(G116), .C2(new_n803), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1052), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1045), .B1(new_n1070), .B2(new_n759), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n682), .B2(new_n754), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n1035), .B2(new_n738), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1036), .A2(new_n1073), .ZN(G393));
  NAND3_X1  g0874(.A1(new_n1013), .A2(KEYINPUT109), .A3(new_n1011), .ZN(new_n1075));
  OR3_X1    g0875(.A1(new_n1012), .A2(KEYINPUT109), .A3(new_n683), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n690), .B(new_n1014), .C1(new_n1077), .C2(new_n999), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n247), .A2(new_n744), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n755), .B1(new_n215), .B2(new_n227), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n457), .A2(new_n763), .B1(new_n768), .B2(new_n450), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n781), .A2(new_n837), .B1(new_n804), .B2(G322), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1082), .B(new_n277), .C1(new_n373), .C2(new_n783), .ZN(new_n1083));
  XOR2_X1   g0883(.A(new_n1083), .B(KEYINPUT112), .Z(new_n1084));
  AOI211_X1 g0884(.A(new_n1081), .B(new_n1084), .C1(G294), .C2(new_n786), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n842), .A2(new_n787), .B1(new_n791), .B2(new_n984), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT52), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n846), .A2(new_n791), .B1(new_n787), .B2(new_n775), .ZN(new_n1088));
  XOR2_X1   g0888(.A(new_n1088), .B(KEYINPUT110), .Z(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(KEYINPUT51), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1089), .A2(KEYINPUT51), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(G68), .A2(new_n781), .B1(new_n804), .B2(G143), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1092), .B(new_n334), .C1(new_n209), .C2(new_n783), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n1093), .B(KEYINPUT111), .Z(new_n1094));
  NOR2_X1   g0894(.A1(new_n763), .A2(new_n333), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n769), .B2(G50), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n310), .B2(new_n785), .ZN(new_n1097));
  NOR3_X1   g0897(.A1(new_n1091), .A2(new_n1094), .A3(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n1085), .A2(new_n1087), .B1(new_n1090), .B2(new_n1098), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n739), .B1(new_n1079), .B2(new_n1080), .C1(new_n1099), .C2(new_n759), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(new_n754), .B2(new_n1004), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n1077), .B2(new_n738), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1078), .A2(new_n1102), .ZN(G390));
  AOI21_X1  g0903(.A(new_n695), .B1(new_n945), .B2(new_n713), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n825), .B1(new_n923), .B2(new_n915), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n673), .B(new_n825), .C1(new_n932), .C2(new_n935), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n824), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n924), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n903), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1109), .A2(new_n1110), .B1(new_n902), .B2(new_n911), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n924), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n678), .B(new_n823), .C1(new_n729), .C2(new_n730), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1112), .B1(new_n1113), .B2(new_n824), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n889), .A2(new_n891), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n901), .B1(new_n1115), .B2(KEYINPUT38), .ZN(new_n1116));
  NOR3_X1   g0916(.A1(new_n1114), .A2(new_n1116), .A3(new_n903), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1106), .B1(new_n1111), .B2(new_n1117), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n957), .B(new_n719), .C1(new_n625), .C2(new_n673), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1119), .A2(G330), .A3(new_n827), .A4(new_n924), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n1113), .A2(new_n824), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1110), .B(new_n951), .C1(new_n1121), .C2(new_n1112), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n902), .A2(new_n911), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n903), .B1(new_n913), .B2(new_n924), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1120), .B(new_n1122), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1118), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1119), .A2(G330), .A3(new_n827), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1112), .A2(new_n1127), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n913), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n924), .B1(new_n1104), .B2(new_n827), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1121), .A2(new_n1120), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n1128), .A2(new_n1129), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1104), .A2(new_n434), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1132), .A2(new_n939), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1033), .B1(new_n1126), .B2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n1135), .B2(new_n1126), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1118), .A2(new_n1125), .A3(new_n738), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n833), .B1(new_n834), .B2(new_n310), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(G97), .A2(new_n786), .B1(new_n769), .B2(G107), .ZN(new_n1140));
  INV_X1    g0940(.A(G283), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n1140), .B1(new_n457), .B2(new_n787), .C1(new_n1141), .C2(new_n791), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n277), .B1(new_n780), .B2(new_n209), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n783), .A2(new_n207), .B1(new_n774), .B2(new_n839), .ZN(new_n1144));
  NOR4_X1   g0944(.A1(new_n1142), .A2(new_n1095), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1145));
  OR2_X1    g0945(.A1(new_n1145), .A2(KEYINPUT114), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n334), .B1(new_n783), .B2(new_n790), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(G125), .B2(new_n804), .ZN(new_n1148));
  XOR2_X1   g0948(.A(new_n1148), .B(KEYINPUT113), .Z(new_n1149));
  NAND2_X1  g0949(.A1(new_n781), .A2(G150), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1150), .B(KEYINPUT53), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G159), .B2(new_n762), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n973), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n769), .A2(new_n1153), .B1(new_n800), .B2(G128), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(KEYINPUT54), .B(G143), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n786), .A2(new_n1156), .B1(new_n788), .B2(G132), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1149), .A2(new_n1152), .A3(new_n1154), .A4(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1146), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(KEYINPUT114), .B2(new_n1145), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n1139), .B1(new_n759), .B2(new_n1160), .C1(new_n1123), .C2(new_n753), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n1138), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT115), .ZN(new_n1163));
  AND2_X1   g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1137), .B1(new_n1164), .B2(new_n1165), .ZN(G378));
  INV_X1    g0966(.A(KEYINPUT117), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n361), .A2(new_n363), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n354), .A2(new_n671), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1168), .B(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1171));
  XOR2_X1   g0971(.A(new_n1170), .B(new_n1171), .Z(new_n1172));
  NAND4_X1  g0972(.A1(new_n949), .A2(G330), .A3(new_n952), .A4(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1170), .B(new_n1171), .ZN(new_n1174));
  OAI211_X1 g0974(.A(KEYINPUT40), .B(new_n1105), .C1(new_n956), .C2(new_n958), .ZN(new_n1175));
  OAI21_X1  g0975(.A(G330), .B1(new_n1175), .B2(new_n1116), .ZN(new_n1176));
  AOI21_X1  g0976(.A(KEYINPUT40), .B1(new_n914), .B2(new_n946), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1174), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  AND3_X1   g0978(.A1(new_n927), .A2(new_n1173), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1112), .B1(new_n828), .B2(new_n824), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n1180), .A2(new_n914), .B1(new_n631), .B2(new_n671), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n1173), .A2(new_n1178), .B1(new_n912), .B2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1167), .B1(new_n1179), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n939), .A2(new_n1134), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(KEYINPUT119), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT119), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n939), .A2(new_n1186), .A3(new_n1134), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1185), .B(new_n1187), .C1(new_n1126), .C2(new_n1135), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1181), .A2(new_n912), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n948), .B(new_n941), .C1(new_n713), .C2(new_n945), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n695), .B1(new_n1190), .B2(new_n951), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1172), .B1(new_n1191), .B2(new_n949), .ZN(new_n1192));
  NOR3_X1   g0992(.A1(new_n1176), .A2(new_n1177), .A3(new_n1174), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1189), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n927), .A2(new_n1173), .A3(new_n1178), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1194), .A2(KEYINPUT117), .A3(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1183), .A2(new_n1188), .A3(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT57), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1198), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1033), .B1(new_n1200), .B2(new_n1188), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1183), .A2(new_n1196), .A3(new_n738), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n834), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n739), .B1(new_n1204), .B2(G50), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n769), .A2(G97), .B1(new_n788), .B2(G107), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n457), .B2(new_n791), .C1(new_n367), .C2(new_n785), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n277), .A2(new_n252), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n1046), .A2(new_n1208), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n783), .A2(new_n213), .B1(new_n774), .B2(new_n1141), .ZN(new_n1210));
  NOR4_X1   g1010(.A1(new_n1207), .A2(new_n971), .A3(new_n1209), .A4(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(G50), .B1(new_n281), .B2(new_n252), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1211), .A2(KEYINPUT58), .B1(new_n1208), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n769), .A2(G132), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n786), .A2(G137), .B1(new_n788), .B2(G128), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n762), .A2(G150), .B1(new_n781), .B2(new_n1156), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n800), .A2(G125), .ZN(new_n1217));
  AND4_X1   g1017(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .A4(new_n1217), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT116), .Z(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1220), .A2(KEYINPUT59), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n281), .B(new_n252), .C1(new_n783), .C2(new_n775), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(G124), .B2(new_n804), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT59), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1223), .B1(new_n1219), .B2(new_n1224), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1213), .B1(KEYINPUT58), .B2(new_n1211), .C1(new_n1221), .C2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1205), .B1(new_n1226), .B2(new_n751), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n1172), .B2(new_n753), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1203), .A2(KEYINPUT118), .A3(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(KEYINPUT118), .B1(new_n1203), .B2(new_n1228), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1202), .B1(new_n1229), .B2(new_n1230), .ZN(G375));
  AOI211_X1 g1031(.A(new_n633), .B(new_n1133), .C1(new_n938), .C2(new_n929), .ZN(new_n1232));
  OAI21_X1  g1032(.A(KEYINPUT121), .B1(new_n1232), .B2(new_n1132), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1132), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT121), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1234), .A2(new_n1184), .A3(new_n1235), .ZN(new_n1236));
  XOR2_X1   g1036(.A(new_n1017), .B(KEYINPUT120), .Z(new_n1237));
  NAND4_X1  g1037(.A1(new_n1233), .A2(new_n1236), .A3(new_n1135), .A4(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1112), .A2(new_n752), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n850), .A2(new_n791), .B1(new_n768), .B2(new_n1155), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(G159), .A2(new_n781), .B1(new_n804), .B2(G128), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1241), .B(new_n334), .C1(new_n213), .C2(new_n783), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n1240), .B(new_n1242), .C1(new_n788), .C2(new_n1153), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n790), .A2(new_n763), .B1(new_n785), .B2(new_n846), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n1244), .B(KEYINPUT122), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n277), .B1(new_n783), .B2(new_n333), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n780), .A2(new_n215), .B1(new_n774), .B2(new_n450), .ZN(new_n1247));
  NOR3_X1   g1047(.A1(new_n1051), .A2(new_n1246), .A3(new_n1247), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n457), .A2(new_n768), .B1(new_n791), .B2(new_n839), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n373), .A2(new_n785), .B1(new_n787), .B2(new_n1141), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n1243), .A2(new_n1245), .B1(new_n1248), .B2(new_n1251), .ZN(new_n1252));
  OAI221_X1 g1052(.A(new_n739), .B1(G68), .B2(new_n1204), .C1(new_n1252), .C2(new_n759), .ZN(new_n1253));
  XOR2_X1   g1053(.A(new_n1253), .B(KEYINPUT123), .Z(new_n1254));
  AOI22_X1  g1054(.A1(new_n1132), .A2(new_n738), .B1(new_n1239), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1238), .A2(new_n1255), .ZN(G381));
  INV_X1    g1056(.A(G390), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(G396), .A2(G393), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1257), .A2(new_n1258), .A3(new_n855), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1137), .A2(new_n1162), .ZN(new_n1260));
  OR2_X1    g1060(.A1(new_n1260), .A2(G381), .ZN(new_n1261));
  OR4_X1    g1061(.A1(G387), .A2(new_n1259), .A3(new_n1261), .A4(G375), .ZN(G407));
  INV_X1    g1062(.A(new_n1260), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n672), .A2(G213), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1263), .A2(new_n1265), .ZN(new_n1266));
  OAI211_X1 g1066(.A(G407), .B(G213), .C1(G375), .C2(new_n1266), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1267), .B(KEYINPUT124), .ZN(G409));
  NAND2_X1  g1068(.A1(new_n1135), .A2(KEYINPUT60), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1233), .A2(new_n1269), .A3(new_n1236), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1232), .A2(new_n1132), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1033), .B1(new_n1271), .B2(KEYINPUT60), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1270), .A2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(G384), .B1(new_n1273), .B2(new_n1255), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1255), .ZN(new_n1275));
  AOI211_X1 g1075(.A(new_n855), .B(new_n1275), .C1(new_n1270), .C2(new_n1272), .ZN(new_n1276));
  INV_X1    g1076(.A(G2897), .ZN(new_n1277));
  OAI22_X1  g1077(.A1(new_n1274), .A2(new_n1276), .B1(new_n1277), .B2(new_n1264), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1273), .A2(new_n1255), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n855), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1273), .A2(G384), .A3(new_n1255), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1264), .A2(new_n1277), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1280), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1278), .A2(new_n1283), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(new_n1284), .B(KEYINPUT125), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1202), .B(G378), .C1(new_n1229), .C2(new_n1230), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n738), .B1(new_n1179), .B2(new_n1182), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1237), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1228), .B(new_n1287), .C1(new_n1197), .C2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1263), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1286), .A2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n1264), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1285), .A2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1265), .B1(new_n1286), .B2(new_n1290), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1274), .A2(new_n1276), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1294), .A2(KEYINPUT63), .A3(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1291), .A2(new_n1264), .A3(new_n1295), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT63), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1257), .A2(G387), .ZN(new_n1300));
  OAI211_X1 g1100(.A(G390), .B(new_n995), .C1(new_n1019), .C2(new_n1031), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(G393), .B(new_n820), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1302), .A2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1300), .A2(new_n1301), .A3(new_n1303), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1307), .A2(KEYINPUT61), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1293), .A2(new_n1296), .A3(new_n1299), .A4(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1306), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1303), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT127), .ZN(new_n1312));
  NOR3_X1   g1112(.A1(new_n1310), .A2(new_n1311), .A3(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(KEYINPUT127), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT61), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1316), .B1(new_n1294), .B2(new_n1284), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT62), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1297), .A2(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1294), .A2(KEYINPUT62), .A3(new_n1295), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1317), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT126), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1315), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1278), .A2(new_n1283), .ZN(new_n1324));
  AOI21_X1  g1124(.A(KEYINPUT61), .B1(new_n1292), .B2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1320), .ZN(new_n1326));
  AOI21_X1  g1126(.A(KEYINPUT62), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1327));
  OAI211_X1 g1127(.A(new_n1322), .B(new_n1325), .C1(new_n1326), .C2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1328), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1309), .B1(new_n1323), .B2(new_n1329), .ZN(G405));
  NAND2_X1  g1130(.A1(G375), .A2(new_n1263), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(new_n1286), .ZN(new_n1332));
  XNOR2_X1  g1132(.A(new_n1332), .B(new_n1295), .ZN(new_n1333));
  XNOR2_X1  g1133(.A(new_n1333), .B(new_n1307), .ZN(G402));
endmodule


