//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 0 1 1 0 1 1 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 1 0 1 0 0 0 0 1 0 1 0 1 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:54 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1278, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  OR3_X1    g0007(.A1(new_n207), .A2(KEYINPUT65), .A3(G13), .ZN(new_n208));
  OAI21_X1  g0008(.A(KEYINPUT65), .B1(new_n207), .B2(G13), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT66), .Z(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  XNOR2_X1  g0013(.A(KEYINPUT67), .B(G244), .ZN(new_n214));
  AND2_X1   g0014(.A1(new_n214), .A2(G77), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G87), .A2(G250), .ZN(new_n219));
  NAND4_X1  g0019(.A1(new_n216), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n207), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(new_n203), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G50), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(new_n221), .A2(KEYINPUT1), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n221), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n213), .A2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT68), .ZN(new_n240));
  XOR2_X1   g0040(.A(G50), .B(G58), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G87), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G97), .B(G107), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  XNOR2_X1  g0046(.A(KEYINPUT3), .B(G33), .ZN(new_n247));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n247), .A2(G222), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(G1698), .ZN(new_n250));
  INV_X1    g0050(.A(G223), .ZN(new_n251));
  OAI221_X1 g0051(.A(new_n249), .B1(new_n202), .B2(new_n247), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  AND2_X1   g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(new_n222), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(KEYINPUT69), .B1(new_n253), .B2(new_n222), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT69), .ZN(new_n258));
  NAND4_X1  g0058(.A1(new_n257), .A2(new_n258), .A3(G1), .A4(G13), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G41), .A2(G45), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(G1), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n260), .A2(G274), .A3(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(KEYINPUT71), .B1(new_n261), .B2(G1), .ZN(new_n264));
  OR3_X1    g0064(.A1(new_n261), .A2(KEYINPUT71), .A3(G1), .ZN(new_n265));
  AND3_X1   g0065(.A1(new_n260), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT70), .B(G226), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n255), .A2(new_n263), .A3(new_n268), .ZN(new_n269));
  OR2_X1    g0069(.A1(new_n269), .A2(G179), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT73), .ZN(new_n271));
  OR2_X1    g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n271), .ZN(new_n273));
  INV_X1    g0073(.A(G1), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G13), .A3(G20), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G50), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n222), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n280), .B1(new_n274), .B2(G20), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n278), .B1(new_n282), .B2(new_n277), .ZN(new_n283));
  INV_X1    g0083(.A(new_n201), .ZN(new_n284));
  OAI21_X1  g0084(.A(G20), .B1(new_n284), .B2(new_n225), .ZN(new_n285));
  INV_X1    g0085(.A(G150), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n223), .A2(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(KEYINPUT72), .A2(G58), .ZN(new_n290));
  XOR2_X1   g0090(.A(new_n290), .B(KEYINPUT8), .Z(new_n291));
  OAI221_X1 g0091(.A(new_n285), .B1(new_n286), .B2(new_n288), .C1(new_n289), .C2(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n283), .B1(new_n292), .B2(new_n280), .ZN(new_n293));
  INV_X1    g0093(.A(G169), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n293), .B1(new_n294), .B2(new_n269), .ZN(new_n295));
  AND3_X1   g0095(.A1(new_n272), .A2(new_n273), .A3(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n247), .A2(G238), .A3(G1698), .ZN(new_n297));
  INV_X1    g0097(.A(G107), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n247), .A2(new_n248), .ZN(new_n299));
  INV_X1    g0099(.A(G232), .ZN(new_n300));
  OAI221_X1 g0100(.A(new_n297), .B1(new_n298), .B2(new_n247), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n254), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n266), .A2(new_n214), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n302), .A2(new_n263), .A3(new_n303), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n304), .A2(G179), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n276), .A2(new_n202), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(new_n282), .B2(new_n202), .ZN(new_n307));
  INV_X1    g0107(.A(new_n280), .ZN(new_n308));
  XOR2_X1   g0108(.A(KEYINPUT8), .B(G58), .Z(new_n309));
  AOI22_X1  g0109(.A1(new_n309), .A2(new_n287), .B1(G20), .B2(G77), .ZN(new_n310));
  XNOR2_X1  g0110(.A(KEYINPUT15), .B(G87), .ZN(new_n311));
  OR2_X1    g0111(.A1(new_n311), .A2(new_n289), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n308), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n307), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n304), .A2(new_n294), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n305), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT74), .B(G200), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n304), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G190), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n320), .B(new_n314), .C1(new_n321), .C2(new_n304), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n317), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n269), .A2(new_n319), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n293), .B1(KEYINPUT75), .B2(KEYINPUT9), .ZN(new_n325));
  AND3_X1   g0125(.A1(new_n325), .A2(KEYINPUT75), .A3(KEYINPUT9), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n325), .B1(KEYINPUT75), .B2(KEYINPUT9), .ZN(new_n327));
  OAI221_X1 g0127(.A(new_n324), .B1(new_n321), .B2(new_n269), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n328), .A2(KEYINPUT10), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(KEYINPUT10), .ZN(new_n330));
  AOI211_X1 g0130(.A(new_n296), .B(new_n323), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT77), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n266), .A2(G238), .ZN(new_n333));
  NAND2_X1  g0133(.A1(G33), .A2(G97), .ZN(new_n334));
  INV_X1    g0134(.A(G226), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n334), .B1(new_n299), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n250), .A2(new_n300), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n254), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n333), .A2(new_n338), .A3(new_n263), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT13), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT13), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n333), .A2(new_n338), .A3(new_n341), .A4(new_n263), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n340), .A2(G190), .A3(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n288), .A2(new_n277), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n289), .A2(new_n202), .B1(new_n223), .B2(G68), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n280), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n346), .A2(KEYINPUT11), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(KEYINPUT11), .ZN(new_n348));
  INV_X1    g0148(.A(G68), .ZN(new_n349));
  OAI22_X1  g0149(.A1(new_n347), .A2(new_n348), .B1(new_n349), .B2(new_n282), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT76), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT12), .ZN(new_n352));
  AOI211_X1 g0152(.A(new_n351), .B(new_n352), .C1(new_n276), .C2(new_n349), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n276), .A2(new_n349), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n354), .A2(KEYINPUT12), .ZN(new_n355));
  AOI21_X1  g0155(.A(KEYINPUT76), .B1(new_n354), .B2(KEYINPUT12), .ZN(new_n356));
  NOR3_X1   g0156(.A1(new_n353), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n350), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n343), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G200), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n360), .B1(new_n340), .B2(new_n342), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n332), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n361), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n363), .A2(KEYINPUT77), .A3(new_n358), .A4(new_n343), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT78), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n362), .A2(new_n364), .A3(KEYINPUT78), .ZN(new_n368));
  INV_X1    g0168(.A(new_n358), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n294), .B1(new_n340), .B2(new_n342), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT14), .ZN(new_n371));
  AND2_X1   g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n340), .A2(G179), .A3(new_n342), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(new_n370), .B2(new_n371), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n369), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n367), .A2(new_n368), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G33), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT3), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT3), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(G33), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(KEYINPUT7), .B1(new_n382), .B2(new_n223), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT7), .ZN(new_n384));
  AOI211_X1 g0184(.A(new_n384), .B(G20), .C1(new_n379), .C2(new_n381), .ZN(new_n385));
  OAI21_X1  g0185(.A(G68), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT16), .ZN(new_n387));
  INV_X1    g0187(.A(G58), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n388), .A2(new_n349), .ZN(new_n389));
  OAI21_X1  g0189(.A(G20), .B1(new_n389), .B2(new_n203), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n287), .A2(G159), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n386), .A2(new_n387), .A3(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n384), .B1(new_n247), .B2(G20), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n380), .A2(G33), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n378), .A2(KEYINPUT3), .ZN(new_n397));
  OAI211_X1 g0197(.A(KEYINPUT7), .B(new_n223), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n349), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(KEYINPUT16), .B1(new_n399), .B2(new_n392), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n393), .A2(KEYINPUT79), .A3(new_n387), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n394), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n386), .A2(KEYINPUT79), .A3(new_n387), .A4(new_n393), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(new_n280), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n291), .A2(new_n275), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(new_n281), .B2(new_n291), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n406), .B(KEYINPUT80), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n260), .A2(G232), .A3(new_n264), .A4(new_n265), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n263), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT81), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n409), .A2(KEYINPUT81), .A3(new_n263), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n247), .A2(G226), .A3(G1698), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n379), .A2(new_n381), .A3(G223), .A4(new_n248), .ZN(new_n415));
  NAND2_X1  g0215(.A1(G33), .A2(G87), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n254), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n412), .A2(new_n413), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(G169), .ZN(new_n420));
  AOI21_X1  g0220(.A(KEYINPUT81), .B1(new_n409), .B2(new_n263), .ZN(new_n421));
  AND2_X1   g0221(.A1(new_n417), .A2(new_n254), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n423), .A2(G179), .A3(new_n413), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n408), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT18), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT18), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n408), .A2(new_n425), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT17), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n404), .A2(new_n407), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n412), .A2(G190), .A3(new_n413), .A4(new_n418), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n360), .B1(new_n423), .B2(new_n413), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n430), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n409), .A2(KEYINPUT81), .A3(new_n263), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n437), .A2(new_n421), .A3(new_n422), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n432), .B1(new_n438), .B2(new_n360), .ZN(new_n439));
  NOR3_X1   g0239(.A1(new_n408), .A2(new_n439), .A3(KEYINPUT17), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n427), .B(new_n429), .C1(new_n436), .C2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n331), .A2(new_n377), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n274), .A2(G33), .ZN(new_n445));
  AND3_X1   g0245(.A1(new_n308), .A2(new_n275), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(KEYINPUT25), .B1(new_n276), .B2(new_n298), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n276), .A2(KEYINPUT25), .A3(new_n298), .ZN(new_n449));
  AOI22_X1  g0249(.A1(G107), .A2(new_n446), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT87), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n379), .A2(new_n381), .A3(new_n223), .A4(G87), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT22), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT22), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n247), .A2(new_n454), .A3(new_n223), .A4(G87), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G33), .A2(G116), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(G20), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT23), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n459), .B1(new_n223), .B2(G107), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n298), .A2(KEYINPUT23), .A3(G20), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n458), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n456), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT24), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT24), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n456), .A2(new_n465), .A3(new_n462), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n451), .B1(new_n467), .B2(new_n280), .ZN(new_n468));
  AND3_X1   g0268(.A1(new_n456), .A2(new_n465), .A3(new_n462), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n465), .B1(new_n456), .B2(new_n462), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n451), .B(new_n280), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n450), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n254), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n379), .A2(new_n381), .A3(G257), .A4(G1698), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT88), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT88), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n247), .A2(new_n477), .A3(G257), .A4(G1698), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n379), .A2(new_n381), .A3(G250), .A4(new_n248), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G294), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n474), .B1(new_n484), .B2(KEYINPUT89), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n482), .B1(new_n476), .B2(new_n478), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT89), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G41), .ZN(new_n489));
  OR2_X1    g0289(.A1(new_n489), .A2(KEYINPUT5), .ZN(new_n490));
  INV_X1    g0290(.A(G45), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(G1), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n489), .A2(KEYINPUT5), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n490), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n260), .A2(new_n494), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n485), .A2(new_n488), .B1(G264), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(G179), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n260), .A2(G274), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n490), .A2(KEYINPUT83), .A3(new_n492), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n274), .B(G45), .C1(new_n489), .C2(KEYINPUT5), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT83), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n500), .A2(new_n503), .A3(new_n493), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n499), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n496), .A2(new_n497), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n484), .A2(KEYINPUT89), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n508), .A2(new_n254), .A3(new_n488), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n495), .A2(G264), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n509), .A2(new_n506), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n294), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n473), .A2(new_n507), .A3(new_n512), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n499), .A2(new_n505), .B1(new_n495), .B2(G257), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n379), .A2(new_n381), .A3(G244), .A4(new_n248), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT4), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n247), .A2(KEYINPUT4), .A3(G244), .A4(new_n248), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G283), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n247), .A2(G250), .A3(G1698), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n517), .A2(new_n518), .A3(new_n519), .A4(new_n520), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n521), .A2(KEYINPUT82), .A3(new_n254), .ZN(new_n522));
  AOI21_X1  g0322(.A(KEYINPUT82), .B1(new_n521), .B2(new_n254), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n497), .B(new_n514), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n275), .A2(G97), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n308), .A2(new_n275), .A3(new_n445), .ZN(new_n527));
  INV_X1    g0327(.A(G97), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT6), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n244), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n298), .A2(KEYINPUT6), .A3(G97), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n533), .A2(G20), .B1(G77), .B2(new_n287), .ZN(new_n534));
  OAI21_X1  g0334(.A(G107), .B1(new_n383), .B2(new_n385), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n529), .B1(new_n536), .B2(new_n280), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n521), .A2(new_n254), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n514), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n537), .B1(new_n294), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n514), .A2(G190), .A3(new_n538), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n541), .A2(new_n537), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n514), .B1(new_n522), .B2(new_n523), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G200), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n524), .A2(new_n540), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n446), .A2(G116), .ZN(new_n546));
  INV_X1    g0346(.A(G116), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n276), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n519), .B(new_n223), .C1(G33), .C2(new_n528), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT86), .ZN(new_n550));
  XNOR2_X1  g0350(.A(new_n549), .B(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n308), .B1(G20), .B2(new_n547), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n551), .A2(KEYINPUT20), .A3(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(KEYINPUT20), .B1(new_n551), .B2(new_n552), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n546), .B(new_n548), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n247), .A2(G264), .A3(G1698), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n382), .A2(G303), .ZN(new_n558));
  INV_X1    g0358(.A(G257), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n557), .B(new_n558), .C1(new_n299), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n254), .ZN(new_n561));
  INV_X1    g0361(.A(G270), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n260), .A2(new_n494), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n561), .B(new_n506), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n556), .A2(KEYINPUT21), .A3(G169), .A4(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT21), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n546), .A2(new_n548), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n551), .A2(new_n552), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT20), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n567), .B1(new_n570), .B2(new_n553), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n560), .A2(new_n254), .ZN(new_n572));
  OAI22_X1  g0372(.A1(new_n504), .A2(new_n498), .B1(new_n563), .B2(new_n562), .ZN(new_n573));
  OAI21_X1  g0373(.A(G169), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n566), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n572), .A2(new_n573), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n556), .A2(G179), .A3(new_n576), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n565), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n556), .B1(G190), .B2(new_n576), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(new_n360), .B2(new_n576), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n513), .A2(new_n545), .A3(new_n578), .A4(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n509), .A2(new_n321), .A3(new_n506), .A4(new_n510), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT90), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n582), .A2(new_n583), .B1(new_n511), .B2(new_n360), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n496), .A2(KEYINPUT90), .A3(new_n321), .A4(new_n506), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n473), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n247), .A2(new_n223), .A3(G68), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT19), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n223), .B1(new_n334), .B2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(G87), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n590), .A2(new_n528), .A3(new_n298), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n588), .B1(new_n289), .B2(new_n528), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n587), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n280), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n311), .A2(new_n276), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n595), .B(new_n596), .C1(new_n311), .C2(new_n527), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n379), .A2(new_n381), .A3(G238), .A4(new_n248), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n379), .A2(new_n381), .A3(G244), .A4(G1698), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n598), .A2(new_n599), .A3(new_n457), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n254), .ZN(new_n601));
  NOR3_X1   g0401(.A1(new_n491), .A2(G1), .A3(G274), .ZN(new_n602));
  AOI21_X1  g0402(.A(G250), .B1(new_n274), .B2(G45), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n260), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT84), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT84), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n601), .A2(new_n608), .A3(new_n605), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n294), .A3(new_n609), .ZN(new_n610));
  AOI221_X4 g0410(.A(KEYINPUT84), .B1(new_n260), .B2(new_n604), .C1(new_n600), .C2(new_n254), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n608), .B1(new_n601), .B2(new_n605), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n497), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n610), .A2(new_n613), .A3(KEYINPUT85), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT85), .B1(new_n610), .B2(new_n613), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n597), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(G190), .B1(new_n611), .B2(new_n612), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n446), .A2(G87), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n595), .A2(new_n596), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n607), .A2(new_n609), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n617), .B(new_n619), .C1(new_n620), .C2(new_n318), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n581), .A2(new_n586), .A3(new_n622), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n444), .A2(new_n623), .ZN(G372));
  INV_X1    g0424(.A(new_n606), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n613), .B(new_n597), .C1(G169), .C2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT91), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n619), .B(new_n628), .C1(new_n318), .C2(new_n625), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n595), .A2(new_n596), .A3(new_n618), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n318), .B1(new_n601), .B2(new_n605), .ZN(new_n631));
  OAI21_X1  g0431(.A(KEYINPUT91), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n629), .A2(new_n617), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n626), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n536), .A2(new_n280), .ZN(new_n635));
  INV_X1    g0435(.A(new_n529), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n538), .ZN(new_n638));
  OAI22_X1  g0438(.A1(new_n504), .A2(new_n498), .B1(new_n563), .B2(new_n559), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n294), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n524), .A2(new_n637), .A3(new_n640), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n634), .A2(KEYINPUT26), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n641), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n616), .A2(new_n621), .A3(new_n643), .ZN(new_n644));
  AOI211_X1 g0444(.A(new_n627), .B(new_n642), .C1(KEYINPUT26), .C2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n513), .A2(new_n578), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n582), .A2(new_n583), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n511), .A2(new_n360), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(new_n585), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n473), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT82), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n538), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n521), .A2(KEYINPUT82), .A3(new_n254), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n360), .B1(new_n655), .B2(new_n514), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n541), .A2(new_n537), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n641), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n658), .A2(new_n634), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n646), .A2(new_n651), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n645), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n444), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n427), .A2(new_n429), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n362), .A2(new_n364), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n375), .B1(new_n664), .B2(new_n317), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n431), .A2(new_n435), .A3(new_n430), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n419), .A2(G200), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n404), .A2(new_n667), .A3(new_n407), .A4(new_n432), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(KEYINPUT17), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n663), .B1(new_n665), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n329), .A2(new_n330), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n296), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n662), .A2(new_n674), .ZN(G369));
  AND2_X1   g0475(.A1(new_n223), .A2(G13), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n274), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(G213), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n513), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n586), .B1(new_n473), .B2(new_n682), .ZN(new_n685));
  INV_X1    g0485(.A(new_n513), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n565), .A2(new_n575), .A3(new_n577), .ZN(new_n688));
  INV_X1    g0488(.A(new_n682), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT92), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n684), .B1(new_n687), .B2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n687), .A2(new_n683), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n556), .A2(new_n682), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n688), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n688), .A2(new_n695), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(new_n580), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(G330), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n694), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n693), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT93), .ZN(G399));
  INV_X1    g0503(.A(new_n210), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(G41), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n591), .A2(G116), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n705), .A2(new_n274), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n708), .B1(new_n227), .B2(new_n705), .ZN(new_n709));
  XOR2_X1   g0509(.A(new_n709), .B(KEYINPUT28), .Z(new_n710));
  AOI21_X1  g0510(.A(new_n682), .B1(new_n645), .B2(new_n660), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(KEYINPUT29), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n660), .A2(new_n626), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT26), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n634), .A2(new_n714), .A3(new_n641), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n644), .A2(new_n714), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n715), .B1(new_n716), .B2(KEYINPUT98), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT98), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n644), .A2(new_n718), .A3(new_n714), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n713), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(KEYINPUT99), .B1(new_n720), .B2(new_n682), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT99), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n644), .A2(new_n718), .A3(new_n714), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n718), .B1(new_n644), .B2(new_n714), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n723), .A2(new_n724), .A3(new_n715), .ZN(new_n725));
  OAI211_X1 g0525(.A(new_n722), .B(new_n689), .C1(new_n725), .C2(new_n713), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n721), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n712), .B1(new_n727), .B2(KEYINPUT29), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT94), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n254), .B1(new_n486), .B2(new_n487), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n484), .A2(KEYINPUT89), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n510), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n611), .A2(new_n612), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n729), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n496), .A2(KEYINPUT94), .A3(new_n620), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n539), .A2(new_n564), .A3(new_n497), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n734), .A2(new_n735), .A3(KEYINPUT30), .A4(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(KEYINPUT95), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n576), .A2(G179), .A3(new_n514), .A4(new_n538), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n620), .A2(new_n509), .A3(new_n510), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n739), .B1(new_n729), .B2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT95), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n741), .A2(new_n742), .A3(KEYINPUT30), .A4(new_n735), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n738), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT30), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT96), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n576), .A2(G179), .A3(new_n625), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n750), .A2(new_n511), .A3(new_n543), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n745), .A2(KEYINPUT96), .A3(new_n746), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n744), .A2(new_n749), .A3(new_n751), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n682), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT97), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT31), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  AND3_X1   g0557(.A1(new_n745), .A2(KEYINPUT96), .A3(new_n746), .ZN(new_n758));
  AOI21_X1  g0558(.A(KEYINPUT96), .B1(new_n745), .B2(new_n746), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n751), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n761), .B1(new_n738), .B2(new_n743), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n689), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(KEYINPUT97), .B1(new_n763), .B2(KEYINPUT31), .ZN(new_n764));
  NOR4_X1   g0564(.A1(new_n581), .A2(new_n622), .A3(new_n586), .A4(new_n682), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n762), .A2(new_n747), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n689), .A2(new_n756), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n757), .A2(new_n764), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n728), .B1(G330), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n710), .B1(new_n770), .B2(G1), .ZN(G364));
  NOR2_X1   g0571(.A1(new_n223), .A2(G190), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n772), .A2(new_n497), .A3(new_n360), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n773), .A2(KEYINPUT101), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(KEYINPUT101), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G159), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT32), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n321), .A2(G179), .A3(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n223), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n528), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n497), .A2(new_n360), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(new_n772), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n382), .B(new_n782), .C1(G68), .C2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n223), .A2(new_n497), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n787), .A2(new_n321), .A3(new_n360), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n223), .A2(new_n321), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n783), .A2(new_n789), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n788), .A2(new_n202), .B1(new_n790), .B2(new_n277), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n787), .A2(G190), .A3(new_n360), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n791), .B1(G58), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n319), .A2(new_n497), .A3(new_n772), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G107), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n319), .A2(new_n497), .A3(new_n789), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G87), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n786), .A2(new_n794), .A3(new_n797), .A4(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n788), .ZN(new_n802));
  INV_X1    g0602(.A(new_n790), .ZN(new_n803));
  AOI22_X1  g0603(.A1(G311), .A2(new_n802), .B1(new_n803), .B2(G326), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n247), .B1(new_n793), .B2(G322), .ZN(new_n805));
  INV_X1    g0605(.A(G317), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(KEYINPUT33), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n806), .A2(KEYINPUT33), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n785), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n781), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(G294), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n804), .A2(new_n805), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n777), .A2(G329), .B1(G303), .B2(new_n799), .ZN(new_n813));
  INV_X1    g0613(.A(G283), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n814), .B2(new_n795), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n779), .A2(new_n801), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n222), .B1(G20), .B2(new_n294), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(G13), .A2(G33), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n820), .A2(G20), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(new_n817), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n210), .A2(new_n247), .ZN(new_n823));
  INV_X1    g0623(.A(G355), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n823), .A2(new_n824), .B1(G116), .B2(new_n210), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT100), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n242), .A2(new_n491), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n704), .A2(new_n247), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(G45), .B2(new_n226), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n827), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n825), .A2(new_n826), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n822), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n274), .B1(new_n676), .B2(G45), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n705), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n818), .A2(new_n833), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(new_n698), .B2(new_n821), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n700), .A2(new_n836), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n698), .A2(new_n699), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(G396));
  OAI21_X1  g0642(.A(new_n322), .B1(new_n314), .B2(new_n689), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n317), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n317), .A2(new_n682), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n711), .B(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n769), .A2(G330), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n836), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n850), .B2(new_n849), .ZN(new_n852));
  INV_X1    g0652(.A(new_n836), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n817), .A2(new_n819), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(KEYINPUT102), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n853), .B1(new_n856), .B2(new_n202), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n795), .A2(new_n590), .ZN(new_n858));
  OR2_X1    g0658(.A1(new_n785), .A2(KEYINPUT103), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n785), .A2(KEYINPUT103), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n858), .B1(new_n862), .B2(G283), .ZN(new_n863));
  INV_X1    g0663(.A(G311), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n863), .B1(new_n298), .B2(new_n798), .C1(new_n864), .C2(new_n776), .ZN(new_n865));
  INV_X1    g0665(.A(G303), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n382), .B1(new_n790), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(G294), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n792), .A2(new_n868), .B1(new_n788), .B2(new_n547), .ZN(new_n869));
  NOR4_X1   g0669(.A1(new_n865), .A2(new_n782), .A3(new_n867), .A4(new_n869), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n793), .A2(G143), .B1(new_n785), .B2(G150), .ZN(new_n871));
  INV_X1    g0671(.A(G137), .ZN(new_n872));
  INV_X1    g0672(.A(G159), .ZN(new_n873));
  OAI221_X1 g0673(.A(new_n871), .B1(new_n872), .B2(new_n790), .C1(new_n873), .C2(new_n788), .ZN(new_n874));
  XOR2_X1   g0674(.A(KEYINPUT104), .B(KEYINPUT34), .Z(new_n875));
  XNOR2_X1  g0675(.A(new_n874), .B(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n796), .A2(G68), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n877), .B1(new_n277), .B2(new_n798), .C1(new_n388), .C2(new_n781), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(G132), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n247), .B1(new_n776), .B2(new_n880), .ZN(new_n881));
  XOR2_X1   g0681(.A(new_n881), .B(KEYINPUT105), .Z(new_n882));
  AOI21_X1  g0682(.A(new_n870), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n817), .ZN(new_n884));
  OAI221_X1 g0684(.A(new_n857), .B1(new_n883), .B2(new_n884), .C1(new_n848), .C2(new_n820), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n852), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(G384));
  OAI211_X1 g0687(.A(G116), .B(new_n224), .C1(new_n533), .C2(KEYINPUT35), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n888), .B1(KEYINPUT35), .B2(new_n533), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n889), .B(KEYINPUT36), .ZN(new_n890));
  OR3_X1    g0690(.A1(new_n226), .A2(new_n202), .A3(new_n389), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n201), .A2(G68), .ZN(new_n892));
  AOI211_X1 g0692(.A(new_n274), .B(G13), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n369), .A2(new_n682), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n376), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n365), .A2(new_n375), .A3(new_n895), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n623), .A2(new_n689), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n763), .B2(KEYINPUT31), .ZN(new_n901));
  AOI211_X1 g0701(.A(new_n756), .B(new_n689), .C1(new_n760), .C2(new_n762), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n848), .B(new_n899), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT38), .ZN(new_n905));
  INV_X1    g0705(.A(new_n680), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n408), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n442), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT37), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT108), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n909), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n426), .A2(new_n907), .A3(new_n668), .ZN(new_n912));
  XOR2_X1   g0712(.A(new_n911), .B(new_n912), .Z(new_n913));
  OAI21_X1  g0713(.A(new_n905), .B1(new_n908), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n308), .B1(new_n394), .B2(new_n400), .ZN(new_n915));
  INV_X1    g0715(.A(new_n406), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n917), .A2(new_n680), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n436), .A2(new_n440), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n918), .B1(new_n919), .B2(new_n663), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(KEYINPUT106), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT107), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n420), .A2(new_n424), .A3(new_n680), .ZN(new_n923));
  INV_X1    g0723(.A(new_n917), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n431), .A2(new_n435), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n922), .B1(new_n925), .B2(new_n909), .ZN(new_n926));
  INV_X1    g0726(.A(new_n923), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n668), .B1(new_n927), .B2(new_n917), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n928), .A2(KEYINPUT107), .A3(KEYINPUT37), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n926), .B(new_n929), .C1(KEYINPUT37), .C2(new_n912), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT106), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n441), .A2(new_n931), .A3(new_n918), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n921), .A2(new_n930), .A3(KEYINPUT38), .A4(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n914), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n904), .A2(KEYINPUT40), .A3(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT40), .ZN(new_n936));
  INV_X1    g0736(.A(new_n918), .ZN(new_n937));
  AND3_X1   g0737(.A1(new_n408), .A2(new_n425), .A3(new_n428), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n428), .B1(new_n408), .B2(new_n425), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI211_X1 g0740(.A(KEYINPUT106), .B(new_n937), .C1(new_n940), .C2(new_n670), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n931), .B1(new_n441), .B2(new_n918), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(KEYINPUT38), .B1(new_n943), .B2(new_n930), .ZN(new_n944));
  AND4_X1   g0744(.A1(KEYINPUT38), .A2(new_n921), .A3(new_n930), .A4(new_n932), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n936), .B1(new_n946), .B2(new_n903), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n947), .A2(KEYINPUT110), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT110), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n921), .A2(new_n930), .A3(new_n932), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n905), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n933), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n765), .B1(new_n754), .B2(new_n756), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n763), .A2(KEYINPUT31), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n847), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n952), .A2(new_n955), .A3(new_n899), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n949), .B1(new_n956), .B2(new_n936), .ZN(new_n957));
  OAI211_X1 g0757(.A(G330), .B(new_n935), .C1(new_n948), .C2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n754), .A2(new_n756), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n959), .A2(new_n954), .A3(new_n900), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n444), .A2(G330), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT111), .Z(new_n963));
  AND3_X1   g0763(.A1(new_n904), .A2(KEYINPUT40), .A3(new_n934), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n947), .A2(KEYINPUT110), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n956), .A2(new_n949), .A3(new_n936), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n967), .A2(new_n444), .A3(new_n960), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n963), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n952), .A2(KEYINPUT39), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT39), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n914), .A2(new_n933), .A3(new_n971), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n375), .A2(new_n682), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n845), .B1(new_n711), .B2(new_n848), .ZN(new_n978));
  INV_X1    g0778(.A(new_n898), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(new_n376), .B2(new_n896), .ZN(new_n980));
  NOR3_X1   g0780(.A1(new_n946), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(new_n663), .B2(new_n680), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n977), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n969), .B(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n674), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n727), .A2(KEYINPUT29), .ZN(new_n986));
  INV_X1    g0786(.A(new_n712), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n986), .A2(new_n444), .A3(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT109), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n728), .A2(KEYINPUT109), .A3(new_n444), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n985), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n984), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n274), .B2(new_n676), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n984), .A2(new_n992), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n894), .B1(new_n994), .B2(new_n995), .ZN(G367));
  INV_X1    g0796(.A(new_n829), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n822), .B1(new_n210), .B2(new_n311), .C1(new_n997), .C2(new_n237), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n836), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n777), .A2(G137), .B1(G58), .B2(new_n799), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n1000), .B1(new_n202), .B2(new_n795), .C1(new_n873), .C2(new_n861), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n284), .A2(new_n802), .B1(new_n803), .B2(G143), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n810), .A2(G68), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n382), .B1(new_n793), .B2(G150), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n792), .A2(new_n866), .B1(new_n788), .B2(new_n814), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n247), .B(new_n1006), .C1(G311), .C2(new_n803), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n799), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT46), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n798), .B2(new_n547), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n810), .A2(G107), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1007), .A2(new_n1008), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n796), .A2(G97), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n776), .B2(new_n806), .C1(new_n861), .C2(new_n868), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n1001), .A2(new_n1005), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT47), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n884), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n999), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n821), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n689), .A2(new_n619), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n634), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n627), .A2(new_n1021), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1019), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n545), .B1(new_n537), .B2(new_n689), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n643), .A2(new_n682), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n684), .B(new_n1028), .C1(new_n687), .C2(new_n691), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT45), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1029), .B(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1028), .ZN(new_n1032));
  AOI21_X1  g0832(.A(KEYINPUT44), .B1(new_n692), .B2(new_n1032), .ZN(new_n1033));
  AND3_X1   g0833(.A1(new_n692), .A2(KEYINPUT44), .A3(new_n1032), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1031), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT112), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n701), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n701), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1035), .A2(new_n1036), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n691), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n694), .B(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(new_n700), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n770), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n770), .B1(new_n1041), .B2(new_n1045), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n705), .B(KEYINPUT41), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n835), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n694), .A2(new_n1042), .A3(new_n1028), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1049), .A2(KEYINPUT42), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n686), .B1(new_n656), .B2(new_n657), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n682), .B1(new_n1051), .B2(new_n641), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n1049), .B2(KEYINPUT42), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n1050), .A2(new_n1053), .B1(KEYINPUT43), .B2(new_n1024), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n1024), .A2(KEYINPUT43), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n701), .A2(new_n1032), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1059));
  AND3_X1   g0859(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1058), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1025), .B1(new_n1048), .B2(new_n1063), .ZN(G387));
  NAND2_X1  g0864(.A1(new_n1044), .A2(new_n835), .ZN(new_n1065));
  AOI211_X1 g0865(.A(G45), .B(new_n707), .C1(G68), .C2(G77), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n1066), .A2(KEYINPUT113), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(KEYINPUT113), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n309), .A2(new_n277), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT50), .Z(new_n1070));
  NAND3_X1  g0870(.A1(new_n1067), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1071), .B(new_n829), .C1(new_n234), .C2(new_n491), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1072), .B1(G107), .B2(new_n210), .C1(new_n706), .C2(new_n823), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n853), .B1(new_n1073), .B2(new_n822), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n799), .A2(G77), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1013), .B(new_n1075), .C1(new_n286), .C2(new_n776), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n247), .B1(new_n788), .B2(new_n349), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n792), .A2(new_n277), .B1(new_n790), .B2(new_n873), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n291), .A2(new_n784), .B1(new_n311), .B2(new_n781), .ZN(new_n1079));
  NOR4_X1   g0879(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n798), .A2(new_n868), .B1(new_n814), .B2(new_n781), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(G303), .A2(new_n802), .B1(new_n803), .B2(G322), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n806), .B2(new_n792), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(G311), .B2(new_n862), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1081), .B1(new_n1084), .B2(KEYINPUT48), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT114), .Z(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(KEYINPUT48), .B2(new_n1084), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT49), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n247), .B1(new_n777), .B2(G326), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n547), .B2(new_n795), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1080), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n1074), .B1(new_n694), .B2(new_n1020), .C1(new_n1093), .C2(new_n884), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1045), .A2(new_n705), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n770), .A2(new_n1044), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1065), .B(new_n1094), .C1(new_n1095), .C2(new_n1096), .ZN(G393));
  AOI22_X1  g0897(.A1(new_n862), .A2(G303), .B1(new_n777), .B2(G322), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n814), .B2(new_n798), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n792), .A2(new_n864), .B1(new_n790), .B2(new_n806), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT52), .Z(new_n1101));
  AOI21_X1  g0901(.A(new_n247), .B1(new_n802), .B2(G294), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n797), .B(new_n1102), .C1(new_n547), .C2(new_n781), .ZN(new_n1103));
  NOR3_X1   g0903(.A1(new_n1099), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n793), .A2(G159), .B1(new_n803), .B2(G150), .ZN(new_n1105));
  XOR2_X1   g0905(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n1106));
  AOI22_X1  g0906(.A1(new_n777), .A2(G143), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n861), .A2(new_n201), .B1(new_n349), .B2(new_n798), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n382), .B1(new_n802), .B2(new_n309), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n202), .B2(new_n781), .ZN(new_n1111));
  NOR4_X1   g0911(.A1(new_n1108), .A2(new_n1109), .A3(new_n858), .A4(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n817), .B1(new_n1104), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n822), .B1(new_n210), .B2(new_n528), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n829), .B2(new_n245), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n836), .B1(new_n1115), .B2(KEYINPUT115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(KEYINPUT115), .B2(new_n1115), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1113), .B(new_n1117), .C1(new_n1028), .C2(new_n1020), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1035), .B(new_n1039), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n705), .B1(new_n1041), .B2(new_n1045), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n1119), .A2(new_n1045), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n1118), .B1(new_n834), .B2(new_n1119), .C1(new_n1120), .C2(new_n1121), .ZN(G390));
  AOI21_X1  g0922(.A(new_n853), .B1(new_n856), .B2(new_n291), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n862), .A2(G107), .B1(new_n777), .B2(G294), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n382), .B1(new_n790), .B2(new_n814), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n792), .A2(new_n547), .B1(new_n788), .B2(new_n528), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n1125), .B(new_n1126), .C1(G77), .C2(new_n810), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1124), .A2(new_n800), .A3(new_n877), .A4(new_n1127), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n798), .A2(new_n286), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT53), .ZN(new_n1130));
  INV_X1    g0930(.A(G128), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n792), .A2(new_n880), .B1(new_n790), .B2(new_n1131), .ZN(new_n1132));
  XOR2_X1   g0932(.A(KEYINPUT54), .B(G143), .Z(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n247), .B1(new_n1134), .B2(new_n788), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n1132), .B(new_n1135), .C1(G159), .C2(new_n810), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n862), .A2(G137), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n777), .A2(G125), .B1(new_n284), .B2(new_n796), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1130), .A2(new_n1136), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  AND2_X1   g0939(.A1(new_n1128), .A2(new_n1139), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n1123), .B1(new_n884), .B2(new_n1140), .C1(new_n974), .C2(new_n820), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n721), .A2(new_n726), .A3(new_n846), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT117), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n980), .B(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1142), .A2(new_n1144), .A3(new_n844), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n976), .B1(new_n914), .B2(new_n933), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n769), .A2(G330), .A3(new_n848), .A4(new_n899), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n975), .B1(new_n978), .B2(new_n980), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1149), .A2(new_n970), .A3(new_n972), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1147), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n973), .A2(new_n1149), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n904), .A2(G330), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1151), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1141), .B1(new_n1154), .B2(new_n834), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n705), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n990), .A2(new_n991), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n960), .A2(G330), .A3(new_n848), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n980), .B(KEYINPUT117), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1142), .A2(new_n844), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1160), .A2(new_n1161), .A3(new_n1148), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n769), .A2(G330), .A3(new_n848), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n980), .A2(new_n1163), .B1(new_n904), .B2(G330), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1162), .B1(new_n1164), .B2(new_n978), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1157), .A2(new_n1165), .A3(new_n674), .A4(new_n961), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1156), .B1(new_n1166), .B2(new_n1154), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1153), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(new_n1148), .B2(new_n1152), .ZN(new_n1169));
  AOI21_X1  g0969(.A(KEYINPUT109), .B1(new_n728), .B2(new_n444), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT29), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(new_n721), .B2(new_n726), .ZN(new_n1172));
  NOR4_X1   g0972(.A1(new_n1172), .A2(new_n989), .A3(new_n443), .A4(new_n712), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n674), .B(new_n961), .C1(new_n1170), .C2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1169), .A2(new_n1175), .A3(new_n1165), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1155), .B1(new_n1167), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(G378));
  NAND2_X1  g0978(.A1(new_n977), .A2(new_n982), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n296), .ZN(new_n1182));
  AOI21_X1  g0982(.A(KEYINPUT121), .B1(new_n673), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n293), .A2(new_n680), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n673), .A2(KEYINPUT121), .A3(new_n1182), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1184), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1186), .B1(new_n1184), .B2(new_n1187), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1181), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1190), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1192), .A2(new_n1180), .A3(new_n1188), .ZN(new_n1193));
  AND2_X1   g0993(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n958), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(new_n967), .B2(G330), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1179), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n958), .A2(new_n1194), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n967), .A2(G330), .A3(new_n1196), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n983), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1198), .A2(new_n835), .A3(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n853), .B1(new_n856), .B2(new_n201), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n247), .A2(G41), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(G33), .A2(G41), .ZN(new_n1205));
  OR3_X1    g1005(.A1(new_n1204), .A2(G50), .A3(new_n1205), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n777), .A2(G283), .B1(G58), .B2(new_n796), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n792), .A2(new_n298), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT118), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1207), .A2(new_n1075), .A3(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n781), .A2(new_n349), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n790), .A2(new_n547), .B1(new_n784), .B2(new_n528), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1204), .B1(new_n311), .B2(new_n788), .ZN(new_n1213));
  NOR4_X1   g1013(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1206), .B1(new_n1214), .B2(KEYINPUT58), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1215), .A2(KEYINPUT119), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n793), .A2(G128), .B1(new_n802), .B2(G137), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(G125), .A2(new_n803), .B1(new_n785), .B2(G132), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1219), .B1(new_n286), .B2(new_n781), .C1(new_n798), .C2(new_n1134), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1222));
  OR2_X1    g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(G124), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1205), .B1(new_n795), .B2(new_n873), .C1(new_n776), .C2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1223), .A2(new_n1226), .B1(KEYINPUT58), .B2(new_n1214), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1216), .A2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(KEYINPUT119), .B2(new_n1215), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1203), .B1(new_n884), .B2(new_n1229), .C1(new_n1194), .C2(new_n820), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n1202), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1163), .A2(new_n980), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n1153), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n978), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n1159), .A2(new_n1158), .B1(new_n1142), .B2(new_n844), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1233), .A2(new_n1234), .B1(new_n1235), .B2(new_n1148), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1175), .B1(new_n1154), .B2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1198), .A2(new_n1201), .A3(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT57), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1198), .A2(KEYINPUT57), .A3(new_n1201), .A4(new_n1237), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n705), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1231), .B1(new_n1240), .B2(new_n1242), .ZN(G375));
  NAND2_X1  g1043(.A1(new_n1174), .A2(new_n1236), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1166), .A2(new_n1244), .A3(new_n1047), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1159), .A2(new_n819), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n836), .B1(new_n855), .B2(G68), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n861), .A2(new_n547), .B1(new_n776), .B2(new_n866), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n793), .A2(G283), .B1(new_n803), .B2(G294), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1249), .B(new_n382), .C1(new_n298), .C2(new_n788), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n781), .A2(new_n311), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n202), .A2(new_n795), .B1(new_n798), .B2(new_n528), .ZN(new_n1252));
  NOR4_X1   g1052(.A1(new_n1248), .A2(new_n1250), .A3(new_n1251), .A4(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  OR2_X1    g1054(.A1(new_n1254), .A2(KEYINPUT122), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n862), .A2(new_n1133), .B1(G58), .B2(new_n796), .ZN(new_n1256));
  OAI221_X1 g1056(.A(new_n247), .B1(new_n788), .B2(new_n286), .C1(new_n872), .C2(new_n792), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(G50), .B2(new_n810), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n803), .A2(G132), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1259), .B(KEYINPUT123), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n777), .A2(G128), .B1(G159), .B2(new_n799), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1256), .A2(new_n1258), .A3(new_n1260), .A4(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1254), .A2(KEYINPUT122), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1255), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1247), .B1(new_n1264), .B2(new_n817), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n1165), .A2(new_n835), .B1(new_n1246), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1245), .A2(new_n1266), .ZN(G381));
  INV_X1    g1067(.A(G390), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n886), .ZN(new_n1269));
  OR2_X1    g1069(.A1(G393), .A2(G396), .ZN(new_n1270));
  NOR4_X1   g1070(.A1(new_n1269), .A2(G381), .A3(G387), .A4(new_n1270), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(new_n1271), .B(KEYINPUT124), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1202), .A2(new_n1230), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1241), .A2(new_n705), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1273), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1272), .A2(new_n1177), .A3(new_n1276), .ZN(G407));
  NAND3_X1  g1077(.A1(new_n1276), .A2(new_n681), .A3(new_n1177), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(G407), .A2(G213), .A3(new_n1278), .ZN(G409));
  NAND4_X1  g1079(.A1(new_n1198), .A2(new_n1047), .A3(new_n1201), .A4(new_n1237), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1280), .A2(new_n1177), .A3(new_n1202), .A4(new_n1230), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n681), .A2(G213), .ZN(new_n1282));
  AND2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1283), .B1(new_n1276), .B2(new_n1177), .ZN(new_n1284));
  OAI21_X1  g1084(.A(KEYINPUT60), .B1(new_n1174), .B2(new_n1236), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1156), .B1(new_n1285), .B2(new_n1244), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT125), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1174), .A2(KEYINPUT60), .A3(new_n1236), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1286), .A2(new_n1287), .A3(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1287), .B1(new_n1286), .B2(new_n1288), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1266), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n886), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1285), .A2(new_n1244), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1293), .A2(new_n705), .A3(new_n1288), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(KEYINPUT125), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1286), .A2(new_n1287), .A3(new_n1288), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1297), .A2(G384), .A3(new_n1266), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1292), .A2(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(KEYINPUT62), .B1(new_n1284), .B2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n681), .A2(G213), .A3(G2897), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(G384), .B1(new_n1297), .B2(new_n1266), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1266), .ZN(new_n1304));
  AOI211_X1 g1104(.A(new_n886), .B(new_n1304), .C1(new_n1295), .C2(new_n1296), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1302), .B1(new_n1303), .B2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1292), .A2(new_n1298), .A3(new_n1301), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1306), .A2(new_n1284), .A3(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT61), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1303), .A2(new_n1305), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1311), .B1(G375), .B2(G378), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT62), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1310), .A2(new_n1312), .A3(new_n1313), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1300), .A2(new_n1308), .A3(new_n1309), .A4(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(G393), .A2(G396), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1270), .A2(new_n1316), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(G387), .A2(new_n1268), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n770), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1040), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1039), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1319), .B1(new_n1322), .B2(new_n1044), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1047), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n834), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(new_n1062), .ZN(new_n1326));
  AOI21_X1  g1126(.A(G390), .B1(new_n1326), .B2(new_n1025), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1317), .B1(new_n1318), .B2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(G387), .A2(new_n1268), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1326), .A2(new_n1025), .A3(G390), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1329), .A2(new_n1330), .A3(new_n1270), .A4(new_n1316), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1328), .A2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1315), .A2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT126), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1308), .A2(new_n1334), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1328), .A2(new_n1309), .A3(new_n1331), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(G375), .A2(G378), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1337), .A2(new_n1292), .A3(new_n1298), .A4(new_n1283), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT63), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1336), .B1(new_n1338), .B2(new_n1339), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1310), .A2(new_n1312), .A3(KEYINPUT63), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1306), .A2(new_n1284), .A3(new_n1307), .A4(KEYINPUT126), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1335), .A2(new_n1340), .A3(new_n1341), .A4(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1333), .A2(new_n1343), .ZN(G405));
  NAND2_X1  g1144(.A1(new_n1299), .A2(KEYINPUT127), .ZN(new_n1345));
  OAI211_X1 g1145(.A(new_n1331), .B(new_n1328), .C1(new_n1299), .C2(KEYINPUT127), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT127), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1332), .A2(new_n1310), .A3(new_n1347), .ZN(new_n1348));
  XNOR2_X1  g1148(.A(G375), .B(new_n1177), .ZN(new_n1349));
  AND4_X1   g1149(.A1(new_n1345), .A2(new_n1346), .A3(new_n1348), .A4(new_n1349), .ZN(new_n1350));
  AOI22_X1  g1150(.A1(new_n1346), .A2(new_n1348), .B1(new_n1349), .B2(new_n1345), .ZN(new_n1351));
  NOR2_X1   g1151(.A1(new_n1350), .A2(new_n1351), .ZN(G402));
endmodule


