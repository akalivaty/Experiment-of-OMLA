

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U547 ( .A1(n536), .A2(n516), .ZN(n801) );
  OR2_X1 U548 ( .A1(n945), .A2(n639), .ZN(n640) );
  NOR2_X1 U549 ( .A1(n586), .A2(n512), .ZN(n596) );
  AND2_X2 U550 ( .A1(n524), .A2(G2105), .ZN(n590) );
  AND2_X1 U551 ( .A1(n526), .A2(G2104), .ZN(n587) );
  XNOR2_X1 U552 ( .A(KEYINPUT65), .B(KEYINPUT23), .ZN(n588) );
  INV_X1 U553 ( .A(KEYINPUT5), .ZN(n546) );
  NAND2_X1 U554 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U555 ( .A1(n679), .A2(n671), .ZN(n601) );
  INV_X1 U556 ( .A(KEYINPUT97), .ZN(n685) );
  NOR2_X1 U557 ( .A1(G164), .A2(G1384), .ZN(n727) );
  NOR2_X1 U558 ( .A1(G543), .A2(G651), .ZN(n800) );
  BUF_X1 U559 ( .A(n584), .Z(n894) );
  INV_X1 U560 ( .A(KEYINPUT66), .ZN(n593) );
  INV_X1 U561 ( .A(KEYINPUT100), .ZN(n742) );
  XNOR2_X1 U562 ( .A(n548), .B(n547), .ZN(n549) );
  INV_X1 U563 ( .A(G2104), .ZN(n524) );
  AND2_X1 U564 ( .A1(n887), .A2(G113), .ZN(n512) );
  NOR2_X1 U565 ( .A1(n708), .A2(n689), .ZN(n513) );
  INV_X1 U566 ( .A(KEYINPUT27), .ZN(n644) );
  XNOR2_X1 U567 ( .A(n645), .B(n644), .ZN(n646) );
  NOR2_X1 U568 ( .A1(G299), .A2(n651), .ZN(n648) );
  XNOR2_X1 U569 ( .A(n603), .B(KEYINPUT30), .ZN(n604) );
  INV_X1 U570 ( .A(KEYINPUT93), .ZN(n662) );
  INV_X1 U571 ( .A(KEYINPUT32), .ZN(n674) );
  AND2_X1 U572 ( .A1(n673), .A2(n672), .ZN(n675) );
  INV_X1 U573 ( .A(n727), .ZN(n599) );
  INV_X1 U574 ( .A(n643), .ZN(n642) );
  BUF_X1 U575 ( .A(n642), .Z(n665) );
  INV_X1 U576 ( .A(KEYINPUT12), .ZN(n614) );
  XNOR2_X1 U577 ( .A(n614), .B(KEYINPUT73), .ZN(n615) );
  NAND2_X1 U578 ( .A1(n526), .A2(n524), .ZN(n525) );
  XNOR2_X1 U579 ( .A(n616), .B(n615), .ZN(n618) );
  XNOR2_X1 U580 ( .A(n546), .B(KEYINPUT76), .ZN(n547) );
  XNOR2_X1 U581 ( .A(n594), .B(n593), .ZN(n595) );
  NAND2_X1 U582 ( .A1(n596), .A2(n595), .ZN(n598) );
  XNOR2_X1 U583 ( .A(n598), .B(n597), .ZN(n762) );
  NOR2_X1 U584 ( .A1(n532), .A2(n531), .ZN(G164) );
  NAND2_X1 U585 ( .A1(G91), .A2(n800), .ZN(n515) );
  XOR2_X1 U586 ( .A(KEYINPUT0), .B(G543), .Z(n536) );
  INV_X1 U587 ( .A(G651), .ZN(n516) );
  NAND2_X1 U588 ( .A1(G78), .A2(n801), .ZN(n514) );
  NAND2_X1 U589 ( .A1(n515), .A2(n514), .ZN(n521) );
  NOR2_X1 U590 ( .A1(G543), .A2(n516), .ZN(n518) );
  XNOR2_X1 U591 ( .A(KEYINPUT1), .B(KEYINPUT69), .ZN(n517) );
  XNOR2_X1 U592 ( .A(n518), .B(n517), .ZN(n804) );
  NAND2_X1 U593 ( .A1(n804), .A2(G65), .ZN(n519) );
  XOR2_X1 U594 ( .A(KEYINPUT70), .B(n519), .Z(n520) );
  NOR2_X1 U595 ( .A1(n521), .A2(n520), .ZN(n523) );
  NOR2_X2 U596 ( .A1(n536), .A2(G651), .ZN(n805) );
  NAND2_X1 U597 ( .A1(n805), .A2(G53), .ZN(n522) );
  NAND2_X1 U598 ( .A1(n523), .A2(n522), .ZN(G299) );
  XNOR2_X2 U599 ( .A(n525), .B(KEYINPUT17), .ZN(n584) );
  NAND2_X1 U600 ( .A1(G138), .A2(n584), .ZN(n528) );
  INV_X1 U601 ( .A(G2105), .ZN(n526) );
  BUF_X1 U602 ( .A(n587), .Z(n891) );
  NAND2_X1 U603 ( .A1(G102), .A2(n891), .ZN(n527) );
  NAND2_X1 U604 ( .A1(n528), .A2(n527), .ZN(n532) );
  NAND2_X1 U605 ( .A1(G126), .A2(n590), .ZN(n530) );
  AND2_X1 U606 ( .A1(G2104), .A2(G2105), .ZN(n887) );
  NAND2_X1 U607 ( .A1(G114), .A2(n887), .ZN(n529) );
  NAND2_X1 U608 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U609 ( .A1(G49), .A2(n805), .ZN(n534) );
  NAND2_X1 U610 ( .A1(G74), .A2(G651), .ZN(n533) );
  NAND2_X1 U611 ( .A1(n534), .A2(n533), .ZN(n535) );
  NOR2_X1 U612 ( .A1(n804), .A2(n535), .ZN(n538) );
  NAND2_X1 U613 ( .A1(n536), .A2(G87), .ZN(n537) );
  NAND2_X1 U614 ( .A1(n538), .A2(n537), .ZN(G288) );
  NAND2_X1 U615 ( .A1(n805), .A2(G51), .ZN(n539) );
  XOR2_X1 U616 ( .A(KEYINPUT77), .B(n539), .Z(n541) );
  NAND2_X1 U617 ( .A1(n804), .A2(G63), .ZN(n540) );
  NAND2_X1 U618 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U619 ( .A(KEYINPUT6), .B(n542), .ZN(n550) );
  NAND2_X1 U620 ( .A1(n800), .A2(G89), .ZN(n543) );
  XNOR2_X1 U621 ( .A(n543), .B(KEYINPUT4), .ZN(n545) );
  NAND2_X1 U622 ( .A1(G76), .A2(n801), .ZN(n544) );
  NAND2_X1 U623 ( .A1(n545), .A2(n544), .ZN(n548) );
  NOR2_X1 U624 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U625 ( .A(KEYINPUT7), .B(n551), .Z(G168) );
  NAND2_X1 U626 ( .A1(G64), .A2(n804), .ZN(n553) );
  NAND2_X1 U627 ( .A1(G52), .A2(n805), .ZN(n552) );
  NAND2_X1 U628 ( .A1(n553), .A2(n552), .ZN(n558) );
  NAND2_X1 U629 ( .A1(G90), .A2(n800), .ZN(n555) );
  NAND2_X1 U630 ( .A1(G77), .A2(n801), .ZN(n554) );
  NAND2_X1 U631 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U632 ( .A(KEYINPUT9), .B(n556), .Z(n557) );
  NOR2_X1 U633 ( .A1(n558), .A2(n557), .ZN(G171) );
  XOR2_X1 U634 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U635 ( .A1(G88), .A2(n800), .ZN(n560) );
  NAND2_X1 U636 ( .A1(G75), .A2(n801), .ZN(n559) );
  NAND2_X1 U637 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U638 ( .A(KEYINPUT82), .B(n561), .ZN(n565) );
  NAND2_X1 U639 ( .A1(G62), .A2(n804), .ZN(n563) );
  NAND2_X1 U640 ( .A1(G50), .A2(n805), .ZN(n562) );
  NAND2_X1 U641 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U642 ( .A1(n565), .A2(n564), .ZN(G166) );
  XNOR2_X1 U643 ( .A(KEYINPUT87), .B(G166), .ZN(G303) );
  XOR2_X1 U644 ( .A(KEYINPUT80), .B(KEYINPUT2), .Z(n567) );
  NAND2_X1 U645 ( .A1(G73), .A2(n801), .ZN(n566) );
  XNOR2_X1 U646 ( .A(n567), .B(n566), .ZN(n571) );
  NAND2_X1 U647 ( .A1(G86), .A2(n800), .ZN(n569) );
  NAND2_X1 U648 ( .A1(G61), .A2(n804), .ZN(n568) );
  NAND2_X1 U649 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U650 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U651 ( .A(KEYINPUT81), .B(n572), .Z(n574) );
  NAND2_X1 U652 ( .A1(n805), .A2(G48), .ZN(n573) );
  NAND2_X1 U653 ( .A1(n574), .A2(n573), .ZN(G305) );
  NAND2_X1 U654 ( .A1(G85), .A2(n800), .ZN(n576) );
  NAND2_X1 U655 ( .A1(G72), .A2(n801), .ZN(n575) );
  NAND2_X1 U656 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U657 ( .A(KEYINPUT68), .B(n577), .Z(n581) );
  NAND2_X1 U658 ( .A1(G60), .A2(n804), .ZN(n579) );
  NAND2_X1 U659 ( .A1(G47), .A2(n805), .ZN(n578) );
  AND2_X1 U660 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U661 ( .A1(n581), .A2(n580), .ZN(G290) );
  NOR2_X1 U662 ( .A1(G1976), .A2(G288), .ZN(n955) );
  INV_X1 U663 ( .A(n955), .ZN(n583) );
  INV_X1 U664 ( .A(KEYINPUT33), .ZN(n582) );
  AND2_X1 U665 ( .A1(n583), .A2(n582), .ZN(n688) );
  NAND2_X1 U666 ( .A1(n584), .A2(G137), .ZN(n585) );
  XNOR2_X1 U667 ( .A(n585), .B(KEYINPUT67), .ZN(n586) );
  NAND2_X1 U668 ( .A1(G101), .A2(n587), .ZN(n589) );
  XNOR2_X1 U669 ( .A(n589), .B(n588), .ZN(n592) );
  NAND2_X1 U670 ( .A1(G125), .A2(n590), .ZN(n591) );
  NAND2_X1 U671 ( .A1(n592), .A2(n591), .ZN(n594) );
  INV_X1 U672 ( .A(KEYINPUT64), .ZN(n597) );
  NAND2_X1 U673 ( .A1(n762), .A2(G40), .ZN(n726) );
  NOR2_X2 U674 ( .A1(n726), .A2(n599), .ZN(n643) );
  NOR2_X1 U675 ( .A1(G2084), .A2(n642), .ZN(n677) );
  INV_X1 U676 ( .A(n677), .ZN(n602) );
  INV_X1 U677 ( .A(G8), .ZN(n671) );
  NOR2_X1 U678 ( .A1(n671), .A2(G1966), .ZN(n600) );
  AND2_X1 U679 ( .A1(n642), .A2(n600), .ZN(n679) );
  NOR2_X1 U680 ( .A1(n604), .A2(G168), .ZN(n609) );
  INV_X1 U681 ( .A(G1961), .ZN(n949) );
  NAND2_X1 U682 ( .A1(n665), .A2(n949), .ZN(n607) );
  BUF_X1 U683 ( .A(n643), .Z(n605) );
  XNOR2_X1 U684 ( .A(KEYINPUT25), .B(G2078), .ZN(n1000) );
  NAND2_X1 U685 ( .A1(n605), .A2(n1000), .ZN(n606) );
  NAND2_X1 U686 ( .A1(n607), .A2(n606), .ZN(n657) );
  NOR2_X1 U687 ( .A1(G171), .A2(n657), .ZN(n608) );
  NOR2_X1 U688 ( .A1(n609), .A2(n608), .ZN(n610) );
  XOR2_X1 U689 ( .A(n610), .B(KEYINPUT31), .Z(n661) );
  NAND2_X1 U690 ( .A1(n643), .A2(G1996), .ZN(n611) );
  XNOR2_X1 U691 ( .A(n611), .B(KEYINPUT26), .ZN(n613) );
  NAND2_X1 U692 ( .A1(n642), .A2(G1341), .ZN(n612) );
  NAND2_X1 U693 ( .A1(n613), .A2(n612), .ZN(n626) );
  NAND2_X1 U694 ( .A1(G81), .A2(n800), .ZN(n616) );
  NAND2_X1 U695 ( .A1(G68), .A2(n801), .ZN(n617) );
  NAND2_X1 U696 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U697 ( .A(KEYINPUT13), .B(n619), .ZN(n625) );
  NAND2_X1 U698 ( .A1(G56), .A2(n804), .ZN(n620) );
  XOR2_X1 U699 ( .A(KEYINPUT14), .B(n620), .Z(n623) );
  NAND2_X1 U700 ( .A1(n805), .A2(G43), .ZN(n621) );
  XOR2_X1 U701 ( .A(KEYINPUT74), .B(n621), .Z(n622) );
  NOR2_X1 U702 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X1 U703 ( .A1(n625), .A2(n624), .ZN(n946) );
  NOR2_X1 U704 ( .A1(n626), .A2(n946), .ZN(n639) );
  NAND2_X1 U705 ( .A1(G92), .A2(n800), .ZN(n628) );
  NAND2_X1 U706 ( .A1(G79), .A2(n801), .ZN(n627) );
  NAND2_X1 U707 ( .A1(n628), .A2(n627), .ZN(n632) );
  NAND2_X1 U708 ( .A1(G66), .A2(n804), .ZN(n630) );
  NAND2_X1 U709 ( .A1(G54), .A2(n805), .ZN(n629) );
  NAND2_X1 U710 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U711 ( .A1(n632), .A2(n631), .ZN(n633) );
  XOR2_X1 U712 ( .A(KEYINPUT15), .B(n633), .Z(n945) );
  NAND2_X1 U713 ( .A1(n639), .A2(n945), .ZN(n638) );
  NAND2_X1 U714 ( .A1(n665), .A2(G1348), .ZN(n634) );
  XNOR2_X1 U715 ( .A(n634), .B(KEYINPUT90), .ZN(n636) );
  NAND2_X1 U716 ( .A1(n605), .A2(G2067), .ZN(n635) );
  NAND2_X1 U717 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U718 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U719 ( .A1(n641), .A2(n640), .ZN(n650) );
  NAND2_X1 U720 ( .A1(G1956), .A2(n642), .ZN(n647) );
  NAND2_X1 U721 ( .A1(n643), .A2(G2072), .ZN(n645) );
  NAND2_X1 U722 ( .A1(n647), .A2(n646), .ZN(n651) );
  XNOR2_X1 U723 ( .A(n648), .B(KEYINPUT91), .ZN(n649) );
  NAND2_X1 U724 ( .A1(n650), .A2(n649), .ZN(n654) );
  NAND2_X1 U725 ( .A1(G299), .A2(n651), .ZN(n652) );
  XNOR2_X1 U726 ( .A(n652), .B(KEYINPUT28), .ZN(n653) );
  NAND2_X1 U727 ( .A1(n654), .A2(n653), .ZN(n656) );
  XOR2_X1 U728 ( .A(KEYINPUT92), .B(KEYINPUT29), .Z(n655) );
  XNOR2_X1 U729 ( .A(n656), .B(n655), .ZN(n659) );
  NAND2_X1 U730 ( .A1(n657), .A2(G171), .ZN(n658) );
  NAND2_X1 U731 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U732 ( .A1(n661), .A2(n660), .ZN(n663) );
  XNOR2_X1 U733 ( .A(n663), .B(n662), .ZN(n676) );
  NAND2_X1 U734 ( .A1(n676), .A2(G286), .ZN(n673) );
  NAND2_X1 U735 ( .A1(G8), .A2(n665), .ZN(n708) );
  NOR2_X1 U736 ( .A1(G1971), .A2(n708), .ZN(n664) );
  XNOR2_X1 U737 ( .A(n664), .B(KEYINPUT94), .ZN(n667) );
  NOR2_X1 U738 ( .A1(n665), .A2(G2090), .ZN(n666) );
  NOR2_X1 U739 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U740 ( .A1(n668), .A2(G303), .ZN(n669) );
  XOR2_X1 U741 ( .A(KEYINPUT95), .B(n669), .Z(n670) );
  OR2_X1 U742 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U743 ( .A(n675), .B(n674), .ZN(n682) );
  NAND2_X1 U744 ( .A1(G8), .A2(n677), .ZN(n678) );
  NAND2_X1 U745 ( .A1(n676), .A2(n678), .ZN(n680) );
  NOR2_X1 U746 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X2 U747 ( .A1(n682), .A2(n681), .ZN(n698) );
  NOR2_X1 U748 ( .A1(G1971), .A2(G303), .ZN(n683) );
  XNOR2_X1 U749 ( .A(KEYINPUT96), .B(n683), .ZN(n684) );
  NOR2_X2 U750 ( .A1(n698), .A2(n684), .ZN(n686) );
  XNOR2_X1 U751 ( .A(n686), .B(n685), .ZN(n687) );
  NAND2_X1 U752 ( .A1(n688), .A2(n687), .ZN(n696) );
  XNOR2_X1 U753 ( .A(G1981), .B(G305), .ZN(n965) );
  NAND2_X1 U754 ( .A1(G1976), .A2(G288), .ZN(n953) );
  INV_X1 U755 ( .A(n953), .ZN(n689) );
  NOR2_X1 U756 ( .A1(KEYINPUT33), .A2(n513), .ZN(n690) );
  NOR2_X1 U757 ( .A1(n965), .A2(n690), .ZN(n694) );
  NOR2_X1 U758 ( .A1(KEYINPUT33), .A2(KEYINPUT97), .ZN(n691) );
  NOR2_X1 U759 ( .A1(n708), .A2(n691), .ZN(n692) );
  NAND2_X1 U760 ( .A1(n955), .A2(n692), .ZN(n693) );
  AND2_X1 U761 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U762 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U763 ( .A(n697), .B(KEYINPUT98), .ZN(n704) );
  INV_X1 U764 ( .A(n698), .ZN(n701) );
  NOR2_X1 U765 ( .A1(G2090), .A2(G303), .ZN(n699) );
  NAND2_X1 U766 ( .A1(G8), .A2(n699), .ZN(n700) );
  NAND2_X1 U767 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U768 ( .A1(n702), .A2(n708), .ZN(n703) );
  NAND2_X1 U769 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U770 ( .A(n705), .B(KEYINPUT99), .ZN(n710) );
  NOR2_X1 U771 ( .A1(G1981), .A2(G305), .ZN(n706) );
  XOR2_X1 U772 ( .A(n706), .B(KEYINPUT24), .Z(n707) );
  OR2_X1 U773 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U774 ( .A1(n710), .A2(n709), .ZN(n741) );
  NAND2_X1 U775 ( .A1(G131), .A2(n894), .ZN(n712) );
  NAND2_X1 U776 ( .A1(G119), .A2(n590), .ZN(n711) );
  NAND2_X1 U777 ( .A1(n712), .A2(n711), .ZN(n716) );
  NAND2_X1 U778 ( .A1(G95), .A2(n891), .ZN(n714) );
  NAND2_X1 U779 ( .A1(G107), .A2(n887), .ZN(n713) );
  NAND2_X1 U780 ( .A1(n714), .A2(n713), .ZN(n715) );
  OR2_X1 U781 ( .A1(n716), .A2(n715), .ZN(n884) );
  AND2_X1 U782 ( .A1(n884), .A2(G1991), .ZN(n725) );
  NAND2_X1 U783 ( .A1(G141), .A2(n894), .ZN(n718) );
  NAND2_X1 U784 ( .A1(G129), .A2(n590), .ZN(n717) );
  NAND2_X1 U785 ( .A1(n718), .A2(n717), .ZN(n721) );
  NAND2_X1 U786 ( .A1(n891), .A2(G105), .ZN(n719) );
  XOR2_X1 U787 ( .A(KEYINPUT38), .B(n719), .Z(n720) );
  NOR2_X1 U788 ( .A1(n721), .A2(n720), .ZN(n723) );
  NAND2_X1 U789 ( .A1(n887), .A2(G117), .ZN(n722) );
  NAND2_X1 U790 ( .A1(n723), .A2(n722), .ZN(n874) );
  AND2_X1 U791 ( .A1(G1996), .A2(n874), .ZN(n724) );
  NOR2_X1 U792 ( .A1(n725), .A2(n724), .ZN(n927) );
  NOR2_X1 U793 ( .A1(n727), .A2(n726), .ZN(n757) );
  INV_X1 U794 ( .A(n757), .ZN(n728) );
  NOR2_X1 U795 ( .A1(n927), .A2(n728), .ZN(n751) );
  XNOR2_X1 U796 ( .A(KEYINPUT89), .B(n751), .ZN(n739) );
  XNOR2_X1 U797 ( .A(G2067), .B(KEYINPUT37), .ZN(n746) );
  XNOR2_X1 U798 ( .A(KEYINPUT88), .B(KEYINPUT34), .ZN(n732) );
  NAND2_X1 U799 ( .A1(G140), .A2(n894), .ZN(n730) );
  NAND2_X1 U800 ( .A1(G104), .A2(n891), .ZN(n729) );
  NAND2_X1 U801 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U802 ( .A(n732), .B(n731), .ZN(n737) );
  NAND2_X1 U803 ( .A1(G128), .A2(n590), .ZN(n734) );
  NAND2_X1 U804 ( .A1(G116), .A2(n887), .ZN(n733) );
  NAND2_X1 U805 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U806 ( .A(KEYINPUT35), .B(n735), .Z(n736) );
  NOR2_X1 U807 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U808 ( .A(KEYINPUT36), .B(n738), .ZN(n903) );
  NOR2_X1 U809 ( .A1(n746), .A2(n903), .ZN(n930) );
  NAND2_X1 U810 ( .A1(n757), .A2(n930), .ZN(n754) );
  AND2_X1 U811 ( .A1(n739), .A2(n754), .ZN(n740) );
  NAND2_X1 U812 ( .A1(n741), .A2(n740), .ZN(n743) );
  XNOR2_X1 U813 ( .A(n743), .B(n742), .ZN(n745) );
  XNOR2_X1 U814 ( .A(G1986), .B(G290), .ZN(n951) );
  NAND2_X1 U815 ( .A1(n951), .A2(n757), .ZN(n744) );
  NAND2_X1 U816 ( .A1(n745), .A2(n744), .ZN(n760) );
  NAND2_X1 U817 ( .A1(n903), .A2(n746), .ZN(n747) );
  XNOR2_X1 U818 ( .A(n747), .B(KEYINPUT102), .ZN(n936) );
  NOR2_X1 U819 ( .A1(G1996), .A2(n874), .ZN(n923) );
  NOR2_X1 U820 ( .A1(G1986), .A2(G290), .ZN(n748) );
  NOR2_X1 U821 ( .A1(G1991), .A2(n884), .ZN(n932) );
  NOR2_X1 U822 ( .A1(n748), .A2(n932), .ZN(n749) );
  XOR2_X1 U823 ( .A(KEYINPUT101), .B(n749), .Z(n750) );
  NOR2_X1 U824 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U825 ( .A1(n923), .A2(n752), .ZN(n753) );
  XNOR2_X1 U826 ( .A(KEYINPUT39), .B(n753), .ZN(n755) );
  NAND2_X1 U827 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U828 ( .A1(n936), .A2(n756), .ZN(n758) );
  NAND2_X1 U829 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U830 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U831 ( .A(n761), .B(KEYINPUT40), .ZN(G329) );
  BUF_X1 U832 ( .A(n762), .Z(G160) );
  XOR2_X1 U833 ( .A(G2443), .B(KEYINPUT106), .Z(n764) );
  XNOR2_X1 U834 ( .A(G1348), .B(G1341), .ZN(n763) );
  XNOR2_X1 U835 ( .A(n764), .B(n763), .ZN(n774) );
  XOR2_X1 U836 ( .A(G2446), .B(KEYINPUT105), .Z(n766) );
  XNOR2_X1 U837 ( .A(G2430), .B(G2438), .ZN(n765) );
  XNOR2_X1 U838 ( .A(n766), .B(n765), .ZN(n770) );
  XOR2_X1 U839 ( .A(KEYINPUT104), .B(KEYINPUT103), .Z(n768) );
  XNOR2_X1 U840 ( .A(G2435), .B(G2454), .ZN(n767) );
  XNOR2_X1 U841 ( .A(n768), .B(n767), .ZN(n769) );
  XOR2_X1 U842 ( .A(n770), .B(n769), .Z(n772) );
  XNOR2_X1 U843 ( .A(G2427), .B(G2451), .ZN(n771) );
  XNOR2_X1 U844 ( .A(n772), .B(n771), .ZN(n773) );
  XNOR2_X1 U845 ( .A(n774), .B(n773), .ZN(n775) );
  AND2_X1 U846 ( .A1(n775), .A2(G14), .ZN(G401) );
  AND2_X1 U847 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U848 ( .A(G132), .ZN(G219) );
  INV_X1 U849 ( .A(G57), .ZN(G237) );
  XOR2_X1 U850 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n778) );
  NAND2_X1 U851 ( .A1(G7), .A2(G661), .ZN(n776) );
  XOR2_X1 U852 ( .A(n776), .B(KEYINPUT10), .Z(n917) );
  NAND2_X1 U853 ( .A1(G567), .A2(n917), .ZN(n777) );
  XNOR2_X1 U854 ( .A(n778), .B(n777), .ZN(G234) );
  INV_X1 U855 ( .A(G860), .ZN(n783) );
  OR2_X1 U856 ( .A1(n946), .A2(n783), .ZN(G153) );
  XNOR2_X1 U857 ( .A(G171), .B(KEYINPUT75), .ZN(G301) );
  NAND2_X1 U858 ( .A1(G868), .A2(G301), .ZN(n780) );
  OR2_X1 U859 ( .A1(n945), .A2(G868), .ZN(n779) );
  NAND2_X1 U860 ( .A1(n780), .A2(n779), .ZN(G284) );
  INV_X1 U861 ( .A(G868), .ZN(n819) );
  NOR2_X1 U862 ( .A1(G286), .A2(n819), .ZN(n782) );
  NOR2_X1 U863 ( .A1(G868), .A2(G299), .ZN(n781) );
  NOR2_X1 U864 ( .A1(n782), .A2(n781), .ZN(G297) );
  NAND2_X1 U865 ( .A1(n783), .A2(G559), .ZN(n784) );
  NAND2_X1 U866 ( .A1(n784), .A2(n945), .ZN(n785) );
  XNOR2_X1 U867 ( .A(n785), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U868 ( .A1(G868), .A2(n946), .ZN(n786) );
  XNOR2_X1 U869 ( .A(KEYINPUT78), .B(n786), .ZN(n789) );
  NAND2_X1 U870 ( .A1(G868), .A2(n945), .ZN(n787) );
  NOR2_X1 U871 ( .A1(G559), .A2(n787), .ZN(n788) );
  NOR2_X1 U872 ( .A1(n789), .A2(n788), .ZN(G282) );
  NAND2_X1 U873 ( .A1(G123), .A2(n590), .ZN(n790) );
  XNOR2_X1 U874 ( .A(n790), .B(KEYINPUT18), .ZN(n792) );
  NAND2_X1 U875 ( .A1(n891), .A2(G99), .ZN(n791) );
  NAND2_X1 U876 ( .A1(n792), .A2(n791), .ZN(n796) );
  NAND2_X1 U877 ( .A1(G135), .A2(n894), .ZN(n794) );
  NAND2_X1 U878 ( .A1(G111), .A2(n887), .ZN(n793) );
  NAND2_X1 U879 ( .A1(n794), .A2(n793), .ZN(n795) );
  NOR2_X1 U880 ( .A1(n796), .A2(n795), .ZN(n931) );
  XOR2_X1 U881 ( .A(n931), .B(G2096), .Z(n797) );
  NOR2_X1 U882 ( .A1(G2100), .A2(n797), .ZN(n798) );
  XNOR2_X1 U883 ( .A(KEYINPUT79), .B(n798), .ZN(G156) );
  NAND2_X1 U884 ( .A1(n945), .A2(G559), .ZN(n817) );
  XNOR2_X1 U885 ( .A(n946), .B(n817), .ZN(n799) );
  NOR2_X1 U886 ( .A1(n799), .A2(G860), .ZN(n810) );
  NAND2_X1 U887 ( .A1(G93), .A2(n800), .ZN(n803) );
  NAND2_X1 U888 ( .A1(G80), .A2(n801), .ZN(n802) );
  NAND2_X1 U889 ( .A1(n803), .A2(n802), .ZN(n809) );
  NAND2_X1 U890 ( .A1(G67), .A2(n804), .ZN(n807) );
  NAND2_X1 U891 ( .A1(G55), .A2(n805), .ZN(n806) );
  NAND2_X1 U892 ( .A1(n807), .A2(n806), .ZN(n808) );
  OR2_X1 U893 ( .A1(n809), .A2(n808), .ZN(n820) );
  XOR2_X1 U894 ( .A(n810), .B(n820), .Z(G145) );
  XOR2_X1 U895 ( .A(G166), .B(KEYINPUT19), .Z(n811) );
  XNOR2_X1 U896 ( .A(G288), .B(n811), .ZN(n814) );
  XOR2_X1 U897 ( .A(G290), .B(G305), .Z(n812) );
  XNOR2_X1 U898 ( .A(n946), .B(n812), .ZN(n813) );
  XNOR2_X1 U899 ( .A(n814), .B(n813), .ZN(n816) );
  XOR2_X1 U900 ( .A(G299), .B(n820), .Z(n815) );
  XNOR2_X1 U901 ( .A(n816), .B(n815), .ZN(n906) );
  XOR2_X1 U902 ( .A(n906), .B(n817), .Z(n818) );
  NAND2_X1 U903 ( .A1(G868), .A2(n818), .ZN(n822) );
  NAND2_X1 U904 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U905 ( .A1(n822), .A2(n821), .ZN(G295) );
  NAND2_X1 U906 ( .A1(G2078), .A2(G2084), .ZN(n823) );
  XOR2_X1 U907 ( .A(KEYINPUT20), .B(n823), .Z(n824) );
  NAND2_X1 U908 ( .A1(G2090), .A2(n824), .ZN(n825) );
  XNOR2_X1 U909 ( .A(KEYINPUT21), .B(n825), .ZN(n826) );
  NAND2_X1 U910 ( .A1(n826), .A2(G2072), .ZN(G158) );
  XOR2_X1 U911 ( .A(KEYINPUT83), .B(G44), .Z(n827) );
  XNOR2_X1 U912 ( .A(KEYINPUT3), .B(n827), .ZN(G218) );
  XNOR2_X1 U913 ( .A(KEYINPUT71), .B(G82), .ZN(G220) );
  NAND2_X1 U914 ( .A1(G69), .A2(G120), .ZN(n828) );
  NOR2_X1 U915 ( .A1(G237), .A2(n828), .ZN(n829) );
  NAND2_X1 U916 ( .A1(G108), .A2(n829), .ZN(n844) );
  NAND2_X1 U917 ( .A1(G567), .A2(n844), .ZN(n836) );
  NOR2_X1 U918 ( .A1(G219), .A2(G220), .ZN(n830) );
  XOR2_X1 U919 ( .A(KEYINPUT84), .B(n830), .Z(n831) );
  XNOR2_X1 U920 ( .A(n831), .B(KEYINPUT22), .ZN(n832) );
  NOR2_X1 U921 ( .A1(G218), .A2(n832), .ZN(n833) );
  XOR2_X1 U922 ( .A(KEYINPUT85), .B(n833), .Z(n834) );
  NAND2_X1 U923 ( .A1(G96), .A2(n834), .ZN(n843) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n843), .ZN(n835) );
  NAND2_X1 U925 ( .A1(n836), .A2(n835), .ZN(n845) );
  NAND2_X1 U926 ( .A1(G661), .A2(G483), .ZN(n837) );
  XNOR2_X1 U927 ( .A(KEYINPUT86), .B(n837), .ZN(n838) );
  NOR2_X1 U928 ( .A1(n845), .A2(n838), .ZN(n842) );
  NAND2_X1 U929 ( .A1(n842), .A2(G36), .ZN(G176) );
  NAND2_X1 U930 ( .A1(G2106), .A2(n917), .ZN(G217) );
  NAND2_X1 U931 ( .A1(G15), .A2(G2), .ZN(n839) );
  XNOR2_X1 U932 ( .A(KEYINPUT107), .B(n839), .ZN(n840) );
  NAND2_X1 U933 ( .A1(n840), .A2(G661), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n841) );
  NAND2_X1 U935 ( .A1(n842), .A2(n841), .ZN(G188) );
  INV_X1 U937 ( .A(G120), .ZN(G236) );
  INV_X1 U938 ( .A(G96), .ZN(G221) );
  INV_X1 U939 ( .A(G69), .ZN(G235) );
  NOR2_X1 U940 ( .A1(n844), .A2(n843), .ZN(G325) );
  INV_X1 U941 ( .A(G325), .ZN(G261) );
  INV_X1 U942 ( .A(n845), .ZN(G319) );
  XOR2_X1 U943 ( .A(G1976), .B(G1971), .Z(n847) );
  XNOR2_X1 U944 ( .A(G1981), .B(G1966), .ZN(n846) );
  XNOR2_X1 U945 ( .A(n847), .B(n846), .ZN(n857) );
  XOR2_X1 U946 ( .A(KEYINPUT110), .B(KEYINPUT109), .Z(n849) );
  XNOR2_X1 U947 ( .A(G1991), .B(G2474), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(n853) );
  XNOR2_X1 U949 ( .A(G1956), .B(n949), .ZN(n851) );
  XNOR2_X1 U950 ( .A(G1996), .B(G1986), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U952 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U953 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U955 ( .A(n857), .B(n856), .Z(G229) );
  XOR2_X1 U956 ( .A(G2096), .B(KEYINPUT43), .Z(n859) );
  XNOR2_X1 U957 ( .A(G2090), .B(KEYINPUT42), .ZN(n858) );
  XNOR2_X1 U958 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U959 ( .A(n860), .B(G2678), .Z(n862) );
  XNOR2_X1 U960 ( .A(G2067), .B(G2072), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U962 ( .A(KEYINPUT108), .B(G2100), .Z(n864) );
  XNOR2_X1 U963 ( .A(G2078), .B(G2084), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n864), .B(n863), .ZN(n865) );
  XNOR2_X1 U965 ( .A(n866), .B(n865), .ZN(G227) );
  NAND2_X1 U966 ( .A1(G124), .A2(n590), .ZN(n867) );
  XNOR2_X1 U967 ( .A(n867), .B(KEYINPUT44), .ZN(n869) );
  NAND2_X1 U968 ( .A1(n891), .A2(G100), .ZN(n868) );
  NAND2_X1 U969 ( .A1(n869), .A2(n868), .ZN(n873) );
  NAND2_X1 U970 ( .A1(G136), .A2(n894), .ZN(n871) );
  NAND2_X1 U971 ( .A1(G112), .A2(n887), .ZN(n870) );
  NAND2_X1 U972 ( .A1(n871), .A2(n870), .ZN(n872) );
  NOR2_X1 U973 ( .A1(n873), .A2(n872), .ZN(G162) );
  XOR2_X1 U974 ( .A(G162), .B(n931), .Z(n876) );
  XOR2_X1 U975 ( .A(G164), .B(n874), .Z(n875) );
  XNOR2_X1 U976 ( .A(n876), .B(n875), .ZN(n901) );
  NAND2_X1 U977 ( .A1(G130), .A2(n590), .ZN(n878) );
  NAND2_X1 U978 ( .A1(G118), .A2(n887), .ZN(n877) );
  NAND2_X1 U979 ( .A1(n878), .A2(n877), .ZN(n883) );
  NAND2_X1 U980 ( .A1(G142), .A2(n894), .ZN(n880) );
  NAND2_X1 U981 ( .A1(G106), .A2(n891), .ZN(n879) );
  NAND2_X1 U982 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U983 ( .A(n881), .B(KEYINPUT45), .Z(n882) );
  NOR2_X1 U984 ( .A1(n883), .A2(n882), .ZN(n885) );
  XNOR2_X1 U985 ( .A(n885), .B(n884), .ZN(n886) );
  XOR2_X1 U986 ( .A(n886), .B(KEYINPUT46), .Z(n899) );
  NAND2_X1 U987 ( .A1(G127), .A2(n590), .ZN(n889) );
  NAND2_X1 U988 ( .A1(G115), .A2(n887), .ZN(n888) );
  NAND2_X1 U989 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U990 ( .A(n890), .B(KEYINPUT47), .ZN(n893) );
  NAND2_X1 U991 ( .A1(G103), .A2(n891), .ZN(n892) );
  NAND2_X1 U992 ( .A1(n893), .A2(n892), .ZN(n897) );
  NAND2_X1 U993 ( .A1(n894), .A2(G139), .ZN(n895) );
  XOR2_X1 U994 ( .A(KEYINPUT112), .B(n895), .Z(n896) );
  NOR2_X1 U995 ( .A1(n897), .A2(n896), .ZN(n918) );
  XNOR2_X1 U996 ( .A(n918), .B(KEYINPUT48), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U998 ( .A(n901), .B(n900), .Z(n902) );
  XNOR2_X1 U999 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U1000 ( .A(n904), .B(G160), .ZN(n905) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n905), .ZN(G395) );
  XOR2_X1 U1002 ( .A(KEYINPUT113), .B(n906), .Z(n908) );
  XNOR2_X1 U1003 ( .A(G171), .B(G286), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(n908), .B(n907), .ZN(n909) );
  XNOR2_X1 U1005 ( .A(n909), .B(n945), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n910), .ZN(G397) );
  NOR2_X1 U1007 ( .A1(G229), .A2(G227), .ZN(n911) );
  XOR2_X1 U1008 ( .A(KEYINPUT49), .B(n911), .Z(n912) );
  NAND2_X1 U1009 ( .A1(G319), .A2(n912), .ZN(n913) );
  NOR2_X1 U1010 ( .A1(G401), .A2(n913), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(KEYINPUT114), .B(n914), .ZN(n916) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n915) );
  NAND2_X1 U1013 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(G108), .ZN(G238) );
  INV_X1 U1016 ( .A(n917), .ZN(G223) );
  XNOR2_X1 U1017 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n1027) );
  INV_X1 U1018 ( .A(KEYINPUT55), .ZN(n1018) );
  XNOR2_X1 U1019 ( .A(KEYINPUT52), .B(KEYINPUT116), .ZN(n941) );
  XOR2_X1 U1020 ( .A(G2072), .B(n918), .Z(n920) );
  XOR2_X1 U1021 ( .A(G164), .B(G2078), .Z(n919) );
  NOR2_X1 U1022 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1023 ( .A(KEYINPUT50), .B(n921), .ZN(n926) );
  XOR2_X1 U1024 ( .A(G2090), .B(G162), .Z(n922) );
  NOR2_X1 U1025 ( .A1(n923), .A2(n922), .ZN(n924) );
  XOR2_X1 U1026 ( .A(KEYINPUT51), .B(n924), .Z(n925) );
  NAND2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n939) );
  XNOR2_X1 U1028 ( .A(G2084), .B(G160), .ZN(n928) );
  NAND2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1030 ( .A1(n930), .A2(n929), .ZN(n934) );
  NOR2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1033 ( .A(KEYINPUT115), .B(n935), .ZN(n937) );
  NAND2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1036 ( .A(n941), .B(n940), .ZN(n942) );
  NAND2_X1 U1037 ( .A1(n1018), .A2(n942), .ZN(n943) );
  NAND2_X1 U1038 ( .A1(n943), .A2(G29), .ZN(n1025) );
  XNOR2_X1 U1039 ( .A(KEYINPUT56), .B(KEYINPUT121), .ZN(n944) );
  XOR2_X1 U1040 ( .A(G16), .B(n944), .Z(n970) );
  XOR2_X1 U1041 ( .A(G1348), .B(n945), .Z(n948) );
  XNOR2_X1 U1042 ( .A(n946), .B(G1341), .ZN(n947) );
  NOR2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n962) );
  XNOR2_X1 U1044 ( .A(G171), .B(n949), .ZN(n950) );
  NOR2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n957) );
  XOR2_X1 U1046 ( .A(G1956), .B(G299), .Z(n952) );
  NAND2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1049 ( .A1(n957), .A2(n956), .ZN(n960) );
  XNOR2_X1 U1050 ( .A(G1971), .B(G303), .ZN(n958) );
  XNOR2_X1 U1051 ( .A(KEYINPUT122), .B(n958), .ZN(n959) );
  NOR2_X1 U1052 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1053 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1054 ( .A(KEYINPUT123), .B(n963), .ZN(n968) );
  XOR2_X1 U1055 ( .A(G1966), .B(G168), .Z(n964) );
  NOR2_X1 U1056 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1057 ( .A(KEYINPUT57), .B(n966), .Z(n967) );
  NAND2_X1 U1058 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1059 ( .A1(n970), .A2(n969), .ZN(n996) );
  INV_X1 U1060 ( .A(G16), .ZN(n994) );
  XOR2_X1 U1061 ( .A(G1986), .B(KEYINPUT124), .Z(n971) );
  XNOR2_X1 U1062 ( .A(G24), .B(n971), .ZN(n975) );
  XNOR2_X1 U1063 ( .A(G1971), .B(G22), .ZN(n973) );
  XNOR2_X1 U1064 ( .A(G23), .B(G1976), .ZN(n972) );
  NOR2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1067 ( .A(KEYINPUT58), .B(n976), .Z(n990) );
  XOR2_X1 U1068 ( .A(G1966), .B(G21), .Z(n978) );
  XOR2_X1 U1069 ( .A(G1961), .B(G5), .Z(n977) );
  NAND2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n988) );
  XOR2_X1 U1071 ( .A(G1348), .B(KEYINPUT59), .Z(n979) );
  XNOR2_X1 U1072 ( .A(G4), .B(n979), .ZN(n981) );
  XNOR2_X1 U1073 ( .A(G20), .B(G1956), .ZN(n980) );
  NOR2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n985) );
  XNOR2_X1 U1075 ( .A(G1981), .B(G6), .ZN(n983) );
  XNOR2_X1 U1076 ( .A(G19), .B(G1341), .ZN(n982) );
  NOR2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(KEYINPUT60), .B(n986), .ZN(n987) );
  NOR2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1082 ( .A(n991), .B(KEYINPUT125), .ZN(n992) );
  XNOR2_X1 U1083 ( .A(KEYINPUT61), .B(n992), .ZN(n993) );
  NAND2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n1021) );
  XNOR2_X1 U1086 ( .A(G2084), .B(G34), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(n997), .B(KEYINPUT54), .ZN(n999) );
  XNOR2_X1 U1088 ( .A(G35), .B(G2090), .ZN(n998) );
  NOR2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1016) );
  XNOR2_X1 U1090 ( .A(G27), .B(n1000), .ZN(n1007) );
  XNOR2_X1 U1091 ( .A(G2067), .B(G26), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(G2072), .B(G33), .ZN(n1001) );
  NOR2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1094 ( .A(KEYINPUT118), .B(n1003), .Z(n1005) );
  XNOR2_X1 U1095 ( .A(G1996), .B(G32), .ZN(n1004) );
  NOR2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1098 ( .A(KEYINPUT119), .B(n1008), .ZN(n1009) );
  NAND2_X1 U1099 ( .A1(n1009), .A2(G28), .ZN(n1012) );
  XOR2_X1 U1100 ( .A(G25), .B(G1991), .Z(n1010) );
  XNOR2_X1 U1101 ( .A(KEYINPUT117), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1103 ( .A(n1013), .B(KEYINPUT53), .Z(n1014) );
  XNOR2_X1 U1104 ( .A(KEYINPUT120), .B(n1014), .ZN(n1015) );
  NAND2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1106 ( .A(n1018), .B(n1017), .Z(n1019) );
  NOR2_X1 U1107 ( .A1(G29), .A2(n1019), .ZN(n1020) );
  NOR2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1109 ( .A1(G11), .A2(n1022), .ZN(n1023) );
  XOR2_X1 U1110 ( .A(KEYINPUT126), .B(n1023), .Z(n1024) );
  NAND2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1112 ( .A(n1027), .B(n1026), .Z(G150) );
  INV_X1 U1113 ( .A(G150), .ZN(G311) );
endmodule

