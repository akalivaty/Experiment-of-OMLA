

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n638, n639, n640, n641, n642,
         n643, n644, n646, n647, n648, n649, n650, n651, n652, n653, n655,
         n656, n657, n658, n659, n660, n661, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755;

  AND2_X1 U366 ( .A1(n348), .A2(n347), .ZN(n646) );
  INV_X1 U367 ( .A(n737), .ZN(n344) );
  INV_X1 U368 ( .A(n737), .ZN(n347) );
  INV_X1 U369 ( .A(n737), .ZN(n350) );
  INV_X1 U370 ( .A(n737), .ZN(n353) );
  INV_X1 U371 ( .A(n635), .ZN(n346) );
  INV_X1 U372 ( .A(n643), .ZN(n349) );
  INV_X1 U373 ( .A(n660), .ZN(n352) );
  INV_X1 U374 ( .A(n652), .ZN(n355) );
  INV_X1 U375 ( .A(n693), .ZN(n576) );
  XNOR2_X1 U376 ( .A(n458), .B(n457), .ZN(n617) );
  XNOR2_X1 U377 ( .A(G122), .B(G104), .ZN(n498) );
  INV_X1 U378 ( .A(KEYINPUT87), .ZN(n429) );
  XNOR2_X2 U379 ( .A(n616), .B(n615), .ZN(n368) );
  AND2_X2 U380 ( .A1(n345), .A2(n344), .ZN(n640) );
  XNOR2_X1 U381 ( .A(n636), .B(n346), .ZN(n345) );
  XNOR2_X1 U382 ( .A(n644), .B(n349), .ZN(n348) );
  AND2_X2 U383 ( .A1(n351), .A2(n350), .ZN(n664) );
  XNOR2_X1 U384 ( .A(n661), .B(n352), .ZN(n351) );
  AND2_X2 U385 ( .A1(n354), .A2(n353), .ZN(n655) );
  XNOR2_X1 U386 ( .A(n653), .B(n355), .ZN(n354) );
  XNOR2_X2 U387 ( .A(n699), .B(KEYINPUT6), .ZN(n553) );
  XNOR2_X2 U388 ( .A(n356), .B(KEYINPUT45), .ZN(n611) );
  NAND2_X2 U389 ( .A1(n371), .A2(n362), .ZN(n356) );
  INV_X1 U390 ( .A(G104), .ZN(n441) );
  INV_X1 U391 ( .A(G110), .ZN(n438) );
  INV_X1 U392 ( .A(G953), .ZN(n448) );
  AND2_X2 U393 ( .A1(n375), .A2(n547), .ZN(n371) );
  AND2_X1 U394 ( .A1(n604), .A2(n603), .ZN(n741) );
  NOR2_X1 U395 ( .A1(n406), .A2(KEYINPUT44), .ZN(n405) );
  NAND2_X1 U396 ( .A1(n625), .A2(n623), .ZN(n406) );
  NOR2_X1 U397 ( .A1(n527), .A2(n369), .ZN(n543) );
  NOR2_X1 U398 ( .A1(n555), .A2(n373), .ZN(n593) );
  XNOR2_X1 U399 ( .A(n592), .B(n370), .ZN(n676) );
  XNOR2_X1 U400 ( .A(n382), .B(KEYINPUT19), .ZN(n578) );
  NOR2_X1 U401 ( .A1(n540), .A2(n539), .ZN(n592) );
  NAND2_X1 U402 ( .A1(n376), .A2(n381), .ZN(n382) );
  XNOR2_X1 U403 ( .A(n656), .B(n659), .ZN(n660) );
  XNOR2_X1 U404 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U405 ( .A(n634), .B(KEYINPUT62), .ZN(n635) );
  OR2_X1 U406 ( .A1(n656), .A2(n378), .ZN(n377) );
  XNOR2_X1 U407 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U408 ( .A(n433), .B(n432), .ZN(n471) );
  NOR2_X1 U409 ( .A1(n753), .A2(n755), .ZN(n416) );
  AND2_X1 U410 ( .A1(n372), .A2(n583), .ZN(n385) );
  NOR2_X1 U411 ( .A1(n361), .A2(n682), .ZN(n372) );
  NAND2_X1 U412 ( .A1(n379), .A2(n606), .ZN(n378) );
  XNOR2_X1 U413 ( .A(n465), .B(n464), .ZN(n693) );
  XNOR2_X1 U414 ( .A(n463), .B(n462), .ZN(n464) );
  OR2_X1 U415 ( .A1(n634), .A2(G902), .ZN(n413) );
  XNOR2_X1 U416 ( .A(n401), .B(n591), .ZN(n599) );
  NAND2_X1 U417 ( .A1(n409), .A2(n459), .ZN(n408) );
  INV_X1 U418 ( .A(G469), .ZN(n409) );
  NAND2_X1 U419 ( .A1(G902), .A2(G469), .ZN(n411) );
  XNOR2_X1 U420 ( .A(n455), .B(G140), .ZN(n492) );
  XNOR2_X1 U421 ( .A(G125), .B(KEYINPUT10), .ZN(n455) );
  XNOR2_X1 U422 ( .A(n383), .B(n414), .ZN(n604) );
  XNOR2_X1 U423 ( .A(n416), .B(KEYINPUT46), .ZN(n415) );
  NOR2_X1 U424 ( .A1(n576), .A2(n357), .ZN(n392) );
  NAND2_X1 U425 ( .A1(n482), .A2(n549), .ZN(n380) );
  XOR2_X1 U426 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n451) );
  XNOR2_X1 U427 ( .A(G128), .B(G146), .ZN(n450) );
  XNOR2_X1 U428 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U429 ( .A(n475), .B(n476), .ZN(n477) );
  NAND2_X1 U430 ( .A1(n561), .A2(n363), .ZN(n373) );
  NAND2_X1 U431 ( .A1(n554), .A2(n676), .ZN(n555) );
  XNOR2_X1 U432 ( .A(n567), .B(KEYINPUT30), .ZN(n388) );
  NOR2_X1 U433 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U434 ( .A1(n406), .A2(KEYINPUT44), .ZN(n402) );
  XNOR2_X1 U435 ( .A(G146), .B(KEYINPUT4), .ZN(n421) );
  XNOR2_X1 U436 ( .A(KEYINPUT18), .B(G125), .ZN(n473) );
  NAND2_X1 U437 ( .A1(G237), .A2(G234), .ZN(n484) );
  AND2_X1 U438 ( .A1(n377), .A2(n365), .ZN(n376) );
  XNOR2_X1 U439 ( .A(n438), .B(G107), .ZN(n468) );
  XNOR2_X1 U440 ( .A(KEYINPUT3), .B(G119), .ZN(n432) );
  XNOR2_X1 U441 ( .A(G116), .B(G113), .ZN(n430) );
  INV_X1 U442 ( .A(G134), .ZN(n420) );
  XNOR2_X1 U443 ( .A(G116), .B(G107), .ZN(n507) );
  XOR2_X1 U444 ( .A(KEYINPUT100), .B(G122), .Z(n508) );
  XNOR2_X1 U445 ( .A(G146), .B(G113), .ZN(n495) );
  XNOR2_X1 U446 ( .A(KEYINPUT97), .B(KEYINPUT11), .ZN(n490) );
  NOR2_X1 U447 ( .A1(n741), .A2(n684), .ZN(n685) );
  XNOR2_X1 U448 ( .A(n391), .B(n390), .ZN(n389) );
  INV_X1 U449 ( .A(KEYINPUT28), .ZN(n390) );
  INV_X1 U450 ( .A(n740), .ZN(n457) );
  XNOR2_X1 U451 ( .A(n400), .B(n399), .ZN(n753) );
  INV_X1 U452 ( .A(KEYINPUT40), .ZN(n399) );
  XNOR2_X1 U453 ( .A(n387), .B(n386), .ZN(n750) );
  INV_X1 U454 ( .A(KEYINPUT107), .ZN(n386) );
  INV_X1 U455 ( .A(KEYINPUT103), .ZN(n523) );
  NOR2_X1 U456 ( .A1(n538), .A2(n537), .ZN(n679) );
  INV_X1 U457 ( .A(KEYINPUT105), .ZN(n370) );
  NOR2_X1 U458 ( .A1(n731), .A2(G953), .ZN(n732) );
  OR2_X1 U459 ( .A1(n692), .A2(n575), .ZN(n357) );
  OR2_X1 U460 ( .A1(G902), .A2(n734), .ZN(n358) );
  XOR2_X1 U461 ( .A(n492), .B(n491), .Z(n359) );
  XOR2_X1 U462 ( .A(KEYINPUT96), .B(KEYINPUT12), .Z(n360) );
  AND2_X1 U463 ( .A1(n582), .A2(n581), .ZN(n361) );
  AND2_X1 U464 ( .A1(n403), .A2(n402), .ZN(n362) );
  AND2_X1 U465 ( .A1(n552), .A2(n707), .ZN(n363) );
  INV_X1 U466 ( .A(n606), .ZN(n549) );
  XNOR2_X1 U467 ( .A(KEYINPUT15), .B(G902), .ZN(n606) );
  INV_X1 U468 ( .A(G902), .ZN(n459) );
  AND2_X1 U469 ( .A1(n603), .A2(KEYINPUT2), .ZN(n364) );
  AND2_X1 U470 ( .A1(n380), .A2(n707), .ZN(n365) );
  AND2_X1 U471 ( .A1(n377), .A2(n380), .ZN(n366) );
  INV_X1 U472 ( .A(KEYINPUT1), .ZN(n397) );
  XNOR2_X1 U473 ( .A(n616), .B(n615), .ZN(n367) );
  XNOR2_X1 U474 ( .A(n616), .B(n615), .ZN(n733) );
  NAND2_X2 U475 ( .A1(n614), .A2(n688), .ZN(n616) );
  NOR2_X1 U476 ( .A1(n570), .A2(n388), .ZN(n590) );
  AND2_X2 U477 ( .A1(n412), .A2(n411), .ZN(n410) );
  OR2_X2 U478 ( .A1(n647), .A2(n408), .ZN(n407) );
  NAND2_X1 U479 ( .A1(n395), .A2(n410), .ZN(n394) );
  BUF_X1 U480 ( .A(n522), .Z(n369) );
  NAND2_X1 U481 ( .A1(n396), .A2(n394), .ZN(n522) );
  NAND2_X1 U482 ( .A1(n410), .A2(n407), .ZN(n393) );
  AND2_X2 U483 ( .A1(n407), .A2(n397), .ZN(n395) );
  XNOR2_X1 U484 ( .A(n531), .B(n466), .ZN(n374) );
  NOR2_X2 U485 ( .A1(n717), .A2(n535), .ZN(n417) );
  NAND2_X1 U486 ( .A1(n393), .A2(KEYINPUT1), .ZN(n396) );
  NOR2_X1 U487 ( .A1(n374), .A2(n553), .ZN(n467) );
  NAND2_X1 U488 ( .A1(n404), .A2(n405), .ZN(n375) );
  NAND2_X1 U489 ( .A1(n366), .A2(n381), .ZN(n562) );
  INV_X1 U490 ( .A(n482), .ZN(n379) );
  NAND2_X1 U491 ( .A1(n656), .A2(n482), .ZN(n381) );
  NAND2_X1 U492 ( .A1(n384), .A2(n415), .ZN(n383) );
  XNOR2_X1 U493 ( .A(n385), .B(KEYINPUT70), .ZN(n384) );
  NAND2_X1 U494 ( .A1(n590), .A2(n572), .ZN(n387) );
  NAND2_X1 U495 ( .A1(n389), .A2(n398), .ZN(n577) );
  NAND2_X1 U496 ( .A1(n699), .A2(n392), .ZN(n391) );
  NAND2_X1 U497 ( .A1(n407), .A2(n410), .ZN(n398) );
  NAND2_X1 U498 ( .A1(n696), .A2(n398), .ZN(n568) );
  NOR2_X1 U499 ( .A1(n535), .A2(n519), .ZN(n521) );
  NAND2_X1 U500 ( .A1(n604), .A2(n364), .ZN(n610) );
  NAND2_X1 U501 ( .A1(n599), .A2(n592), .ZN(n400) );
  NAND2_X1 U502 ( .A1(n590), .A2(n708), .ZN(n401) );
  NAND2_X1 U503 ( .A1(n751), .A2(KEYINPUT44), .ZN(n403) );
  INV_X1 U504 ( .A(n751), .ZN(n404) );
  XNOR2_X2 U505 ( .A(n518), .B(KEYINPUT35), .ZN(n751) );
  NAND2_X1 U506 ( .A1(n647), .A2(G469), .ZN(n412) );
  AND2_X2 U507 ( .A1(n522), .A2(n696), .ZN(n531) );
  XNOR2_X2 U508 ( .A(n413), .B(n437), .ZN(n699) );
  INV_X1 U509 ( .A(KEYINPUT48), .ZN(n414) );
  XNOR2_X1 U510 ( .A(n417), .B(KEYINPUT34), .ZN(n517) );
  XNOR2_X1 U511 ( .A(n467), .B(KEYINPUT33), .ZN(n717) );
  XOR2_X1 U512 ( .A(G110), .B(G119), .Z(n418) );
  XNOR2_X1 U513 ( .A(n442), .B(n441), .ZN(n443) );
  INV_X1 U514 ( .A(n575), .ZN(n560) );
  XOR2_X1 U515 ( .A(n444), .B(n443), .Z(n445) );
  AND2_X1 U516 ( .A1(n693), .A2(n560), .ZN(n561) );
  INV_X1 U517 ( .A(KEYINPUT22), .ZN(n520) );
  INV_X1 U518 ( .A(KEYINPUT125), .ZN(n621) );
  XNOR2_X2 U519 ( .A(G143), .B(KEYINPUT65), .ZN(n419) );
  XNOR2_X2 U520 ( .A(n419), .B(G128), .ZN(n475) );
  XNOR2_X2 U521 ( .A(n475), .B(n420), .ZN(n510) );
  XNOR2_X2 U522 ( .A(n510), .B(KEYINPUT69), .ZN(n424) );
  XNOR2_X1 U523 ( .A(n421), .B(KEYINPUT64), .ZN(n476) );
  INV_X1 U524 ( .A(G131), .ZN(n422) );
  XNOR2_X1 U525 ( .A(n476), .B(n422), .ZN(n423) );
  XNOR2_X2 U526 ( .A(n424), .B(n423), .ZN(n738) );
  XOR2_X1 U527 ( .A(KEYINPUT5), .B(KEYINPUT91), .Z(n426) );
  XNOR2_X1 U528 ( .A(G137), .B(KEYINPUT92), .ZN(n425) );
  XNOR2_X1 U529 ( .A(n426), .B(n425), .ZN(n428) );
  NOR2_X1 U530 ( .A1(G953), .A2(G237), .ZN(n493) );
  NAND2_X1 U531 ( .A1(n493), .A2(G210), .ZN(n427) );
  XNOR2_X1 U532 ( .A(n428), .B(n427), .ZN(n434) );
  XNOR2_X1 U533 ( .A(n429), .B(G101), .ZN(n431) );
  XNOR2_X1 U534 ( .A(n431), .B(n430), .ZN(n433) );
  XNOR2_X1 U535 ( .A(n434), .B(n471), .ZN(n435) );
  XNOR2_X1 U536 ( .A(n738), .B(n435), .ZN(n634) );
  INV_X1 U537 ( .A(KEYINPUT71), .ZN(n436) );
  XNOR2_X1 U538 ( .A(n436), .B(G472), .ZN(n437) );
  XOR2_X1 U539 ( .A(n468), .B(G101), .Z(n440) );
  XOR2_X1 U540 ( .A(G137), .B(KEYINPUT68), .Z(n456) );
  XNOR2_X1 U541 ( .A(G140), .B(n456), .ZN(n439) );
  XNOR2_X1 U542 ( .A(n440), .B(n439), .ZN(n444) );
  NAND2_X1 U543 ( .A1(G227), .A2(n448), .ZN(n442) );
  XNOR2_X2 U544 ( .A(n738), .B(n445), .ZN(n647) );
  NAND2_X1 U545 ( .A1(G234), .A2(n606), .ZN(n446) );
  XNOR2_X1 U546 ( .A(KEYINPUT20), .B(n446), .ZN(n461) );
  NAND2_X1 U547 ( .A1(n461), .A2(G221), .ZN(n447) );
  XNOR2_X1 U548 ( .A(n447), .B(KEYINPUT21), .ZN(n692) );
  NAND2_X1 U549 ( .A1(G234), .A2(n448), .ZN(n449) );
  XOR2_X1 U550 ( .A(KEYINPUT8), .B(n449), .Z(n511) );
  NAND2_X1 U551 ( .A1(G221), .A2(n511), .ZN(n454) );
  XNOR2_X1 U552 ( .A(n418), .B(n450), .ZN(n452) );
  XNOR2_X1 U553 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U554 ( .A(n454), .B(n453), .ZN(n458) );
  XNOR2_X1 U555 ( .A(n492), .B(n456), .ZN(n740) );
  INV_X1 U556 ( .A(n617), .ZN(n460) );
  NAND2_X1 U557 ( .A1(n460), .A2(n459), .ZN(n465) );
  NAND2_X1 U558 ( .A1(n461), .A2(G217), .ZN(n463) );
  XNOR2_X1 U559 ( .A(KEYINPUT90), .B(KEYINPUT25), .ZN(n462) );
  NOR2_X1 U560 ( .A1(n692), .A2(n693), .ZN(n696) );
  INV_X1 U561 ( .A(KEYINPUT104), .ZN(n466) );
  XNOR2_X1 U562 ( .A(n498), .B(KEYINPUT16), .ZN(n469) );
  XNOR2_X1 U563 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U564 ( .A(n471), .B(n470), .ZN(n631) );
  NAND2_X1 U565 ( .A1(n448), .A2(G224), .ZN(n472) );
  XNOR2_X1 U566 ( .A(n472), .B(KEYINPUT17), .ZN(n474) );
  XNOR2_X1 U567 ( .A(n474), .B(n473), .ZN(n478) );
  XNOR2_X1 U568 ( .A(n631), .B(n479), .ZN(n656) );
  INV_X1 U569 ( .A(G237), .ZN(n480) );
  NAND2_X1 U570 ( .A1(n459), .A2(n480), .ZN(n483) );
  NAND2_X1 U571 ( .A1(n483), .A2(G210), .ZN(n481) );
  XNOR2_X1 U572 ( .A(n481), .B(KEYINPUT88), .ZN(n482) );
  NAND2_X1 U573 ( .A1(n483), .A2(G214), .ZN(n707) );
  XOR2_X1 U574 ( .A(KEYINPUT14), .B(KEYINPUT89), .Z(n485) );
  XNOR2_X1 U575 ( .A(n485), .B(n484), .ZN(n486) );
  NAND2_X1 U576 ( .A1(G952), .A2(n486), .ZN(n724) );
  NOR2_X1 U577 ( .A1(n724), .A2(G953), .ZN(n559) );
  NAND2_X1 U578 ( .A1(G902), .A2(n486), .ZN(n556) );
  OR2_X1 U579 ( .A1(n448), .A2(G898), .ZN(n630) );
  NOR2_X1 U580 ( .A1(n556), .A2(n630), .ZN(n487) );
  OR2_X1 U581 ( .A1(n559), .A2(n487), .ZN(n488) );
  NAND2_X1 U582 ( .A1(n578), .A2(n488), .ZN(n489) );
  XNOR2_X2 U583 ( .A(n489), .B(KEYINPUT0), .ZN(n535) );
  XNOR2_X1 U584 ( .A(n360), .B(n490), .ZN(n491) );
  NAND2_X1 U585 ( .A1(G214), .A2(n493), .ZN(n494) );
  XNOR2_X1 U586 ( .A(n359), .B(n494), .ZN(n502) );
  XOR2_X1 U587 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n496) );
  XNOR2_X1 U588 ( .A(n496), .B(n495), .ZN(n500) );
  XOR2_X1 U589 ( .A(G143), .B(G131), .Z(n497) );
  XNOR2_X1 U590 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U591 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U592 ( .A(n502), .B(n501), .ZN(n642) );
  NAND2_X1 U593 ( .A1(n642), .A2(n459), .ZN(n506) );
  XOR2_X1 U594 ( .A(KEYINPUT13), .B(KEYINPUT99), .Z(n504) );
  XNOR2_X1 U595 ( .A(KEYINPUT98), .B(G475), .ZN(n503) );
  XNOR2_X1 U596 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U597 ( .A(n506), .B(n505), .ZN(n539) );
  XNOR2_X1 U598 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U599 ( .A(n510), .B(n509), .ZN(n515) );
  XOR2_X1 U600 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n513) );
  NAND2_X1 U601 ( .A1(G217), .A2(n511), .ZN(n512) );
  XNOR2_X1 U602 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U603 ( .A(n515), .B(n514), .ZN(n734) );
  XNOR2_X1 U604 ( .A(G478), .B(n358), .ZN(n540) );
  INV_X1 U605 ( .A(n540), .ZN(n537) );
  OR2_X1 U606 ( .A1(n539), .A2(n537), .ZN(n571) );
  INV_X1 U607 ( .A(n571), .ZN(n516) );
  NAND2_X1 U608 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U609 ( .A1(n539), .A2(n537), .ZN(n584) );
  INV_X1 U610 ( .A(n692), .ZN(n552) );
  NAND2_X1 U611 ( .A1(n584), .A2(n552), .ZN(n519) );
  XNOR2_X1 U612 ( .A(n521), .B(n520), .ZN(n527) );
  INV_X1 U613 ( .A(n369), .ZN(n594) );
  XNOR2_X1 U614 ( .A(n543), .B(n523), .ZN(n525) );
  BUF_X1 U615 ( .A(n699), .Z(n566) );
  NOR2_X1 U616 ( .A1(n566), .A2(n576), .ZN(n524) );
  NAND2_X1 U617 ( .A1(n525), .A2(n524), .ZN(n625) );
  NOR2_X1 U618 ( .A1(n594), .A2(n576), .ZN(n526) );
  NAND2_X1 U619 ( .A1(n526), .A2(n553), .ZN(n528) );
  NOR2_X1 U620 ( .A1(n528), .A2(n527), .ZN(n530) );
  XOR2_X1 U621 ( .A(KEYINPUT74), .B(KEYINPUT32), .Z(n529) );
  XNOR2_X1 U622 ( .A(n530), .B(n529), .ZN(n623) );
  BUF_X1 U623 ( .A(n531), .Z(n532) );
  NAND2_X1 U624 ( .A1(n566), .A2(n532), .ZN(n703) );
  NOR2_X1 U625 ( .A1(n535), .A2(n703), .ZN(n534) );
  XNOR2_X1 U626 ( .A(KEYINPUT31), .B(KEYINPUT93), .ZN(n533) );
  XNOR2_X1 U627 ( .A(n534), .B(n533), .ZN(n680) );
  OR2_X1 U628 ( .A1(n568), .A2(n566), .ZN(n536) );
  NOR2_X1 U629 ( .A1(n536), .A2(n535), .ZN(n669) );
  NOR2_X1 U630 ( .A1(n680), .A2(n669), .ZN(n541) );
  INV_X1 U631 ( .A(n539), .ZN(n538) );
  XOR2_X1 U632 ( .A(KEYINPUT101), .B(n679), .Z(n598) );
  NOR2_X1 U633 ( .A1(n598), .A2(n592), .ZN(n713) );
  NOR2_X1 U634 ( .A1(n541), .A2(n713), .ZN(n542) );
  XNOR2_X1 U635 ( .A(n542), .B(KEYINPUT102), .ZN(n546) );
  INV_X1 U636 ( .A(n543), .ZN(n545) );
  NAND2_X1 U637 ( .A1(n553), .A2(n576), .ZN(n544) );
  NOR2_X1 U638 ( .A1(n545), .A2(n544), .ZN(n624) );
  NOR2_X1 U639 ( .A1(n546), .A2(n624), .ZN(n547) );
  NAND2_X1 U640 ( .A1(n611), .A2(n549), .ZN(n551) );
  INV_X1 U641 ( .A(KEYINPUT78), .ZN(n550) );
  XNOR2_X1 U642 ( .A(n551), .B(n550), .ZN(n605) );
  INV_X1 U643 ( .A(n553), .ZN(n554) );
  OR2_X1 U644 ( .A1(n448), .A2(n556), .ZN(n557) );
  NOR2_X1 U645 ( .A1(G900), .A2(n557), .ZN(n558) );
  NOR2_X1 U646 ( .A1(n559), .A2(n558), .ZN(n575) );
  INV_X1 U647 ( .A(n562), .ZN(n563) );
  NAND2_X1 U648 ( .A1(n593), .A2(n563), .ZN(n564) );
  XNOR2_X1 U649 ( .A(n564), .B(KEYINPUT36), .ZN(n565) );
  NOR2_X1 U650 ( .A1(n594), .A2(n565), .ZN(n682) );
  NAND2_X1 U651 ( .A1(n699), .A2(n707), .ZN(n567) );
  NOR2_X1 U652 ( .A1(n575), .A2(n568), .ZN(n569) );
  XNOR2_X1 U653 ( .A(n569), .B(KEYINPUT73), .ZN(n570) );
  NOR2_X1 U654 ( .A1(n571), .A2(n562), .ZN(n572) );
  NAND2_X1 U655 ( .A1(n713), .A2(KEYINPUT47), .ZN(n573) );
  NAND2_X1 U656 ( .A1(n750), .A2(n573), .ZN(n574) );
  XNOR2_X1 U657 ( .A(n574), .B(KEYINPUT75), .ZN(n583) );
  XNOR2_X1 U658 ( .A(n577), .B(KEYINPUT108), .ZN(n588) );
  INV_X1 U659 ( .A(n588), .ZN(n579) );
  NAND2_X1 U660 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U661 ( .A(n580), .B(KEYINPUT47), .ZN(n582) );
  INV_X1 U662 ( .A(n580), .ZN(n674) );
  NAND2_X1 U663 ( .A1(n674), .A2(n713), .ZN(n581) );
  INV_X1 U664 ( .A(n584), .ZN(n711) );
  XNOR2_X1 U665 ( .A(KEYINPUT72), .B(KEYINPUT38), .ZN(n585) );
  XNOR2_X1 U666 ( .A(n562), .B(n585), .ZN(n708) );
  NAND2_X1 U667 ( .A1(n708), .A2(n707), .ZN(n714) );
  NOR2_X1 U668 ( .A1(n711), .A2(n714), .ZN(n587) );
  XOR2_X1 U669 ( .A(KEYINPUT109), .B(KEYINPUT41), .Z(n586) );
  XNOR2_X1 U670 ( .A(n587), .B(n586), .ZN(n726) );
  NOR2_X1 U671 ( .A1(n726), .A2(n588), .ZN(n589) );
  XNOR2_X1 U672 ( .A(n589), .B(KEYINPUT42), .ZN(n755) );
  XOR2_X1 U673 ( .A(KEYINPUT83), .B(KEYINPUT39), .Z(n591) );
  NAND2_X1 U674 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U675 ( .A(KEYINPUT43), .B(n595), .ZN(n596) );
  NAND2_X1 U676 ( .A1(n596), .A2(n562), .ZN(n597) );
  XNOR2_X1 U677 ( .A(n597), .B(KEYINPUT106), .ZN(n748) );
  INV_X1 U678 ( .A(n748), .ZN(n602) );
  NAND2_X1 U679 ( .A1(n599), .A2(n598), .ZN(n601) );
  INV_X1 U680 ( .A(KEYINPUT110), .ZN(n600) );
  XNOR2_X1 U681 ( .A(n601), .B(n600), .ZN(n754) );
  NOR2_X1 U682 ( .A1(n602), .A2(n754), .ZN(n603) );
  NAND2_X1 U683 ( .A1(n605), .A2(n741), .ZN(n609) );
  XOR2_X1 U684 ( .A(KEYINPUT80), .B(n606), .Z(n607) );
  NAND2_X1 U685 ( .A1(n607), .A2(KEYINPUT2), .ZN(n608) );
  NAND2_X1 U686 ( .A1(n609), .A2(n608), .ZN(n614) );
  XNOR2_X1 U687 ( .A(n610), .B(KEYINPUT81), .ZN(n613) );
  BUF_X1 U688 ( .A(n611), .Z(n612) );
  NAND2_X1 U689 ( .A1(n613), .A2(n612), .ZN(n688) );
  INV_X1 U690 ( .A(KEYINPUT66), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n368), .A2(G217), .ZN(n618) );
  XNOR2_X1 U692 ( .A(n618), .B(n617), .ZN(n620) );
  INV_X1 U693 ( .A(G952), .ZN(n619) );
  AND2_X1 U694 ( .A1(n619), .A2(G953), .ZN(n737) );
  NOR2_X2 U695 ( .A1(n620), .A2(n737), .ZN(n622) );
  XNOR2_X1 U696 ( .A(n622), .B(n621), .ZN(G66) );
  XNOR2_X1 U697 ( .A(n623), .B(G119), .ZN(G21) );
  XOR2_X1 U698 ( .A(G101), .B(n624), .Z(G3) );
  XNOR2_X1 U699 ( .A(n625), .B(G110), .ZN(G12) );
  NAND2_X1 U700 ( .A1(n612), .A2(n448), .ZN(n629) );
  NAND2_X1 U701 ( .A1(G953), .A2(G224), .ZN(n626) );
  XNOR2_X1 U702 ( .A(KEYINPUT61), .B(n626), .ZN(n627) );
  NAND2_X1 U703 ( .A1(n627), .A2(G898), .ZN(n628) );
  NAND2_X1 U704 ( .A1(n629), .A2(n628), .ZN(n633) );
  NAND2_X1 U705 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U706 ( .A(n633), .B(n632), .Z(G69) );
  NAND2_X1 U707 ( .A1(n367), .A2(G472), .ZN(n636) );
  XNOR2_X1 U708 ( .A(KEYINPUT86), .B(KEYINPUT63), .ZN(n638) );
  XOR2_X1 U709 ( .A(n638), .B(KEYINPUT84), .Z(n639) );
  XNOR2_X1 U710 ( .A(n640), .B(n639), .ZN(G57) );
  NAND2_X1 U711 ( .A1(n368), .A2(G475), .ZN(n644) );
  XOR2_X1 U712 ( .A(KEYINPUT67), .B(KEYINPUT59), .Z(n641) );
  XNOR2_X1 U713 ( .A(n646), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U714 ( .A1(n733), .A2(G469), .ZN(n653) );
  XNOR2_X1 U715 ( .A(n647), .B(KEYINPUT122), .ZN(n651) );
  XOR2_X1 U716 ( .A(KEYINPUT121), .B(KEYINPUT123), .Z(n649) );
  XNOR2_X1 U717 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n648) );
  XNOR2_X1 U718 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U719 ( .A(n655), .B(KEYINPUT124), .ZN(G54) );
  NAND2_X1 U720 ( .A1(n733), .A2(G210), .ZN(n661) );
  XNOR2_X1 U721 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n658) );
  XNOR2_X1 U722 ( .A(KEYINPUT55), .B(KEYINPUT85), .ZN(n657) );
  XNOR2_X1 U723 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U724 ( .A(KEYINPUT82), .B(KEYINPUT56), .ZN(n663) );
  XNOR2_X1 U725 ( .A(n664), .B(n663), .ZN(G51) );
  NAND2_X1 U726 ( .A1(n676), .A2(n669), .ZN(n665) );
  XNOR2_X1 U727 ( .A(n665), .B(G104), .ZN(G6) );
  XOR2_X1 U728 ( .A(KEYINPUT112), .B(KEYINPUT27), .Z(n667) );
  XNOR2_X1 U729 ( .A(G107), .B(KEYINPUT26), .ZN(n666) );
  XNOR2_X1 U730 ( .A(n667), .B(n666), .ZN(n668) );
  XOR2_X1 U731 ( .A(KEYINPUT111), .B(n668), .Z(n671) );
  NAND2_X1 U732 ( .A1(n669), .A2(n679), .ZN(n670) );
  XNOR2_X1 U733 ( .A(n671), .B(n670), .ZN(G9) );
  XOR2_X1 U734 ( .A(G128), .B(KEYINPUT29), .Z(n673) );
  NAND2_X1 U735 ( .A1(n674), .A2(n679), .ZN(n672) );
  XNOR2_X1 U736 ( .A(n673), .B(n672), .ZN(G30) );
  NAND2_X1 U737 ( .A1(n674), .A2(n676), .ZN(n675) );
  XNOR2_X1 U738 ( .A(n675), .B(G146), .ZN(G48) );
  XOR2_X1 U739 ( .A(G113), .B(KEYINPUT113), .Z(n678) );
  NAND2_X1 U740 ( .A1(n676), .A2(n680), .ZN(n677) );
  XNOR2_X1 U741 ( .A(n678), .B(n677), .ZN(G15) );
  NAND2_X1 U742 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U743 ( .A(n681), .B(G116), .ZN(G18) );
  XNOR2_X1 U744 ( .A(G125), .B(n682), .ZN(n683) );
  XNOR2_X1 U745 ( .A(n683), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U746 ( .A(KEYINPUT2), .B(KEYINPUT76), .ZN(n684) );
  OR2_X1 U747 ( .A1(n612), .A2(n684), .ZN(n687) );
  XNOR2_X1 U748 ( .A(n685), .B(KEYINPUT77), .ZN(n686) );
  NAND2_X1 U749 ( .A1(n687), .A2(n686), .ZN(n690) );
  INV_X1 U750 ( .A(n688), .ZN(n689) );
  XNOR2_X1 U751 ( .A(KEYINPUT79), .B(n691), .ZN(n730) );
  NAND2_X1 U752 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U753 ( .A(n694), .B(KEYINPUT115), .ZN(n695) );
  XNOR2_X1 U754 ( .A(KEYINPUT49), .B(n695), .ZN(n701) );
  NOR2_X1 U755 ( .A1(n696), .A2(n369), .ZN(n697) );
  XNOR2_X1 U756 ( .A(n697), .B(KEYINPUT50), .ZN(n698) );
  NOR2_X1 U757 ( .A1(n566), .A2(n698), .ZN(n700) );
  NAND2_X1 U758 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U759 ( .A(n702), .B(KEYINPUT116), .ZN(n704) );
  NAND2_X1 U760 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U761 ( .A(KEYINPUT51), .B(n705), .ZN(n706) );
  NOR2_X1 U762 ( .A1(n726), .A2(n706), .ZN(n720) );
  NOR2_X1 U763 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U764 ( .A(KEYINPUT117), .B(n709), .Z(n710) );
  NOR2_X1 U765 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U766 ( .A(n712), .B(KEYINPUT118), .ZN(n716) );
  NOR2_X1 U767 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U768 ( .A1(n716), .A2(n715), .ZN(n718) );
  BUF_X1 U769 ( .A(n717), .Z(n725) );
  NOR2_X1 U770 ( .A1(n718), .A2(n725), .ZN(n719) );
  NOR2_X1 U771 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U772 ( .A(n721), .B(KEYINPUT52), .Z(n722) );
  XNOR2_X1 U773 ( .A(KEYINPUT119), .B(n722), .ZN(n723) );
  NOR2_X1 U774 ( .A1(n724), .A2(n723), .ZN(n728) );
  NOR2_X1 U775 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U776 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U777 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U778 ( .A(n732), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U779 ( .A1(n367), .A2(G478), .ZN(n735) );
  XNOR2_X1 U780 ( .A(n735), .B(n734), .ZN(n736) );
  NOR2_X1 U781 ( .A1(n737), .A2(n736), .ZN(G63) );
  XOR2_X1 U782 ( .A(n738), .B(KEYINPUT126), .Z(n739) );
  XOR2_X1 U783 ( .A(n740), .B(n739), .Z(n743) );
  XOR2_X1 U784 ( .A(n743), .B(n741), .Z(n742) );
  NAND2_X1 U785 ( .A1(n742), .A2(n448), .ZN(n747) );
  XNOR2_X1 U786 ( .A(G227), .B(n743), .ZN(n744) );
  NAND2_X1 U787 ( .A1(n744), .A2(G900), .ZN(n745) );
  NAND2_X1 U788 ( .A1(G953), .A2(n745), .ZN(n746) );
  NAND2_X1 U789 ( .A1(n747), .A2(n746), .ZN(G72) );
  XNOR2_X1 U790 ( .A(G140), .B(n748), .ZN(n749) );
  XNOR2_X1 U791 ( .A(n749), .B(KEYINPUT114), .ZN(G42) );
  XNOR2_X1 U792 ( .A(n750), .B(G143), .ZN(G45) );
  BUF_X1 U793 ( .A(n751), .Z(n752) );
  XOR2_X1 U794 ( .A(n752), .B(G122), .Z(G24) );
  XOR2_X1 U795 ( .A(G131), .B(n753), .Z(G33) );
  XOR2_X1 U796 ( .A(G134), .B(n754), .Z(G36) );
  XOR2_X1 U797 ( .A(G137), .B(n755), .Z(G39) );
endmodule

