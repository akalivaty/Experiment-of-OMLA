//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1 0 1 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n438, new_n449, new_n452, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n571,
    new_n573, new_n574, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n589, new_n590, new_n592, new_n593, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n635, new_n636, new_n639,
    new_n641, new_n642, new_n643, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1206;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  OR2_X1    g011(.A1(new_n436), .A2(KEYINPUT65), .ZN(new_n437));
  NAND2_X1  g012(.A1(new_n436), .A2(KEYINPUT65), .ZN(new_n438));
  NAND2_X1  g013(.A1(new_n437), .A2(new_n438), .ZN(G220));
  INV_X1    g014(.A(G96), .ZN(G221));
  INV_X1    g015(.A(G69), .ZN(G235));
  INV_X1    g016(.A(G120), .ZN(G236));
  INV_X1    g017(.A(G57), .ZN(G237));
  INV_X1    g018(.A(G108), .ZN(G238));
  NAND4_X1  g019(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT66), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XOR2_X1   g029(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n455));
  XNOR2_X1  g030(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n456), .A2(G2106), .ZN(new_n461));
  INV_X1    g036(.A(G567), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n461), .B1(new_n462), .B2(new_n457), .ZN(new_n463));
  XOR2_X1   g038(.A(new_n463), .B(KEYINPUT68), .Z(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(G125), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(KEYINPUT69), .B1(new_n472), .B2(G2105), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n474), .A2(new_n466), .A3(G2104), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n473), .A2(new_n475), .A3(G101), .ZN(new_n476));
  OAI211_X1 g051(.A(G137), .B(new_n466), .C1(new_n467), .C2(new_n468), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n471), .A2(new_n478), .ZN(G160));
  OR2_X1    g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  MUX2_X1   g059(.A(G100), .B(G112), .S(G2105), .Z(new_n485));
  AOI22_X1  g060(.A1(new_n484), .A2(G124), .B1(G2104), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(G2105), .B1(new_n480), .B2(new_n481), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  INV_X1    g065(.A(KEYINPUT71), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n491), .A2(new_n466), .A3(KEYINPUT4), .A4(G138), .ZN(new_n492));
  NAND2_X1  g067(.A1(G126), .A2(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(new_n482), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT70), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n496), .B1(new_n466), .B2(G114), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n498), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n499));
  OR2_X1    g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n497), .A2(new_n499), .A3(new_n500), .A4(G2104), .ZN(new_n501));
  OAI211_X1 g076(.A(G138), .B(new_n466), .C1(new_n467), .C2(new_n468), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n504), .A2(KEYINPUT71), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n495), .B(new_n501), .C1(new_n503), .C2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  NAND2_X1  g082(.A1(KEYINPUT73), .A2(G543), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(KEYINPUT76), .A3(G62), .ZN(new_n513));
  INV_X1    g088(.A(G75), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g091(.A(KEYINPUT76), .B1(new_n512), .B2(G62), .ZN(new_n517));
  OAI21_X1  g092(.A(G651), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AND2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  OAI211_X1 g095(.A(G50), .B(G543), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n521), .B(new_n522), .ZN(new_n523));
  AND3_X1   g098(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n524));
  AOI21_X1  g099(.A(KEYINPUT5), .B1(KEYINPUT73), .B2(G543), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n524), .A2(new_n525), .B1(new_n519), .B2(new_n520), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT74), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT6), .B(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n512), .A2(KEYINPUT74), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n528), .A2(G88), .A3(new_n530), .ZN(new_n531));
  AND3_X1   g106(.A1(new_n523), .A2(new_n531), .A3(KEYINPUT75), .ZN(new_n532));
  AOI21_X1  g107(.A(KEYINPUT75), .B1(new_n523), .B2(new_n531), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n518), .B1(new_n532), .B2(new_n533), .ZN(G303));
  INV_X1    g109(.A(G303), .ZN(G166));
  INV_X1    g110(.A(new_n520), .ZN(new_n536));
  NAND2_X1  g111(.A1(KEYINPUT6), .A2(G651), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n515), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AND2_X1   g113(.A1(G63), .A2(G651), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n538), .A2(G51), .B1(new_n512), .B2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n528), .A2(G89), .A3(new_n530), .ZN(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT7), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT77), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n542), .A2(KEYINPUT77), .A3(new_n544), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n541), .B1(new_n547), .B2(new_n548), .ZN(G168));
  NAND2_X1  g124(.A1(new_n528), .A2(new_n530), .ZN(new_n550));
  INV_X1    g125(.A(G90), .ZN(new_n551));
  INV_X1    g126(.A(G52), .ZN(new_n552));
  INV_X1    g127(.A(new_n538), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n550), .A2(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(KEYINPUT78), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT78), .ZN(new_n556));
  OAI221_X1 g131(.A(new_n556), .B1(new_n552), .B2(new_n553), .C1(new_n550), .C2(new_n551), .ZN(new_n557));
  NAND2_X1  g132(.A1(G77), .A2(G543), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n524), .A2(new_n525), .ZN(new_n559));
  INV_X1    g134(.A(G64), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n555), .A2(new_n557), .B1(G651), .B2(new_n561), .ZN(G171));
  NAND2_X1  g137(.A1(G68), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G56), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n559), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n565), .A2(G651), .B1(G43), .B2(new_n538), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n528), .A2(G81), .A3(new_n530), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(G153));
  AND3_X1   g145(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G36), .ZN(G176));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT8), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n571), .A2(new_n574), .ZN(G188));
  NAND3_X1  g150(.A1(new_n528), .A2(G91), .A3(new_n530), .ZN(new_n576));
  OAI211_X1 g151(.A(G53), .B(G543), .C1(new_n519), .C2(new_n520), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(KEYINPUT79), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT79), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n529), .A2(new_n579), .A3(G53), .A4(G543), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n580), .A3(KEYINPUT9), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT9), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n577), .A2(KEYINPUT79), .A3(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(G65), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n584), .B1(new_n510), .B2(new_n511), .ZN(new_n585));
  AND2_X1   g160(.A1(G78), .A2(G543), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n576), .A2(new_n581), .A3(new_n583), .A4(new_n587), .ZN(G299));
  NAND2_X1  g163(.A1(new_n555), .A2(new_n557), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n561), .A2(G651), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(G301));
  INV_X1    g166(.A(KEYINPUT80), .ZN(new_n592));
  NAND2_X1  g167(.A1(G168), .A2(new_n592), .ZN(new_n593));
  AND3_X1   g168(.A1(new_n542), .A2(KEYINPUT77), .A3(new_n544), .ZN(new_n594));
  AOI21_X1  g169(.A(KEYINPUT77), .B1(new_n542), .B2(new_n544), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n540), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(KEYINPUT80), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G286));
  NAND3_X1  g174(.A1(new_n528), .A2(G87), .A3(new_n530), .ZN(new_n600));
  INV_X1    g175(.A(G74), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n559), .A2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(G651), .B1(new_n538), .B2(G49), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n600), .A2(new_n603), .ZN(G288));
  OAI211_X1 g179(.A(G48), .B(G543), .C1(new_n519), .C2(new_n520), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(G73), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G61), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n559), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n606), .B1(new_n609), .B2(G651), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n528), .A2(G86), .A3(new_n530), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(G305));
  AOI22_X1  g187(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n613));
  INV_X1    g188(.A(G651), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n528), .A2(G85), .A3(new_n530), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT81), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n538), .A2(G47), .ZN(new_n618));
  AND3_X1   g193(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n617), .B1(new_n616), .B2(new_n618), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n615), .B1(new_n619), .B2(new_n620), .ZN(G290));
  NAND2_X1  g196(.A1(new_n538), .A2(G54), .ZN(new_n622));
  XOR2_X1   g197(.A(KEYINPUT82), .B(G66), .Z(new_n623));
  AOI22_X1  g198(.A1(new_n623), .A2(new_n512), .B1(G79), .B2(G543), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n622), .B1(new_n624), .B2(new_n614), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT10), .ZN(new_n626));
  INV_X1    g201(.A(G92), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n550), .B2(new_n627), .ZN(new_n628));
  NAND4_X1  g203(.A1(new_n528), .A2(new_n530), .A3(KEYINPUT10), .A4(G92), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n625), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n632), .B1(G868), .B2(G171), .ZN(G284));
  AOI21_X1  g208(.A(new_n632), .B1(G868), .B2(G171), .ZN(G321));
  INV_X1    g209(.A(G868), .ZN(new_n635));
  NAND2_X1  g210(.A1(G299), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(new_n598), .B2(new_n635), .ZN(G297));
  OAI21_X1  g212(.A(new_n636), .B1(new_n598), .B2(new_n635), .ZN(G280));
  INV_X1    g213(.A(G559), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n630), .B1(new_n639), .B2(G860), .ZN(G148));
  NAND2_X1  g215(.A1(new_n568), .A2(new_n635), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n630), .A2(new_n639), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT83), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n641), .B1(new_n643), .B2(new_n635), .ZN(G323));
  XNOR2_X1  g219(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g220(.A1(new_n473), .A2(new_n475), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(new_n482), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT12), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT13), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n650), .A2(G2100), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n484), .A2(G123), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT84), .ZN(new_n653));
  MUX2_X1   g228(.A(G99), .B(G111), .S(G2105), .Z(new_n654));
  AOI22_X1  g229(.A1(G135), .A2(new_n487), .B1(new_n654), .B2(G2104), .ZN(new_n655));
  AND2_X1   g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2096), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n650), .A2(G2100), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n651), .A2(new_n657), .A3(new_n658), .ZN(G156));
  XNOR2_X1  g234(.A(G2451), .B(G2454), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT16), .ZN(new_n661));
  XOR2_X1   g236(.A(G2443), .B(G2446), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G1341), .B(G1348), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT15), .B(G2435), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT86), .B(G2438), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2427), .B(G2430), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT85), .B(KEYINPUT14), .Z(new_n672));
  NAND3_X1  g247(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n665), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n665), .A2(new_n673), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n674), .A2(G14), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT87), .Z(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(G401));
  XOR2_X1   g253(.A(G2084), .B(G2090), .Z(new_n679));
  XNOR2_X1  g254(.A(G2072), .B(G2078), .ZN(new_n680));
  XNOR2_X1  g255(.A(G2067), .B(G2678), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT18), .Z(new_n683));
  INV_X1    g258(.A(new_n679), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n680), .A2(KEYINPUT17), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(new_n681), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(new_n684), .B2(new_n685), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n679), .A2(new_n681), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n680), .B1(new_n689), .B2(KEYINPUT17), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n683), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(G2096), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(G2100), .ZN(G227));
  XOR2_X1   g268(.A(G1956), .B(G2474), .Z(new_n694));
  XOR2_X1   g269(.A(G1961), .B(G1966), .Z(new_n695));
  AND2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT89), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1971), .B(G1976), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT90), .B(KEYINPUT20), .Z(new_n702));
  OR2_X1    g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n694), .A2(new_n695), .ZN(new_n705));
  NOR3_X1   g280(.A1(new_n700), .A2(new_n696), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(new_n700), .B2(new_n705), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n703), .A2(new_n704), .A3(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT91), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n708), .B(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(G1991), .B(G1996), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1981), .B(G1986), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n711), .B(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(G229));
  XOR2_X1   g291(.A(KEYINPUT93), .B(G16), .Z(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(G166), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G22), .B2(new_n718), .ZN(new_n720));
  INV_X1    g295(.A(G1971), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n720), .A2(new_n721), .ZN(new_n723));
  NOR2_X1   g298(.A1(G6), .A2(G16), .ZN(new_n724));
  INV_X1    g299(.A(G305), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n724), .B1(new_n725), .B2(G16), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT32), .B(G1981), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n726), .B(new_n727), .Z(new_n728));
  INV_X1    g303(.A(G16), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G23), .ZN(new_n730));
  INV_X1    g305(.A(G288), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(new_n729), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT33), .B(G1976), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT95), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n732), .B(new_n734), .Z(new_n735));
  NAND4_X1  g310(.A1(new_n722), .A2(new_n723), .A3(new_n728), .A4(new_n735), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n736), .A2(KEYINPUT34), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(KEYINPUT34), .ZN(new_n738));
  NOR2_X1   g313(.A1(G25), .A2(G29), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n487), .A2(G131), .ZN(new_n740));
  AND2_X1   g315(.A1(G107), .A2(G2105), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G95), .B2(new_n466), .ZN(new_n742));
  INV_X1    g317(.A(G119), .ZN(new_n743));
  OAI221_X1 g318(.A(new_n740), .B1(new_n472), .B2(new_n742), .C1(new_n743), .C2(new_n483), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT92), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n744), .A2(new_n745), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n739), .B1(new_n749), .B2(G29), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT35), .B(G1991), .Z(new_n751));
  XOR2_X1   g326(.A(new_n750), .B(new_n751), .Z(new_n752));
  OR2_X1    g327(.A1(new_n718), .A2(G24), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G290), .B2(new_n717), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT94), .B(G1986), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n754), .A2(new_n755), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n752), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n737), .A2(new_n738), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(KEYINPUT36), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT36), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n737), .A2(new_n761), .A3(new_n738), .A4(new_n758), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n717), .A2(G20), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT23), .ZN(new_n765));
  INV_X1    g340(.A(G299), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n765), .B1(new_n766), .B2(new_n729), .ZN(new_n767));
  INV_X1    g342(.A(G1956), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(G29), .A2(G35), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G162), .B2(G29), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT29), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G2090), .ZN(new_n773));
  MUX2_X1   g348(.A(G104), .B(G116), .S(G2105), .Z(new_n774));
  AOI22_X1  g349(.A1(new_n484), .A2(G128), .B1(G2104), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n487), .A2(G140), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n777), .A2(G29), .ZN(new_n778));
  INV_X1    g353(.A(G29), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(G26), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT28), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G2067), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n718), .A2(G19), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n569), .B2(new_n718), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1341), .ZN(new_n786));
  INV_X1    g361(.A(G1348), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n630), .A2(G16), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G4), .B2(G16), .ZN(new_n789));
  AOI211_X1 g364(.A(new_n783), .B(new_n786), .C1(new_n787), .C2(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n787), .B2(new_n789), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT96), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n769), .B(new_n773), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n792), .B2(new_n791), .ZN(new_n794));
  NOR2_X1   g369(.A1(G5), .A2(G16), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G171), .B2(G16), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT98), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n797), .A2(G1961), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT99), .Z(new_n799));
  NOR2_X1   g374(.A1(G29), .A2(G33), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT97), .Z(new_n801));
  NAND3_X1  g376(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT25), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n802), .A2(new_n803), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n804), .A2(new_n805), .B1(new_n487), .B2(G139), .ZN(new_n806));
  NAND2_X1  g381(.A1(G115), .A2(G2104), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n467), .A2(new_n468), .ZN(new_n808));
  INV_X1    g383(.A(G127), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n810), .A2(G2105), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n806), .A2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n801), .B1(new_n813), .B2(new_n779), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(G2072), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n779), .A2(G32), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n484), .A2(G129), .B1(G141), .B2(new_n487), .ZN(new_n817));
  NAND3_X1  g392(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT26), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(G105), .B2(new_n646), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n816), .B1(new_n821), .B2(G29), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT27), .B(G1996), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT31), .B(G11), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT30), .B(G28), .Z(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(G29), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(new_n656), .B2(G29), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n815), .A2(new_n824), .A3(new_n828), .ZN(new_n829));
  OR2_X1    g404(.A1(KEYINPUT24), .A2(G34), .ZN(new_n830));
  NAND2_X1  g405(.A1(KEYINPUT24), .A2(G34), .ZN(new_n831));
  AOI21_X1  g406(.A(G29), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(G160), .B2(G29), .ZN(new_n833));
  INV_X1    g408(.A(G2084), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n822), .B2(new_n823), .ZN(new_n836));
  NOR2_X1   g411(.A1(G27), .A2(G29), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(G164), .B2(G29), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(G2078), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n829), .A2(new_n836), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n729), .A2(G21), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(G168), .B2(new_n729), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(G1966), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n797), .A2(G1961), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n842), .A2(G1966), .ZN(new_n846));
  NOR3_X1   g421(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  AND3_X1   g422(.A1(new_n799), .A2(KEYINPUT100), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(KEYINPUT100), .B1(new_n799), .B2(new_n847), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n763), .B(new_n794), .C1(new_n848), .C2(new_n849), .ZN(G150));
  INV_X1    g425(.A(G150), .ZN(G311));
  NAND3_X1  g426(.A1(new_n528), .A2(G93), .A3(new_n530), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n538), .A2(G55), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(KEYINPUT101), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT101), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n852), .A2(new_n856), .A3(new_n853), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(G80), .A2(G543), .ZN(new_n859));
  INV_X1    g434(.A(G67), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n859), .B1(new_n559), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(G651), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n566), .A2(KEYINPUT102), .A3(new_n567), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n858), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  AOI22_X1  g440(.A1(new_n855), .A2(new_n857), .B1(G651), .B2(new_n861), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT102), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n568), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(new_n863), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n865), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n630), .A2(G559), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT38), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n871), .B(new_n873), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n874), .A2(KEYINPUT39), .ZN(new_n875));
  INV_X1    g450(.A(G860), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(KEYINPUT39), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n866), .A2(new_n876), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT37), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(G145));
  XNOR2_X1  g456(.A(new_n821), .B(new_n812), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n748), .A2(new_n648), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n484), .A2(G130), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n487), .A2(G142), .ZN(new_n885));
  MUX2_X1   g460(.A(G106), .B(G118), .S(G2105), .Z(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(G2104), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n884), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n748), .A2(new_n648), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n883), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n889), .B1(new_n883), .B2(new_n890), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n777), .B(G164), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NOR3_X1   g470(.A1(new_n892), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n883), .A2(new_n890), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(new_n888), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n894), .B1(new_n898), .B2(new_n891), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n882), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n489), .B(G160), .Z(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n656), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n895), .B1(new_n892), .B2(new_n893), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n898), .A2(new_n891), .A3(new_n894), .ZN(new_n904));
  INV_X1    g479(.A(new_n882), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n900), .A2(new_n902), .A3(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(G37), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n902), .B1(new_n900), .B2(new_n906), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g487(.A1(new_n866), .A2(new_n635), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(G303), .A2(G305), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n725), .B(new_n518), .C1(new_n532), .C2(new_n533), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(G290), .A2(G288), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n731), .B(new_n615), .C1(new_n619), .C2(new_n620), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n917), .A2(new_n920), .A3(KEYINPUT105), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT105), .B1(new_n917), .B2(new_n920), .ZN(new_n922));
  OAI22_X1  g497(.A1(new_n921), .A2(new_n922), .B1(new_n920), .B2(new_n917), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(KEYINPUT42), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n871), .B(new_n643), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n630), .A2(G299), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n630), .A2(G299), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n926), .B1(KEYINPUT103), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT103), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n630), .A2(new_n929), .A3(G299), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n925), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n926), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT41), .B1(new_n933), .B2(new_n927), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n927), .A2(KEYINPUT103), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n935), .A2(new_n933), .A3(KEYINPUT41), .A4(new_n930), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT104), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n928), .A2(KEYINPUT104), .A3(KEYINPUT41), .A4(new_n930), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n934), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n932), .B1(new_n940), .B2(new_n925), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n924), .B(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n914), .B1(new_n942), .B2(G868), .ZN(G295));
  AOI21_X1  g518(.A(new_n914), .B1(new_n942), .B2(G868), .ZN(G331));
  XOR2_X1   g519(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n945));
  NAND3_X1  g520(.A1(new_n593), .A2(new_n597), .A3(G171), .ZN(new_n946));
  NAND2_X1  g521(.A1(G301), .A2(G168), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n871), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n946), .A2(new_n870), .A3(new_n947), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(new_n931), .A3(new_n950), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n946), .A2(new_n870), .A3(new_n947), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n870), .B1(new_n946), .B2(new_n947), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n923), .B(new_n951), .C1(new_n940), .C2(new_n954), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n955), .A2(new_n908), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n933), .A2(new_n927), .ZN(new_n957));
  OAI211_X1 g532(.A(KEYINPUT41), .B(new_n957), .C1(new_n952), .C2(new_n953), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT41), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n959), .B1(new_n949), .B2(new_n950), .ZN(new_n960));
  INV_X1    g535(.A(new_n931), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n923), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n962), .A2(KEYINPUT108), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n956), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT108), .B1(new_n962), .B2(new_n963), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n945), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n951), .B1(new_n940), .B2(new_n954), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n963), .ZN(new_n969));
  INV_X1    g544(.A(new_n945), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n956), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  XOR2_X1   g546(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n972));
  NAND3_X1  g547(.A1(new_n967), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT43), .B1(new_n965), .B2(new_n966), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n969), .A2(new_n908), .A3(new_n955), .A4(new_n945), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n974), .A2(KEYINPUT44), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n973), .A2(new_n976), .ZN(G397));
  INV_X1    g552(.A(G1384), .ZN(new_n978));
  INV_X1    g553(.A(new_n493), .ZN(new_n979));
  INV_X1    g554(.A(G138), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n980), .A2(G2105), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n979), .B1(new_n505), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n501), .B1(new_n982), .B2(new_n808), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n505), .B1(new_n487), .B2(G138), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n978), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT45), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G40), .ZN(new_n989));
  NOR3_X1   g564(.A1(new_n471), .A2(new_n478), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  XOR2_X1   g566(.A(new_n991), .B(KEYINPUT110), .Z(new_n992));
  XNOR2_X1  g567(.A(new_n777), .B(G2067), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n991), .A2(G1996), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n992), .A2(new_n821), .ZN(new_n997));
  INV_X1    g572(.A(G1996), .ZN(new_n998));
  OAI221_X1 g573(.A(new_n994), .B1(new_n821), .B2(new_n996), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  XOR2_X1   g574(.A(new_n748), .B(new_n751), .Z(new_n1000));
  AOI21_X1  g575(.A(new_n999), .B1(new_n1000), .B2(new_n992), .ZN(new_n1001));
  OR2_X1    g576(.A1(G290), .A2(G1986), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n1002), .B(KEYINPUT109), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n1003), .A2(new_n990), .A3(new_n988), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n1004), .A2(KEYINPUT48), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(KEYINPUT48), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1001), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n995), .A2(KEYINPUT127), .A3(KEYINPUT46), .ZN(new_n1008));
  NAND2_X1  g583(.A1(KEYINPUT127), .A2(KEYINPUT46), .ZN(new_n1009));
  NOR2_X1   g584(.A1(KEYINPUT127), .A2(KEYINPUT46), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1009), .B1(new_n996), .B2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n997), .A2(new_n994), .A3(new_n1008), .A4(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n1012), .B(KEYINPUT47), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n749), .A2(new_n751), .ZN(new_n1014));
  OAI22_X1  g589(.A1(new_n999), .A2(new_n1014), .B1(G2067), .B2(new_n777), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n992), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n1007), .A2(new_n1013), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n985), .A2(KEYINPUT50), .ZN(new_n1018));
  XOR2_X1   g593(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n1019));
  OAI211_X1 g594(.A(new_n978), .B(new_n1019), .C1(new_n983), .C2(new_n984), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1018), .A2(new_n834), .A3(new_n990), .A4(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT115), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1020), .A2(new_n990), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT115), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1023), .A2(new_n1024), .A3(new_n834), .A4(new_n1018), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n506), .A2(KEYINPUT45), .A3(new_n978), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n987), .A2(new_n990), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G1966), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1022), .A2(new_n1025), .A3(new_n1029), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n1030), .A2(new_n598), .A3(G8), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n506), .A2(G160), .A3(G40), .A4(new_n978), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n600), .A2(new_n603), .A3(G1976), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1032), .A2(new_n1033), .A3(G8), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT112), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n1034), .A2(new_n1035), .A3(KEYINPUT52), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1035), .B1(new_n1034), .B2(KEYINPUT52), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT49), .ZN(new_n1039));
  INV_X1    g614(.A(G1981), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n610), .A2(new_n1040), .A3(new_n611), .ZN(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT113), .B(G86), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n528), .A2(new_n530), .A3(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1040), .B1(new_n610), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1039), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1043), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n605), .B1(new_n1047), .B2(new_n614), .ZN(new_n1048));
  OAI21_X1  g623(.A(G1981), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n610), .A2(new_n1040), .A3(new_n611), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(KEYINPUT49), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G125), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(new_n480), .B2(new_n481), .ZN(new_n1053));
  INV_X1    g628(.A(new_n470), .ZN(new_n1054));
  OAI21_X1  g629(.A(G2105), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1055), .A2(G40), .A3(new_n476), .A4(new_n477), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n985), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G8), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1045), .A2(new_n1051), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(G1976), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT52), .B1(G288), .B2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1059), .A2(new_n1033), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1038), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1020), .A2(new_n990), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT50), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1067), .B1(new_n506), .B2(new_n978), .ZN(new_n1068));
  OR3_X1    g643(.A1(new_n1066), .A2(new_n1068), .A3(G2090), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1027), .A2(new_n721), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1058), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1071), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1074), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1056), .B1(new_n985), .B2(new_n986), .ZN(new_n1077));
  AOI21_X1  g652(.A(G1971), .B1(new_n1077), .B2(new_n1026), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1067), .B(new_n978), .C1(new_n983), .C2(new_n984), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n990), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1019), .B1(new_n506), .B2(new_n978), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1080), .A2(new_n1081), .A3(G2090), .ZN(new_n1082));
  OAI21_X1  g657(.A(G8), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1076), .A2(new_n1083), .A3(new_n1072), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1031), .A2(new_n1065), .A3(new_n1075), .A4(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT63), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT116), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1085), .A2(KEYINPUT116), .A3(new_n1086), .ZN(new_n1090));
  NOR3_X1   g665(.A1(new_n1071), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1091), .A2(new_n1086), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1092), .A2(new_n1075), .A3(new_n1065), .A4(new_n1031), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1089), .A2(new_n1090), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1075), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1060), .A2(new_n1061), .A3(new_n731), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n1041), .B(KEYINPUT114), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1095), .A2(new_n1065), .B1(new_n1059), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT62), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT124), .B1(G168), .B2(new_n1058), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT124), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n596), .A2(new_n1102), .A3(G8), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(new_n1030), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1030), .A2(G8), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n596), .A2(new_n1102), .A3(G8), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1102), .B1(new_n596), .B2(G8), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT51), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1106), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1110), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT125), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  AOI211_X1 g689(.A(KEYINPUT125), .B(new_n1110), .C1(new_n1106), .C2(new_n1109), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1100), .B(new_n1105), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1065), .A2(new_n1075), .A3(new_n1084), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1027), .ZN(new_n1118));
  INV_X1    g693(.A(G2078), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1118), .A2(KEYINPUT53), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT118), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1121), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1122));
  INV_X1    g697(.A(G1961), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1018), .A2(KEYINPUT118), .A3(new_n990), .A4(new_n1020), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1122), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT53), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1126), .B1(new_n1027), .B2(G2078), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1120), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(G171), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1117), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1116), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1104), .B1(G8), .B2(new_n1030), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT125), .B1(new_n1132), .B2(new_n1110), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1133), .A2(new_n1134), .A3(new_n1111), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1100), .B1(new_n1135), .B2(new_n1105), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1094), .B(new_n1099), .C1(new_n1131), .C2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1105), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1120), .A2(new_n1125), .A3(G301), .A4(new_n1127), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1129), .A2(KEYINPUT54), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(KEYINPUT54), .B1(new_n1129), .B2(new_n1139), .ZN(new_n1141));
  NOR3_X1   g716(.A1(new_n1140), .A2(new_n1141), .A3(new_n1117), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1138), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT126), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1138), .A2(new_n1142), .A3(KEYINPUT126), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g722(.A(KEYINPUT56), .B(G2072), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1077), .A2(new_n1026), .A3(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n768), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT57), .ZN(new_n1152));
  NAND2_X1  g727(.A1(G299), .A2(new_n1152), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n587), .A2(new_n583), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1154), .A2(KEYINPUT57), .A3(new_n581), .A4(new_n576), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1151), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT117), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n1032), .A2(new_n1159), .A3(G2067), .ZN(new_n1160));
  INV_X1    g735(.A(G2067), .ZN(new_n1161));
  AOI21_X1  g736(.A(KEYINPUT117), .B1(new_n1057), .B2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1122), .A2(new_n787), .A3(new_n1124), .ZN(new_n1164));
  AND2_X1   g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1158), .B1(new_n1165), .B2(new_n631), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1150), .A2(new_n1149), .A3(new_n1156), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1165), .A2(KEYINPUT60), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1163), .A2(new_n1164), .A3(KEYINPUT60), .ZN(new_n1170));
  AOI21_X1  g745(.A(KEYINPUT122), .B1(new_n1170), .B2(new_n630), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1170), .A2(new_n630), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1170), .A2(KEYINPUT122), .A3(new_n630), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1169), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n1176));
  AND3_X1   g751(.A1(new_n1150), .A2(new_n1149), .A3(new_n1156), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1156), .B1(new_n1150), .B2(new_n1149), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1176), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(KEYINPUT120), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT120), .ZN(new_n1181));
  OAI211_X1 g756(.A(new_n1181), .B(new_n1176), .C1(new_n1177), .C2(new_n1178), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1158), .A2(KEYINPUT61), .A3(new_n1167), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT121), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1158), .A2(KEYINPUT121), .A3(KEYINPUT61), .A4(new_n1167), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  OR2_X1    g763(.A1(new_n1027), .A2(G1996), .ZN(new_n1189));
  XOR2_X1   g764(.A(KEYINPUT58), .B(G1341), .Z(new_n1190));
  NAND2_X1  g765(.A1(new_n1032), .A2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n568), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g767(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n1192), .B(new_n1193), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1183), .A2(new_n1188), .A3(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1168), .B1(new_n1175), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1196), .A2(KEYINPUT123), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT123), .ZN(new_n1198));
  OAI211_X1 g773(.A(new_n1198), .B(new_n1168), .C1(new_n1175), .C2(new_n1195), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1137), .B1(new_n1147), .B2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1003), .B1(G1986), .B2(G290), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1001), .B1(new_n991), .B2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1017), .B1(new_n1201), .B2(new_n1203), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g779(.A1(G401), .A2(G229), .A3(new_n464), .A4(G227), .ZN(new_n1206));
  NAND4_X1  g780(.A1(new_n967), .A2(new_n911), .A3(new_n971), .A4(new_n1206), .ZN(G225));
  INV_X1    g781(.A(G225), .ZN(G308));
endmodule


