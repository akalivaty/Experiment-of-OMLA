//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 1 1 1 1 1 1 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:08 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n555, new_n557, new_n558, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n827, new_n828, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1171, new_n1172,
    new_n1173, new_n1174;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT67), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  XNOR2_X1  g030(.A(G325), .B(KEYINPUT68), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  XNOR2_X1  g033(.A(KEYINPUT3), .B(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G125), .ZN(new_n460));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n458), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT3), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT70), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT70), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n469), .A3(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n465), .A2(new_n470), .A3(G137), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n463), .A2(new_n464), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n462), .B1(new_n474), .B2(new_n458), .ZN(G160));
  NAND2_X1  g050(.A1(new_n465), .A2(new_n470), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(new_n458), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n476), .A2(new_n458), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n458), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  NAND3_X1  g061(.A1(new_n465), .A2(new_n470), .A3(G126), .ZN(new_n487));
  NAND2_X1  g062(.A1(G114), .A2(G2104), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n458), .A2(G102), .A3(G2104), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n490), .A2(KEYINPUT71), .A3(new_n491), .ZN(new_n492));
  AND2_X1   g067(.A1(KEYINPUT4), .A2(G138), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n465), .A2(new_n470), .A3(new_n458), .A4(new_n493), .ZN(new_n494));
  AND2_X1   g069(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n495));
  NOR2_X1   g070(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n496));
  OAI211_X1 g071(.A(G138), .B(new_n458), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT71), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n458), .B1(new_n487), .B2(new_n488), .ZN(new_n502));
  INV_X1    g077(.A(new_n491), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n492), .A2(new_n500), .A3(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT72), .B1(new_n507), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT5), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n508), .A2(new_n511), .B1(new_n507), .B2(G543), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OR2_X1    g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  XOR2_X1   g094(.A(KEYINPUT73), .B(G88), .Z(new_n520));
  NAND2_X1  g095(.A1(new_n512), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(G50), .A2(G543), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n519), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n515), .A2(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  NAND3_X1  g100(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n526));
  XOR2_X1   g101(.A(new_n526), .B(KEYINPUT74), .Z(new_n527));
  INV_X1    g102(.A(KEYINPUT75), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n518), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n516), .A2(KEYINPUT75), .A3(new_n517), .ZN(new_n530));
  AND3_X1   g105(.A1(new_n529), .A2(G543), .A3(new_n530), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n512), .A2(new_n518), .ZN(new_n532));
  AOI22_X1  g107(.A1(G51), .A2(new_n531), .B1(new_n532), .B2(G89), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n527), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XOR2_X1   g110(.A(new_n535), .B(KEYINPUT7), .Z(new_n536));
  NOR2_X1   g111(.A1(new_n534), .A2(new_n536), .ZN(G168));
  NAND3_X1  g112(.A1(new_n529), .A2(G543), .A3(new_n530), .ZN(new_n538));
  INV_X1    g113(.A(G52), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n512), .A2(new_n518), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n538), .A2(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n514), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n542), .A2(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  AOI22_X1  g121(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT76), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G651), .ZN(new_n549));
  AOI22_X1  g124(.A1(G43), .A2(new_n531), .B1(new_n532), .B2(G81), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(G860), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT77), .ZN(G153));
  AND3_X1   g129(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G36), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n555), .A2(new_n558), .ZN(G188));
  NAND2_X1  g134(.A1(new_n531), .A2(G53), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT9), .ZN(new_n561));
  XOR2_X1   g136(.A(KEYINPUT79), .B(G65), .Z(new_n562));
  NAND2_X1  g137(.A1(new_n512), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n514), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT78), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n540), .B(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G91), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n568), .A2(new_n571), .ZN(G299));
  INV_X1    g147(.A(G168), .ZN(G286));
  NAND4_X1  g148(.A1(new_n529), .A2(G49), .A3(G543), .A4(new_n530), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT80), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n574), .B(new_n575), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n540), .B(KEYINPUT78), .ZN(new_n578));
  INV_X1    g153(.A(G87), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n576), .B(new_n577), .C1(new_n578), .C2(new_n579), .ZN(G288));
  NAND3_X1  g155(.A1(new_n518), .A2(G48), .A3(G543), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n582), .B2(new_n514), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(G86), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n578), .B2(new_n585), .ZN(G305));
  AOI22_X1  g161(.A1(G47), .A2(new_n531), .B1(new_n532), .B2(G85), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n514), .B2(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n570), .A2(G92), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n591), .B(new_n592), .ZN(new_n593));
  AND2_X1   g168(.A1(new_n512), .A2(G66), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT81), .ZN(new_n596));
  OAI21_X1  g171(.A(G651), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n531), .A2(G54), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n593), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n590), .B1(new_n600), .B2(G868), .ZN(G284));
  OAI21_X1  g176(.A(new_n590), .B1(new_n600), .B2(G868), .ZN(G321));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  NOR2_X1   g178(.A1(G168), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT82), .ZN(new_n605));
  INV_X1    g180(.A(new_n571), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n567), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n605), .B1(G868), .B2(new_n607), .ZN(G297));
  OAI21_X1  g183(.A(new_n605), .B1(G868), .B2(new_n607), .ZN(G280));
  AOI21_X1  g184(.A(new_n599), .B1(G559), .B2(new_n552), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT83), .ZN(G148));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n600), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G868), .ZN(new_n614));
  INV_X1    g189(.A(new_n551), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(G868), .B2(new_n615), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n481), .A2(G123), .ZN(new_n618));
  INV_X1    g193(.A(G135), .ZN(new_n619));
  NOR2_X1   g194(.A1(G99), .A2(G2105), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(new_n458), .B2(G111), .ZN(new_n621));
  OAI221_X1 g196(.A(new_n618), .B1(new_n478), .B2(new_n619), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(G2096), .Z(new_n623));
  NAND3_X1  g198(.A1(new_n472), .A2(new_n459), .A3(new_n458), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(KEYINPUT13), .B(G2100), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n623), .A2(new_n628), .ZN(G156));
  XNOR2_X1  g204(.A(G2451), .B(G2454), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT16), .ZN(new_n631));
  XOR2_X1   g206(.A(G2443), .B(G2446), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G1341), .B(G1348), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NOR2_X1   g210(.A1(KEYINPUT85), .A2(KEYINPUT14), .ZN(new_n636));
  XOR2_X1   g211(.A(KEYINPUT15), .B(G2435), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2438), .ZN(new_n638));
  XOR2_X1   g213(.A(G2427), .B(G2430), .Z(new_n639));
  AOI21_X1  g214(.A(new_n636), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(new_n638), .B2(new_n639), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n641), .B1(KEYINPUT85), .B2(KEYINPUT14), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n635), .B(new_n642), .Z(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(G14), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(G401));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT86), .ZN(new_n647));
  XOR2_X1   g222(.A(G2067), .B(G2678), .Z(new_n648));
  OR2_X1    g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(new_n650), .A3(KEYINPUT17), .ZN(new_n651));
  INV_X1    g226(.A(KEYINPUT18), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2096), .B(G2100), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2072), .B(G2078), .Z(new_n656));
  AOI21_X1  g231(.A(new_n656), .B1(new_n649), .B2(KEYINPUT18), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n655), .B(new_n657), .ZN(G227));
  XNOR2_X1  g233(.A(G1971), .B(G1976), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  XOR2_X1   g235(.A(G1956), .B(G2474), .Z(new_n661));
  XOR2_X1   g236(.A(G1961), .B(G1966), .Z(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n660), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n661), .A2(new_n662), .ZN(new_n666));
  AOI22_X1  g241(.A1(new_n664), .A2(KEYINPUT20), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n666), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n668), .A2(new_n660), .A3(new_n663), .ZN(new_n669));
  OAI211_X1 g244(.A(new_n667), .B(new_n669), .C1(KEYINPUT20), .C2(new_n664), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT87), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G1991), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G1981), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1986), .B(G1996), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n672), .B(new_n676), .ZN(G229));
  INV_X1    g252(.A(G29), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(G27), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n679), .B1(G164), .B2(new_n678), .ZN(new_n680));
  INV_X1    g255(.A(G2078), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(G16), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G21), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(G168), .B2(new_n683), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1966), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(G5), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(G171), .B2(new_n683), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G1961), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT31), .B(G11), .Z(new_n690));
  OR2_X1    g265(.A1(G29), .A2(G33), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n459), .A2(G127), .ZN(new_n692));
  AND2_X1   g267(.A1(G115), .A2(G2104), .ZN(new_n693));
  OAI21_X1  g268(.A(G2105), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT25), .Z(new_n696));
  INV_X1    g271(.A(G139), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n694), .B(new_n696), .C1(new_n478), .C2(new_n697), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n691), .B1(new_n698), .B2(new_n678), .ZN(new_n699));
  INV_X1    g274(.A(G2072), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n622), .A2(new_n678), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n699), .A2(new_n700), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT97), .B(G28), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT30), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(new_n678), .ZN(new_n706));
  NAND4_X1  g281(.A1(new_n701), .A2(new_n702), .A3(new_n703), .A4(new_n706), .ZN(new_n707));
  NOR3_X1   g282(.A1(new_n689), .A2(new_n690), .A3(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G1348), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n683), .A2(G4), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n599), .B2(G16), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n708), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n709), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT98), .ZN(new_n714));
  INV_X1    g289(.A(G35), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(G29), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n715), .A2(G29), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n485), .B2(G29), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n716), .B1(new_n718), .B2(new_n714), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT99), .B(KEYINPUT29), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n713), .B1(new_n721), .B2(G2090), .ZN(new_n722));
  AND2_X1   g297(.A1(KEYINPUT89), .A2(G16), .ZN(new_n723));
  NOR2_X1   g298(.A1(KEYINPUT89), .A2(G16), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G19), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n615), .B2(new_n726), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n728), .A2(G1341), .ZN(new_n729));
  NOR2_X1   g304(.A1(G29), .A2(G32), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n479), .A2(G141), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n481), .A2(G129), .ZN(new_n732));
  NAND3_X1  g307(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT26), .Z(new_n734));
  NAND3_X1  g309(.A1(new_n472), .A2(G105), .A3(new_n458), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n731), .A2(new_n732), .A3(new_n734), .A4(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n730), .B1(new_n737), .B2(G29), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT27), .B(G1996), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G2084), .ZN(new_n741));
  NAND2_X1  g316(.A1(G160), .A2(G29), .ZN(new_n742));
  AND2_X1   g317(.A1(KEYINPUT24), .A2(G34), .ZN(new_n743));
  NOR2_X1   g318(.A1(KEYINPUT24), .A2(G34), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n678), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(KEYINPUT95), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n745), .A2(KEYINPUT95), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n742), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n728), .A2(G1341), .B1(new_n741), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n748), .A2(new_n741), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT96), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n729), .A2(new_n740), .A3(new_n749), .A4(new_n751), .ZN(new_n752));
  OR4_X1    g327(.A1(new_n686), .A2(new_n712), .A3(new_n722), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n481), .A2(G128), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT93), .ZN(new_n755));
  OR2_X1    g330(.A1(G104), .A2(G2105), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n756), .B(G2104), .C1(G116), .C2(new_n458), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n479), .A2(G140), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n755), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n759), .A2(KEYINPUT94), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(KEYINPUT94), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n762), .A2(new_n678), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n678), .A2(G26), .ZN(new_n764));
  OAI21_X1  g339(.A(KEYINPUT28), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n764), .A2(KEYINPUT28), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(G2067), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n726), .A2(G20), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT101), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT23), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G299), .B2(G16), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G1956), .ZN(new_n773));
  INV_X1    g348(.A(G2067), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n765), .A2(new_n774), .A3(new_n766), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n768), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n721), .A2(G2090), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT100), .ZN(new_n778));
  NOR3_X1   g353(.A1(new_n753), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n683), .A2(G23), .ZN(new_n780));
  INV_X1    g355(.A(G288), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n780), .B1(new_n781), .B2(new_n683), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT92), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT33), .B(G1976), .Z(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n783), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(G305), .A2(G16), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n683), .A2(G6), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n789), .A2(KEYINPUT91), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(KEYINPUT91), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT32), .B(G1981), .Z(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G166), .A2(new_n726), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G22), .B2(new_n726), .ZN(new_n796));
  INV_X1    g371(.A(G1971), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(new_n793), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n790), .A2(new_n791), .A3(new_n799), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n796), .A2(new_n797), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n794), .A2(new_n798), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(KEYINPUT34), .B1(new_n786), .B2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n802), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n783), .B(new_n784), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT34), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(G25), .A2(G29), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n479), .A2(G131), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n481), .A2(G119), .ZN(new_n810));
  OR2_X1    g385(.A1(G95), .A2(G2105), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n811), .B(G2104), .C1(G107), .C2(new_n458), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n809), .A2(new_n810), .A3(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n808), .B1(new_n814), .B2(G29), .ZN(new_n815));
  XNOR2_X1  g390(.A(KEYINPUT35), .B(G1991), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT88), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n815), .B(new_n817), .ZN(new_n818));
  MUX2_X1   g393(.A(G24), .B(G290), .S(new_n725), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT90), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G1986), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n803), .A2(new_n807), .A3(new_n818), .A4(new_n821), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n822), .A2(KEYINPUT36), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n822), .A2(KEYINPUT36), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n682), .B(new_n779), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(G311));
  INV_X1    g401(.A(KEYINPUT102), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n822), .B(KEYINPUT36), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n829), .A2(KEYINPUT102), .A3(new_n682), .A4(new_n779), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n830), .ZN(G150));
  INV_X1    g406(.A(G55), .ZN(new_n832));
  INV_X1    g407(.A(G93), .ZN(new_n833));
  OAI22_X1  g408(.A1(new_n538), .A2(new_n832), .B1(new_n540), .B2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT103), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n835), .B1(new_n514), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(G860), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT37), .Z(new_n839));
  NOR2_X1   g414(.A1(new_n599), .A2(new_n612), .ZN(new_n840));
  XNOR2_X1  g415(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT104), .ZN(new_n843));
  AND2_X1   g418(.A1(new_n837), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n615), .B1(new_n837), .B2(new_n843), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n845), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n842), .B(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n839), .B1(new_n849), .B2(G860), .ZN(G145));
  INV_X1    g425(.A(G142), .ZN(new_n851));
  NOR2_X1   g426(.A1(G106), .A2(G2105), .ZN(new_n852));
  OAI21_X1  g427(.A(G2104), .B1(new_n458), .B2(G118), .ZN(new_n853));
  OAI22_X1  g428(.A1(new_n478), .A2(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(G130), .B2(new_n481), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n814), .B(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n626), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n760), .A2(new_n761), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n490), .A2(new_n500), .A3(new_n491), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n698), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n861), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n760), .A2(new_n761), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n862), .A2(new_n737), .A3(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n737), .B1(new_n862), .B2(new_n864), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n858), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n867), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n869), .A2(new_n857), .A3(new_n865), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n868), .A2(new_n870), .A3(KEYINPUT106), .ZN(new_n871));
  XNOR2_X1  g446(.A(G160), .B(KEYINPUT105), .ZN(new_n872));
  XNOR2_X1  g447(.A(G162), .B(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n622), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT106), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n875), .B(new_n858), .C1(new_n866), .C2(new_n867), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n871), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(G37), .ZN(new_n878));
  INV_X1    g453(.A(new_n874), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n868), .A2(new_n870), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n877), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(KEYINPUT107), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT107), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n877), .A2(new_n883), .A3(new_n878), .A4(new_n880), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n882), .A2(KEYINPUT40), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(KEYINPUT40), .B1(new_n882), .B2(new_n884), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(G395));
  XNOR2_X1  g462(.A(new_n599), .B(new_n607), .ZN(new_n888));
  XNOR2_X1  g463(.A(KEYINPUT108), .B(KEYINPUT41), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n599), .B(G299), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n892), .A2(KEYINPUT41), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n848), .B(new_n613), .ZN(new_n895));
  MUX2_X1   g470(.A(new_n894), .B(new_n892), .S(new_n895), .Z(new_n896));
  XOR2_X1   g471(.A(G290), .B(KEYINPUT109), .Z(new_n897));
  AOI21_X1  g472(.A(new_n583), .B1(new_n570), .B2(G86), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(G303), .ZN(new_n899));
  OR2_X1    g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n897), .A2(new_n899), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(G288), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n902), .A2(G288), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(KEYINPUT42), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n896), .B(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(G868), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n837), .A2(new_n603), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(G295));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n910), .ZN(G331));
  XNOR2_X1  g487(.A(G168), .B(G171), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n846), .A2(new_n847), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n913), .B1(new_n846), .B2(new_n847), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n914), .B(new_n916), .C1(new_n891), .C2(new_n893), .ZN(new_n917));
  INV_X1    g492(.A(new_n914), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n888), .B1(new_n918), .B2(new_n915), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n917), .A2(new_n906), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n878), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT110), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n922), .B1(new_n904), .B2(new_n905), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n900), .A2(new_n901), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(new_n781), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n925), .A2(KEYINPUT110), .A3(new_n903), .ZN(new_n926));
  AOI22_X1  g501(.A1(new_n917), .A2(new_n919), .B1(new_n923), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(KEYINPUT43), .B1(new_n921), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n923), .A2(new_n926), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT41), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n892), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n888), .A2(new_n889), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n916), .A2(new_n931), .A3(new_n932), .A4(new_n914), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n919), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n929), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n935), .A2(new_n936), .A3(new_n878), .A4(new_n920), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n928), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n936), .B1(new_n921), .B2(new_n927), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n935), .A2(new_n878), .A3(new_n920), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n939), .B1(new_n936), .B2(new_n940), .ZN(new_n941));
  MUX2_X1   g516(.A(new_n938), .B(new_n941), .S(KEYINPUT44), .Z(G397));
  INV_X1    g517(.A(KEYINPUT113), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n943), .B1(G160), .B2(G40), .ZN(new_n944));
  AOI21_X1  g519(.A(G2105), .B1(new_n471), .B2(new_n473), .ZN(new_n945));
  INV_X1    g520(.A(G40), .ZN(new_n946));
  NOR4_X1   g521(.A1(new_n945), .A2(new_n462), .A3(KEYINPUT113), .A4(new_n946), .ZN(new_n947));
  OR2_X1    g522(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  XOR2_X1   g523(.A(KEYINPUT111), .B(G1384), .Z(new_n949));
  NAND2_X1  g524(.A1(new_n860), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n948), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G1996), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  XOR2_X1   g531(.A(new_n956), .B(KEYINPUT46), .Z(new_n957));
  XNOR2_X1  g532(.A(new_n859), .B(new_n774), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n737), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n957), .B1(new_n959), .B2(new_n954), .ZN(new_n960));
  XOR2_X1   g535(.A(new_n960), .B(KEYINPUT47), .Z(new_n961));
  INV_X1    g536(.A(new_n954), .ZN(new_n962));
  NOR3_X1   g537(.A1(new_n962), .A2(G1986), .A3(G290), .ZN(new_n963));
  XOR2_X1   g538(.A(new_n963), .B(KEYINPUT48), .Z(new_n964));
  XNOR2_X1  g539(.A(new_n736), .B(new_n955), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n958), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n813), .A2(new_n816), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n813), .A2(new_n816), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n964), .B1(new_n969), .B2(new_n962), .ZN(new_n970));
  INV_X1    g545(.A(new_n967), .ZN(new_n971));
  OAI22_X1  g546(.A1(new_n966), .A2(new_n971), .B1(G2067), .B2(new_n859), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n954), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n961), .A2(new_n970), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT114), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n494), .A2(new_n499), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n502), .A2(new_n978), .A3(new_n503), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n977), .B1(new_n979), .B2(G1384), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT45), .ZN(new_n981));
  INV_X1    g556(.A(G1384), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n860), .A2(KEYINPUT114), .A3(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n980), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n944), .A2(new_n947), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n505), .A2(new_n982), .A3(new_n951), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G1966), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT119), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT50), .B1(new_n980), .B2(new_n983), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT50), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n993), .B1(new_n505), .B2(new_n982), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n992), .A2(new_n994), .A3(new_n948), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n741), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n987), .A2(KEYINPUT119), .A3(new_n988), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n991), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n976), .B1(new_n998), .B2(G286), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n991), .A2(new_n996), .A3(G168), .A4(new_n997), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(G8), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n976), .B1(new_n1000), .B2(G8), .ZN(new_n1003));
  OAI21_X1  g578(.A(KEYINPUT62), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n860), .A2(KEYINPUT45), .A3(new_n949), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n985), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n951), .B1(new_n505), .B2(new_n982), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT53), .B1(new_n1008), .B2(new_n681), .ZN(new_n1009));
  INV_X1    g584(.A(G1961), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n980), .A2(new_n983), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n993), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n505), .A2(new_n982), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT50), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1012), .A2(new_n1014), .A3(new_n985), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1009), .B1(new_n1010), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n681), .A2(KEYINPUT53), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1016), .B1(new_n987), .B2(new_n1017), .ZN(new_n1018));
  AND2_X1   g593(.A1(new_n1018), .A2(G171), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1001), .A2(KEYINPUT51), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT62), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1020), .B(new_n1021), .C1(new_n1001), .C2(new_n999), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n781), .A2(G1976), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n979), .A2(new_n977), .A3(G1384), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT114), .B1(new_n860), .B2(new_n982), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n985), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n1023), .A2(new_n1026), .A3(G8), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT116), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1023), .A2(G8), .A3(new_n1026), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1030), .A2(new_n1031), .A3(KEYINPUT52), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT117), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n781), .A2(G1976), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1027), .A2(new_n1034), .A3(new_n1028), .A4(new_n1036), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1023), .A2(new_n1026), .A3(new_n1028), .A4(G8), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT117), .B1(new_n1038), .B2(new_n1035), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  OAI22_X1  g615(.A1(new_n1015), .A2(G2090), .B1(G1971), .B2(new_n1008), .ZN(new_n1041));
  NAND2_X1  g616(.A1(G303), .A2(G8), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT55), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n1044));
  NAND3_X1  g619(.A1(G303), .A2(new_n1044), .A3(G8), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1046), .B(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1041), .A2(new_n1048), .A3(G8), .ZN(new_n1049));
  INV_X1    g624(.A(G1981), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n898), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n583), .B1(G86), .B2(new_n532), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1051), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n1053), .B(KEYINPUT49), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1026), .A2(G8), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1033), .A2(new_n1040), .A3(new_n1049), .A4(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n980), .A2(KEYINPUT50), .A3(new_n983), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n985), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT118), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1013), .A2(KEYINPUT50), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1058), .A2(new_n1063), .A3(new_n985), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1060), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  OAI22_X1  g640(.A1(new_n1065), .A2(G2090), .B1(G1971), .B2(new_n1008), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1066), .A2(G8), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1057), .A2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1004), .A2(new_n1019), .A3(new_n1022), .A4(new_n1068), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1033), .A2(new_n1040), .A3(new_n1056), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n998), .A2(G8), .A3(G168), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT63), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1041), .A2(G8), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1073), .B1(new_n1074), .B2(new_n1046), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1070), .A2(new_n1049), .A3(new_n1072), .A4(new_n1075), .ZN(new_n1076));
  NOR3_X1   g651(.A1(new_n1057), .A2(new_n1067), .A3(new_n1071), .ZN(new_n1077));
  XOR2_X1   g652(.A(KEYINPUT120), .B(KEYINPUT63), .Z(new_n1078));
  OAI21_X1  g653(.A(new_n1076), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1049), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1070), .A2(new_n1080), .ZN(new_n1081));
  AOI211_X1 g656(.A(G1976), .B(G288), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1051), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1055), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1069), .A2(new_n1079), .A3(new_n1081), .A4(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(G1956), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1065), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT121), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n607), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1091));
  NAND2_X1  g666(.A1(KEYINPUT121), .A2(KEYINPUT57), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1091), .B(new_n1092), .C1(new_n567), .C2(new_n606), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT56), .B(G2072), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1008), .A2(new_n1095), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1087), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1026), .A2(G2067), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1098), .B1(new_n1015), .B2(new_n709), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT122), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n1099), .A2(new_n1100), .A3(new_n599), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1011), .A2(new_n774), .A3(new_n985), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(new_n995), .B2(G1348), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT122), .B1(new_n1103), .B2(new_n600), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1064), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1063), .B1(new_n1058), .B2(new_n985), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n1106), .A2(new_n1107), .A3(new_n1061), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1096), .B1(new_n1108), .B2(G1956), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1094), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1097), .B1(new_n1105), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT124), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT123), .B(KEYINPUT58), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n1114), .B(G1341), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  AOI211_X1 g691(.A(new_n1113), .B(new_n1116), .C1(new_n1011), .C2(new_n985), .ZN(new_n1117));
  AOI21_X1  g692(.A(KEYINPUT124), .B1(new_n1026), .B2(new_n1115), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1007), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1120), .A2(new_n955), .A3(new_n985), .A4(new_n1005), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT125), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1026), .A2(new_n1115), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n1113), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1026), .A2(KEYINPUT124), .A3(new_n1115), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1124), .A2(KEYINPUT125), .A3(new_n1121), .A4(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n615), .B1(new_n1122), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT59), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1124), .A2(new_n1121), .A3(new_n1125), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT125), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(new_n1126), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT59), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1133), .A2(new_n1134), .A3(new_n615), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1129), .A2(new_n1135), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1094), .B(new_n1096), .C1(new_n1108), .C2(G1956), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT61), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1087), .A2(KEYINPUT61), .A3(new_n1094), .A4(new_n1096), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT60), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n600), .B1(new_n1103), .B2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1099), .A2(KEYINPUT60), .A3(new_n599), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1103), .A2(new_n1141), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1139), .A2(new_n1140), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  AOI211_X1 g721(.A(KEYINPUT126), .B(new_n1112), .C1(new_n1136), .C2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT126), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1134), .B1(new_n1133), .B2(new_n615), .ZN(new_n1151));
  AOI211_X1 g726(.A(KEYINPUT59), .B(new_n551), .C1(new_n1132), .C2(new_n1126), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1149), .B(new_n1150), .C1(new_n1151), .C2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1112), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1148), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1147), .A2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1020), .B1(new_n1001), .B2(new_n999), .ZN(new_n1157));
  XOR2_X1   g732(.A(G301), .B(KEYINPUT54), .Z(new_n1158));
  AND3_X1   g733(.A1(new_n953), .A2(G40), .A3(G160), .ZN(new_n1159));
  XOR2_X1   g734(.A(KEYINPUT127), .B(G2078), .Z(new_n1160));
  NAND4_X1  g735(.A1(new_n1159), .A2(KEYINPUT53), .A3(new_n1005), .A4(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1016), .A2(new_n1158), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1158), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1018), .A2(new_n1163), .ZN(new_n1164));
  AND4_X1   g739(.A1(new_n1157), .A2(new_n1068), .A3(new_n1162), .A4(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1085), .B1(new_n1156), .B2(new_n1165), .ZN(new_n1166));
  XOR2_X1   g741(.A(G290), .B(G1986), .Z(new_n1167));
  AOI21_X1  g742(.A(new_n962), .B1(new_n969), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n975), .B1(new_n1166), .B2(new_n1168), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g744(.A1(new_n882), .A2(new_n884), .ZN(new_n1171));
  INV_X1    g745(.A(G319), .ZN(new_n1172));
  OR3_X1    g746(.A1(G229), .A2(new_n1172), .A3(G227), .ZN(new_n1173));
  AOI21_X1  g747(.A(new_n1173), .B1(new_n928), .B2(new_n937), .ZN(new_n1174));
  NAND3_X1  g748(.A1(new_n1171), .A2(new_n1174), .A3(new_n644), .ZN(G225));
  INV_X1    g749(.A(G225), .ZN(G308));
endmodule


