//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 1 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 0 0 1 1 0 0 0 0 0 1 1 0 1 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1271, new_n1272, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1334, new_n1335,
    new_n1336, new_n1337;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n210), .B1(new_n203), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  INV_X1    g0017(.A(G107), .ZN(new_n218));
  INV_X1    g0018(.A(G264), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n209), .B1(new_n214), .B2(new_n220), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n206), .A2(G50), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n209), .A2(G13), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n229), .B(G250), .C1(G257), .C2(G264), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT0), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n222), .A2(new_n228), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT65), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n237), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(G50), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n203), .A2(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n245), .B(new_n251), .Z(G351));
  OAI21_X1  g0052(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n253));
  INV_X1    g0053(.A(G150), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n226), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT8), .B(G58), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT67), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n202), .A2(KEYINPUT67), .A3(KEYINPUT8), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n255), .A2(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  OAI221_X1 g0063(.A(new_n253), .B1(new_n254), .B2(new_n256), .C1(new_n261), .C2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n225), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G1), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(G13), .A3(G20), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(G50), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n266), .B1(new_n268), .B2(G20), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n270), .B1(new_n271), .B2(G50), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT3), .B(G33), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G222), .A2(G1698), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(G223), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n275), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G41), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n280), .A2(G1), .A3(G13), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n279), .B(new_n282), .C1(G77), .C2(new_n275), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT66), .ZN(new_n284));
  INV_X1    g0084(.A(G41), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G45), .ZN(new_n287));
  NAND2_X1  g0087(.A1(KEYINPUT66), .A2(G41), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G274), .ZN(new_n290));
  AND2_X1   g0090(.A1(G1), .A2(G13), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n290), .B1(new_n291), .B2(new_n280), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n289), .A2(new_n292), .A3(new_n268), .ZN(new_n293));
  INV_X1    g0093(.A(G226), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n268), .B1(G41), .B2(G45), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n281), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n283), .B(new_n293), .C1(new_n294), .C2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G169), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n300), .B1(G179), .B2(new_n298), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n274), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G190), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n304), .B1(G200), .B2(new_n298), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT9), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n274), .A2(new_n306), .ZN(new_n307));
  NOR3_X1   g0107(.A1(new_n267), .A2(KEYINPUT9), .A3(new_n273), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n305), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT10), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT10), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n311), .B(new_n305), .C1(new_n307), .C2(new_n308), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n302), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n271), .A2(G77), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n314), .B1(G77), .B2(new_n269), .ZN(new_n315));
  NAND2_X1  g0115(.A1(G20), .A2(G77), .ZN(new_n316));
  AND2_X1   g0116(.A1(new_n212), .A2(KEYINPUT15), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n212), .A2(KEYINPUT15), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT68), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  XNOR2_X1  g0119(.A(KEYINPUT15), .B(G87), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT68), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  OAI221_X1 g0123(.A(new_n316), .B1(new_n256), .B2(new_n257), .C1(new_n323), .C2(new_n263), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n315), .B1(new_n324), .B2(new_n266), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n275), .A2(G232), .A3(new_n277), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n275), .A2(G238), .A3(G1698), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n327), .B(new_n328), .C1(new_n218), .C2(new_n275), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n282), .ZN(new_n330));
  INV_X1    g0130(.A(G179), .ZN(new_n331));
  AND2_X1   g0131(.A1(KEYINPUT66), .A2(G41), .ZN(new_n332));
  NOR2_X1   g0132(.A1(KEYINPUT66), .A2(G41), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(G1), .B1(new_n334), .B2(new_n287), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n335), .A2(new_n292), .B1(new_n296), .B2(G244), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n330), .A2(new_n331), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n330), .A2(new_n336), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n299), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n326), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(G200), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n341), .B(new_n325), .C1(new_n303), .C2(new_n338), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g0143(.A(new_n343), .B(KEYINPUT69), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT13), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n294), .A2(G1698), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT3), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G33), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n346), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT70), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n275), .A2(KEYINPUT70), .A3(new_n346), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n348), .A2(new_n349), .A3(G232), .A4(G1698), .ZN(new_n355));
  NAND2_X1  g0155(.A1(G33), .A2(G97), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n281), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n293), .B1(new_n297), .B2(new_n211), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n345), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n335), .A2(new_n292), .B1(new_n296), .B2(G238), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n355), .A2(new_n356), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n362), .B1(new_n352), .B2(new_n353), .ZN(new_n363));
  OAI211_X1 g0163(.A(KEYINPUT13), .B(new_n361), .C1(new_n363), .C2(new_n281), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT14), .B1(new_n365), .B2(new_n299), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT71), .ZN(new_n367));
  OAI22_X1  g0167(.A1(new_n358), .A2(new_n359), .B1(new_n367), .B2(new_n345), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(new_n367), .B2(new_n364), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G179), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT14), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n360), .A2(new_n371), .A3(new_n364), .A4(G169), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n372), .A2(KEYINPUT72), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n372), .A2(KEYINPUT72), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n366), .B(new_n370), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n263), .A2(new_n216), .ZN(new_n376));
  OAI22_X1  g0176(.A1(new_n256), .A2(new_n246), .B1(new_n226), .B2(G68), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n266), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT11), .ZN(new_n379));
  AND2_X1   g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n378), .A2(new_n379), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n271), .A2(G68), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT12), .ZN(new_n383));
  INV_X1    g0183(.A(new_n269), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n383), .B1(new_n384), .B2(new_n203), .ZN(new_n385));
  NOR3_X1   g0185(.A1(new_n269), .A2(KEYINPUT12), .A3(G68), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n382), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NOR3_X1   g0187(.A1(new_n380), .A2(new_n381), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n375), .A2(new_n389), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n369), .A2(G190), .ZN(new_n391));
  INV_X1    g0191(.A(G200), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n388), .B1(new_n365), .B2(new_n392), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n313), .A2(new_n344), .A3(new_n390), .A4(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT16), .ZN(new_n397));
  INV_X1    g0197(.A(G159), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n256), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(G58), .A2(G68), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n204), .A2(new_n205), .A3(new_n400), .ZN(new_n401));
  AOI211_X1 g0201(.A(new_n397), .B(new_n399), .C1(new_n401), .C2(G20), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT7), .ZN(new_n403));
  AND3_X1   g0203(.A1(new_n347), .A2(KEYINPUT73), .A3(G33), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT73), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n404), .B1(new_n275), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n403), .B1(new_n406), .B2(new_n226), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n348), .A2(new_n349), .A3(new_n405), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n347), .A2(KEYINPUT73), .A3(G33), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n408), .A2(new_n403), .A3(new_n226), .A4(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(G68), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n402), .B1(new_n407), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n403), .B1(new_n275), .B2(G20), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n348), .A2(new_n349), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n414), .A2(KEYINPUT7), .A3(new_n226), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n203), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n401), .A2(G20), .ZN(new_n417));
  INV_X1    g0217(.A(new_n399), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n397), .B1(new_n416), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n412), .A2(new_n420), .A3(new_n266), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n261), .A2(new_n271), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n422), .B1(new_n261), .B2(new_n269), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT74), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n281), .A2(G232), .A3(new_n295), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n293), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n426), .B1(new_n293), .B2(new_n427), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OR2_X1    g0231(.A1(G223), .A2(G1698), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n294), .A2(G1698), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  OAI22_X1  g0234(.A1(new_n406), .A2(new_n434), .B1(new_n255), .B2(new_n212), .ZN(new_n435));
  AOI21_X1  g0235(.A(G190), .B1(new_n435), .B2(new_n282), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n434), .B1(new_n408), .B2(new_n409), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n255), .A2(new_n212), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n282), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n335), .A2(new_n292), .B1(new_n296), .B2(G232), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n431), .A2(new_n436), .B1(new_n441), .B2(new_n392), .ZN(new_n442));
  OAI21_X1  g0242(.A(KEYINPUT76), .B1(new_n425), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n441), .A2(new_n392), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n293), .A2(new_n427), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT74), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n446), .A2(new_n303), .A3(new_n428), .A4(new_n439), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT76), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n448), .A2(new_n449), .A3(new_n421), .A4(new_n424), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n443), .A2(KEYINPUT17), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT17), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n448), .A2(new_n452), .A3(new_n421), .A4(new_n424), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT77), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n443), .A2(KEYINPUT77), .A3(KEYINPUT17), .A4(new_n450), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT18), .ZN(new_n458));
  AOI21_X1  g0258(.A(G179), .B1(new_n435), .B2(new_n282), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n431), .A2(new_n459), .B1(new_n441), .B2(new_n299), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n425), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n458), .B1(new_n425), .B2(new_n460), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n461), .A2(new_n462), .A3(KEYINPUT75), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT75), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n265), .A2(new_n225), .ZN(new_n465));
  AOI21_X1  g0265(.A(KEYINPUT7), .B1(new_n414), .B2(new_n226), .ZN(new_n466));
  AOI211_X1 g0266(.A(new_n403), .B(G20), .C1(new_n348), .C2(new_n349), .ZN(new_n467));
  OAI21_X1  g0267(.A(G68), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n399), .B1(new_n401), .B2(G20), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n465), .B1(new_n470), .B2(new_n397), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n423), .B1(new_n471), .B2(new_n412), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n441), .A2(new_n299), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n446), .A2(new_n331), .A3(new_n428), .A4(new_n439), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(KEYINPUT18), .B1(new_n472), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n425), .A2(new_n458), .A3(new_n460), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n464), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n456), .B(new_n457), .C1(new_n463), .C2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n396), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G283), .ZN(new_n481));
  INV_X1    g0281(.A(G97), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n481), .B(new_n226), .C1(G33), .C2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G116), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G20), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n483), .A2(new_n266), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT20), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n483), .A2(KEYINPUT20), .A3(new_n266), .A4(new_n485), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n269), .A2(G116), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n255), .A2(G1), .ZN(new_n492));
  NOR3_X1   g0292(.A1(new_n384), .A2(new_n266), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n491), .B1(new_n493), .B2(G116), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n299), .B1(new_n490), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT5), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n268), .B(G45), .C1(new_n496), .C2(G41), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n496), .B1(new_n332), .B2(new_n333), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n282), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(KEYINPUT5), .B1(new_n286), .B2(new_n288), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(new_n497), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n500), .A2(G270), .B1(new_n502), .B2(new_n292), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n219), .A2(G1698), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n504), .B1(G257), .B2(G1698), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n505), .B1(new_n409), .B2(new_n408), .ZN(new_n506));
  INV_X1    g0306(.A(G303), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n275), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n282), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n495), .A2(new_n510), .A3(KEYINPUT21), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT82), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT82), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n495), .A2(new_n510), .A3(new_n513), .A4(KEYINPUT21), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(KEYINPUT21), .B1(new_n495), .B2(new_n510), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n503), .A2(G179), .A3(new_n509), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n490), .A2(new_n494), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n510), .A2(G200), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n521), .B(new_n518), .C1(new_n303), .C2(new_n510), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n515), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(KEYINPUT83), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT83), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n515), .A2(new_n520), .A3(new_n525), .A4(new_n522), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(KEYINPUT84), .B1(new_n226), .B2(G107), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT23), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT23), .ZN(new_n530));
  OAI211_X1 g0330(.A(KEYINPUT84), .B(new_n530), .C1(new_n226), .C2(G107), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n212), .A2(G20), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n533), .A2(new_n348), .A3(new_n349), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT22), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n262), .A2(G116), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n532), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(KEYINPUT22), .A2(G87), .ZN(new_n539));
  AOI211_X1 g0339(.A(G20), .B(new_n539), .C1(new_n408), .C2(new_n409), .ZN(new_n540));
  OAI21_X1  g0340(.A(KEYINPUT24), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n408), .A2(new_n409), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n542), .A2(KEYINPUT22), .A3(new_n226), .A4(G87), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT24), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n534), .A2(new_n535), .B1(G116), .B2(new_n262), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n543), .A2(new_n544), .A3(new_n532), .A4(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n266), .ZN(new_n548));
  XOR2_X1   g0348(.A(KEYINPUT85), .B(KEYINPUT25), .Z(new_n549));
  NOR2_X1   g0349(.A1(new_n269), .A2(G107), .ZN(new_n550));
  XNOR2_X1  g0350(.A(new_n549), .B(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n493), .A2(G107), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n548), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT86), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n498), .A2(new_n499), .A3(new_n292), .ZN(new_n557));
  OAI211_X1 g0357(.A(G264), .B(new_n281), .C1(new_n501), .C2(new_n497), .ZN(new_n558));
  INV_X1    g0358(.A(G294), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n255), .A2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(G257), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(G1698), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(G250), .B2(G1698), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n560), .B1(new_n542), .B2(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n557), .B(new_n558), .C1(new_n565), .C2(new_n281), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n299), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n563), .B1(new_n409), .B2(new_n408), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n282), .B1(new_n568), .B2(new_n560), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n569), .A2(new_n331), .A3(new_n557), .A4(new_n558), .ZN(new_n570));
  AND2_X1   g0370(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n555), .A2(new_n556), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n553), .B1(new_n547), .B2(new_n266), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n569), .A2(G190), .A3(new_n557), .A4(new_n558), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n566), .A2(G200), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n567), .A2(new_n570), .ZN(new_n577));
  OAI21_X1  g0377(.A(KEYINPUT86), .B1(new_n573), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n572), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n211), .A2(new_n277), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n217), .A2(G1698), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n582), .B1(new_n408), .B2(new_n409), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n255), .A2(new_n484), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n282), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT79), .ZN(new_n586));
  OAI22_X1  g0386(.A1(new_n586), .A2(new_n213), .B1(new_n287), .B2(G1), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n268), .A2(new_n290), .A3(G45), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n213), .A2(KEYINPUT79), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n587), .B(new_n281), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n585), .A2(G179), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n299), .B1(new_n585), .B2(new_n590), .ZN(new_n592));
  OAI21_X1  g0392(.A(KEYINPUT80), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n585), .A2(new_n590), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G169), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT80), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n585), .A2(G179), .A3(new_n590), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT81), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n465), .B(new_n269), .C1(G1), .C2(new_n255), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n599), .B1(new_n323), .B2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n493), .A2(KEYINPUT81), .A3(new_n322), .A4(new_n319), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n323), .A2(new_n384), .ZN(new_n604));
  AOI211_X1 g0404(.A(G20), .B(new_n203), .C1(new_n408), .C2(new_n409), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT19), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n263), .B2(new_n482), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n226), .B1(new_n356), .B2(new_n606), .ZN(new_n608));
  NOR2_X1   g0408(.A1(G97), .A2(G107), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n212), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n266), .B1(new_n605), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n603), .A2(new_n604), .A3(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n593), .A2(new_n598), .A3(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n594), .A2(new_n303), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n392), .B1(new_n585), .B2(new_n590), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n493), .A2(G87), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n613), .A2(new_n619), .A3(new_n604), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(G107), .B1(new_n466), .B2(new_n467), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n256), .A2(new_n216), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT6), .ZN(new_n625));
  AND2_X1   g0425(.A1(G97), .A2(G107), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n625), .B1(new_n626), .B2(new_n609), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT78), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n628), .A2(new_n218), .A3(KEYINPUT6), .A4(G97), .ZN(new_n629));
  NAND2_X1  g0429(.A1(KEYINPUT6), .A2(G97), .ZN(new_n630));
  OAI21_X1  g0430(.A(KEYINPUT78), .B1(new_n630), .B2(G107), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n627), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n624), .B1(new_n632), .B2(G20), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n465), .B1(new_n623), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n384), .A2(new_n482), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n600), .B2(new_n482), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(G250), .A2(G1698), .ZN(new_n638));
  NAND2_X1  g0438(.A1(KEYINPUT4), .A2(G244), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n638), .B1(new_n639), .B2(G1698), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n275), .A2(new_n640), .B1(G33), .B2(G283), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n277), .A2(G244), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n642), .B1(new_n408), .B2(new_n409), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n641), .B1(new_n643), .B2(KEYINPUT4), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n282), .ZN(new_n645));
  OAI211_X1 g0445(.A(G257), .B(new_n281), .C1(new_n501), .C2(new_n497), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n557), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n299), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n647), .B1(new_n282), .B2(new_n644), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n331), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n637), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n649), .A2(G200), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n634), .A2(new_n636), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n651), .A2(G190), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n615), .A2(new_n622), .A3(new_n653), .A4(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n579), .A2(new_n658), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n480), .A2(new_n527), .A3(new_n659), .ZN(G372));
  NOR2_X1   g0460(.A1(new_n461), .A2(new_n462), .ZN(new_n661));
  INV_X1    g0461(.A(new_n390), .ZN(new_n662));
  INV_X1    g0462(.A(new_n340), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n662), .B1(new_n395), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n456), .A2(new_n457), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n661), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n310), .A2(new_n312), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n302), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n480), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n515), .A2(new_n520), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n555), .A2(new_n571), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n603), .A2(new_n604), .A3(new_n613), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT87), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n674), .B1(new_n591), .B2(new_n592), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n595), .A2(KEYINPUT87), .A3(new_n597), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n673), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n616), .A2(new_n620), .A3(new_n617), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AND3_X1   g0479(.A1(new_n576), .A2(new_n653), .A3(new_n657), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n672), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  OAI22_X1  g0482(.A1(new_n651), .A2(G169), .B1(new_n634), .B2(new_n636), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n645), .A2(new_n331), .A3(new_n648), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n615), .A2(new_n685), .A3(new_n622), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(KEYINPUT26), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n591), .A2(new_n592), .A3(new_n674), .ZN(new_n689));
  AOI21_X1  g0489(.A(KEYINPUT87), .B1(new_n595), .B2(new_n597), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n614), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT26), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n691), .A2(new_n692), .A3(new_n685), .A4(new_n622), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n691), .ZN(new_n694));
  OAI21_X1  g0494(.A(KEYINPUT88), .B1(new_n688), .B2(new_n694), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n677), .A2(new_n653), .A3(new_n678), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n677), .B1(new_n696), .B2(new_n692), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT88), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(new_n698), .A3(new_n687), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n682), .B1(new_n695), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n668), .B1(new_n669), .B2(new_n700), .ZN(G369));
  NAND3_X1  g0501(.A1(new_n268), .A2(new_n226), .A3(G13), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n702), .A2(KEYINPUT27), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(KEYINPUT27), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(G213), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT89), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(G343), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(new_n518), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT90), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(new_n670), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n713), .B1(new_n527), .B2(new_n712), .ZN(new_n714));
  INV_X1    g0514(.A(G330), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n579), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(new_n573), .B2(new_n710), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n671), .B2(new_n710), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n670), .A2(new_n709), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(new_n717), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n710), .A2(new_n555), .A3(new_n571), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT91), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n721), .A2(new_n726), .ZN(G399));
  INV_X1    g0527(.A(new_n334), .ZN(new_n728));
  INV_X1    g0528(.A(new_n229), .ZN(new_n729));
  OAI21_X1  g0529(.A(KEYINPUT92), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n728), .A2(KEYINPUT92), .A3(new_n729), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n609), .A2(new_n212), .A3(new_n484), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n733), .A2(new_n268), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n735), .B1(new_n224), .B2(new_n733), .ZN(new_n736));
  XOR2_X1   g0536(.A(new_n736), .B(KEYINPUT28), .Z(new_n737));
  NAND4_X1  g0537(.A1(new_n572), .A2(new_n578), .A3(new_n515), .A4(new_n520), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n738), .A2(new_n680), .A3(new_n679), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n686), .A2(new_n692), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n691), .A2(KEYINPUT26), .A3(new_n685), .A4(new_n622), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n739), .A2(new_n742), .A3(new_n691), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n743), .A2(new_n710), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT29), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n700), .A2(new_n709), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n746), .B1(new_n747), .B2(new_n745), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT93), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT30), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n585), .A2(new_n590), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n651), .A2(new_n751), .A3(new_n558), .A4(new_n569), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n750), .B1(new_n752), .B2(new_n517), .ZN(new_n753));
  AOI21_X1  g0553(.A(G179), .B1(new_n503), .B2(new_n509), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n649), .A2(new_n754), .A3(new_n566), .A4(new_n594), .ZN(new_n755));
  INV_X1    g0555(.A(new_n517), .ZN(new_n756));
  AND4_X1   g0556(.A1(new_n558), .A2(new_n569), .A3(new_n585), .A4(new_n590), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n756), .A2(new_n757), .A3(KEYINPUT30), .A4(new_n651), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n753), .A2(new_n755), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n709), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT31), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n749), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(KEYINPUT31), .B1(new_n759), .B2(new_n709), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n527), .A2(new_n659), .A3(new_n710), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n715), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AND2_X1   g0567(.A1(new_n748), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n737), .B1(new_n768), .B2(G1), .ZN(G364));
  NOR2_X1   g0569(.A1(G13), .A2(G33), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n714), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n225), .B1(G20), .B2(new_n299), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n226), .A2(new_n331), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n775), .A2(G190), .A3(G200), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n226), .A2(G190), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n331), .A2(G200), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n777), .A2(G326), .B1(new_n781), .B2(G311), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G179), .A2(G200), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT96), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n778), .B1(new_n784), .B2(G20), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AND2_X1   g0586(.A1(new_n786), .A2(KEYINPUT98), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(KEYINPUT98), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n782), .B1(new_n789), .B2(new_n559), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(KEYINPUT99), .Z(new_n791));
  NAND3_X1  g0591(.A1(new_n775), .A2(new_n303), .A3(G200), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G317), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(KEYINPUT33), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n794), .A2(KEYINPUT33), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n793), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n392), .A2(G179), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n778), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n275), .B1(new_n800), .B2(G283), .ZN(new_n801));
  INV_X1    g0601(.A(G322), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n226), .A2(new_n303), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(new_n779), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n797), .B(new_n801), .C1(new_n802), .C2(new_n804), .ZN(new_n805));
  NOR3_X1   g0605(.A1(new_n784), .A2(new_n226), .A3(G190), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(G329), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n803), .A2(new_n798), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n808), .A2(KEYINPUT97), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(KEYINPUT97), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n807), .B1(new_n811), .B2(new_n507), .ZN(new_n812));
  NOR3_X1   g0612(.A1(new_n791), .A2(new_n805), .A3(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n789), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(G97), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n806), .A2(G159), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT32), .Z(new_n817));
  OAI22_X1  g0617(.A1(new_n804), .A2(new_n202), .B1(new_n780), .B2(new_n216), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT95), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n792), .A2(new_n203), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n275), .B1(new_n799), .B2(new_n218), .C1(new_n776), .C2(new_n246), .ZN(new_n821));
  INV_X1    g0621(.A(new_n811), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n820), .B(new_n821), .C1(new_n822), .C2(G87), .ZN(new_n823));
  AND4_X1   g0623(.A1(new_n815), .A2(new_n817), .A3(new_n819), .A4(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n774), .B1(new_n813), .B2(new_n824), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n226), .A2(G13), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n268), .B1(new_n826), .B2(G45), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n733), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n729), .A2(new_n414), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n831), .A2(G355), .B1(new_n484), .B2(new_n729), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n251), .A2(new_n287), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n542), .A2(new_n729), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(G45), .B2(new_n223), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n832), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n772), .A2(new_n774), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT94), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n830), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n773), .A2(new_n825), .A3(new_n840), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(KEYINPUT100), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n830), .B1(new_n714), .B2(new_n715), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(new_n715), .B2(new_n714), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(G396));
  AOI21_X1  g0646(.A(new_n698), .B1(new_n697), .B2(new_n687), .ZN(new_n847));
  AND4_X1   g0647(.A1(new_n698), .A2(new_n687), .A3(new_n691), .A4(new_n693), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n681), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n343), .A2(new_n709), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n342), .B1(new_n710), .B2(new_n325), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n340), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n663), .A2(new_n710), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n851), .B1(new_n747), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n767), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n766), .B(new_n851), .C1(new_n747), .C2(new_n856), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n858), .A2(new_n830), .A3(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT101), .ZN(new_n861));
  INV_X1    g0661(.A(new_n774), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n771), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n829), .B1(G77), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(G283), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n792), .A2(new_n865), .B1(new_n776), .B2(new_n507), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n804), .A2(new_n559), .B1(new_n799), .B2(new_n212), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n414), .B1(new_n780), .B2(new_n484), .ZN(new_n868));
  NOR3_X1   g0668(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n822), .A2(G107), .B1(G311), .B2(new_n806), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n815), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n804), .ZN(new_n872));
  AOI22_X1  g0672(.A1(G143), .A2(new_n872), .B1(new_n781), .B2(G159), .ZN(new_n873));
  INV_X1    g0673(.A(G137), .ZN(new_n874));
  OAI221_X1 g0674(.A(new_n873), .B1(new_n874), .B2(new_n776), .C1(new_n254), .C2(new_n792), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT34), .ZN(new_n876));
  OR2_X1    g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n875), .A2(new_n876), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n822), .A2(G50), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n799), .A2(new_n203), .ZN(new_n880));
  AOI211_X1 g0680(.A(new_n406), .B(new_n880), .C1(new_n806), .C2(G132), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n877), .A2(new_n878), .A3(new_n879), .A4(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n789), .A2(new_n202), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n871), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n864), .B1(new_n884), .B2(new_n774), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n856), .B2(new_n771), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n860), .A2(new_n861), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n861), .B1(new_n860), .B2(new_n886), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(G384));
  OR2_X1    g0690(.A1(new_n632), .A2(KEYINPUT35), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n632), .A2(KEYINPUT35), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n891), .A2(G116), .A3(new_n227), .A4(new_n892), .ZN(new_n893));
  XOR2_X1   g0693(.A(new_n893), .B(KEYINPUT36), .Z(new_n894));
  NAND3_X1  g0694(.A1(new_n224), .A2(G77), .A3(new_n400), .ZN(new_n895));
  AOI211_X1 g0695(.A(new_n268), .B(G13), .C1(new_n895), .C2(new_n247), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n850), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n854), .B1(new_n700), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n709), .A2(new_n389), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n390), .A2(new_n395), .A3(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n389), .B(new_n709), .C1(new_n375), .C2(new_n394), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n412), .A2(new_n266), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n408), .A2(new_n226), .A3(new_n409), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT7), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n907), .A2(G68), .A3(new_n410), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT16), .B1(new_n908), .B2(new_n469), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n424), .B1(new_n905), .B2(new_n909), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n910), .A2(new_n706), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n479), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT37), .B1(new_n425), .B2(new_n460), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n425), .A2(new_n706), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n443), .A2(new_n913), .A3(new_n450), .A4(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n475), .A2(new_n707), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n910), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n443), .A2(new_n917), .A3(new_n450), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT102), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n918), .A2(new_n919), .A3(KEYINPUT37), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n919), .B1(new_n918), .B2(KEYINPUT37), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n915), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT38), .B1(new_n912), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n912), .A2(new_n922), .A3(KEYINPUT38), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT103), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n912), .A2(new_n922), .A3(KEYINPUT103), .A4(KEYINPUT38), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n923), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n904), .A2(new_n928), .B1(new_n661), .B2(new_n706), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(KEYINPUT104), .ZN(new_n930));
  XOR2_X1   g0730(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n456), .A2(new_n661), .A3(new_n457), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n933), .A2(new_n425), .A3(new_n706), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n425), .A2(new_n460), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n935), .B(new_n914), .C1(new_n425), .C2(new_n442), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(KEYINPUT37), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n915), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n932), .B1(new_n934), .B2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT39), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n940), .A2(new_n941), .A3(new_n924), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n928), .B2(new_n941), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n662), .A2(new_n710), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT104), .ZN(new_n947));
  OAI221_X1 g0747(.A(new_n947), .B1(new_n661), .B2(new_n706), .C1(new_n904), .C2(new_n928), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n930), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n748), .A2(new_n669), .ZN(new_n950));
  INV_X1    g0750(.A(new_n668), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n949), .B(new_n952), .Z(new_n953));
  INV_X1    g0753(.A(new_n923), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT38), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n918), .A2(KEYINPUT37), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(KEYINPUT102), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n918), .A2(new_n919), .A3(KEYINPUT37), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n955), .B1(new_n959), .B2(new_n915), .ZN(new_n960));
  AOI21_X1  g0760(.A(KEYINPUT103), .B1(new_n960), .B2(new_n912), .ZN(new_n961));
  INV_X1    g0761(.A(new_n927), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n954), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n855), .B1(new_n901), .B2(new_n902), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n760), .A2(new_n761), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n965), .A2(new_n763), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n765), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT40), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AND3_X1   g0770(.A1(new_n912), .A2(new_n922), .A3(KEYINPUT38), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n968), .B1(new_n971), .B2(new_n939), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n963), .A2(new_n970), .B1(new_n972), .B2(KEYINPUT40), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n480), .A2(new_n967), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n715), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n975), .B2(new_n974), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n953), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n268), .B2(new_n826), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n953), .A2(new_n977), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n897), .B1(new_n979), .B2(new_n980), .ZN(G367));
  OAI211_X1 g0781(.A(new_n653), .B(new_n657), .C1(new_n710), .C2(new_n655), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n685), .A2(new_n709), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT107), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(new_n578), .B2(new_n572), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n710), .B1(new_n986), .B2(new_n685), .ZN(new_n987));
  INV_X1    g0787(.A(new_n984), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n723), .A2(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT42), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n710), .A2(new_n621), .ZN(new_n992));
  MUX2_X1   g0792(.A(new_n679), .B(new_n677), .S(new_n992), .Z(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT43), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n991), .B(new_n996), .C1(new_n997), .C2(new_n994), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n991), .B2(new_n996), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n720), .A2(new_n985), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n726), .A2(new_n988), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT44), .Z(new_n1003));
  NOR2_X1   g0803(.A1(new_n726), .A2(new_n988), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT45), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n721), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n723), .B1(new_n719), .B2(new_n722), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n716), .B(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1003), .A2(new_n720), .A3(new_n1005), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1007), .A2(new_n768), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n768), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n733), .B(KEYINPUT41), .ZN(new_n1013));
  AND2_X1   g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1001), .B1(new_n1014), .B2(new_n828), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n789), .A2(new_n218), .B1(new_n865), .B2(new_n780), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT109), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n811), .A2(new_n484), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT46), .Z(new_n1019));
  AOI22_X1  g0819(.A1(new_n793), .A2(G294), .B1(new_n777), .B2(G311), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(G303), .A2(new_n872), .B1(new_n800), .B2(G97), .ZN(new_n1021));
  AND3_X1   g0821(.A1(new_n1020), .A2(new_n406), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n806), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1019), .B(new_n1022), .C1(new_n794), .C2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n789), .A2(new_n203), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n822), .A2(G58), .B1(G137), .B2(new_n806), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n275), .B1(new_n799), .B2(new_n216), .C1(new_n254), .C2(new_n804), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(G143), .B2(new_n777), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n792), .A2(new_n398), .B1(new_n780), .B2(new_n246), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT110), .Z(new_n1030));
  NAND3_X1  g0830(.A1(new_n1026), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n1017), .A2(new_n1024), .B1(new_n1025), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT47), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n862), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n1033), .B2(new_n1032), .ZN(new_n1035));
  AND2_X1   g0835(.A1(new_n241), .A2(new_n834), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n839), .B1(new_n229), .B2(new_n323), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n829), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT108), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n772), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1035), .B(new_n1039), .C1(new_n1040), .C2(new_n993), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1015), .A2(new_n1041), .ZN(G387));
  NAND2_X1  g0842(.A1(new_n1009), .A2(new_n828), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n719), .A2(new_n1040), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n831), .A2(new_n734), .B1(new_n218), .B2(new_n729), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n237), .A2(new_n287), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n257), .A2(G50), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT50), .ZN(new_n1048));
  AOI211_X1 g0848(.A(G45), .B(new_n734), .C1(G68), .C2(G77), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(new_n834), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1045), .B1(new_n1046), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n830), .B1(new_n1052), .B2(new_n839), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n789), .A2(new_n323), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n261), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n822), .A2(G77), .B1(new_n1055), .B2(new_n793), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n254), .B2(new_n1023), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G50), .A2(new_n872), .B1(new_n800), .B2(G97), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n203), .B2(new_n780), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n542), .B1(new_n398), .B2(new_n776), .ZN(new_n1060));
  NOR4_X1   g0860(.A1(new_n1054), .A2(new_n1057), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(G317), .A2(new_n872), .B1(new_n781), .B2(G303), .ZN(new_n1062));
  INV_X1    g0862(.A(G311), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1062), .B1(new_n1063), .B2(new_n792), .C1(new_n802), .C2(new_n776), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT48), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n1064), .A2(new_n1065), .B1(new_n559), .B2(new_n811), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(G283), .B2(new_n814), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT111), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n1065), .B2(new_n1064), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1069), .A2(KEYINPUT49), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n806), .A2(G326), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1071), .B(new_n406), .C1(new_n484), .C2(new_n799), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n1069), .B2(KEYINPUT49), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1061), .B1(new_n1070), .B2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1053), .B1(new_n1074), .B2(new_n862), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n768), .A2(new_n1009), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n733), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n768), .A2(new_n1009), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1043), .B1(new_n1044), .B2(new_n1075), .C1(new_n1077), .C2(new_n1078), .ZN(G393));
  NAND2_X1  g0879(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n1076), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1081), .A2(new_n1011), .A3(new_n733), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT115), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1082), .B(new_n1083), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1080), .A2(new_n827), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n985), .A2(new_n772), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n793), .A2(G303), .B1(new_n781), .B2(G294), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n789), .B2(new_n484), .ZN(new_n1088));
  XOR2_X1   g0888(.A(new_n1088), .B(KEYINPUT113), .Z(new_n1089));
  OAI22_X1  g0889(.A1(new_n776), .A2(new_n794), .B1(new_n804), .B2(new_n1063), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT52), .Z(new_n1091));
  AOI21_X1  g0891(.A(new_n275), .B1(new_n800), .B2(G107), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1092), .B1(new_n1023), .B2(new_n802), .C1(new_n811), .C2(new_n865), .ZN(new_n1093));
  NOR3_X1   g0893(.A1(new_n1089), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n814), .A2(G77), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n257), .A2(new_n780), .B1(new_n799), .B2(new_n212), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n406), .B(new_n1096), .C1(G50), .C2(new_n793), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n822), .A2(G68), .B1(G143), .B2(new_n806), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n776), .A2(new_n254), .B1(new_n804), .B2(new_n398), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT51), .ZN(new_n1100));
  AND4_X1   g0900(.A1(new_n1095), .A2(new_n1097), .A3(new_n1098), .A4(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n774), .B1(new_n1094), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n245), .A2(new_n834), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n839), .B(new_n1103), .C1(new_n482), .C2(new_n229), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT112), .Z(new_n1105));
  NAND3_X1  g0905(.A1(new_n1102), .A2(new_n829), .A3(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT114), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1085), .B1(new_n1086), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1084), .A2(new_n1108), .ZN(G390));
  OAI21_X1  g0909(.A(new_n829), .B1(new_n1055), .B2(new_n863), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n811), .A2(new_n254), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT53), .ZN(new_n1112));
  INV_X1    g0912(.A(G125), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1023), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(G132), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n275), .B1(new_n804), .B2(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(KEYINPUT54), .B(G143), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n1117), .A2(new_n780), .B1(new_n799), .B2(new_n246), .ZN(new_n1118));
  INV_X1    g0918(.A(G128), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n792), .A2(new_n874), .B1(new_n776), .B2(new_n1119), .ZN(new_n1120));
  NOR4_X1   g0920(.A1(new_n1114), .A2(new_n1116), .A3(new_n1118), .A4(new_n1120), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1112), .B(new_n1121), .C1(new_n398), .C2(new_n789), .ZN(new_n1122));
  OR2_X1    g0922(.A1(new_n1122), .A2(KEYINPUT118), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n792), .A2(new_n218), .B1(new_n776), .B2(new_n865), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n804), .A2(new_n484), .B1(new_n780), .B2(new_n482), .ZN(new_n1125));
  NOR4_X1   g0925(.A1(new_n1124), .A2(new_n1125), .A3(new_n275), .A4(new_n880), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n822), .A2(G87), .B1(G294), .B2(new_n806), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1095), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1122), .A2(KEYINPUT118), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1123), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1110), .B1(new_n1130), .B2(new_n774), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n943), .B2(new_n771), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT119), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1132), .B(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n854), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(new_n849), .B2(new_n850), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n903), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n944), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1138), .B(new_n942), .C1(new_n941), .C2(new_n928), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n940), .A2(new_n924), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n743), .A2(new_n710), .A3(new_n853), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n854), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT116), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1141), .A2(KEYINPUT116), .A3(new_n854), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n944), .B(new_n1140), .C1(new_n1146), .C2(new_n1137), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n766), .A2(new_n856), .A3(new_n903), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1139), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n944), .B1(new_n971), .B2(new_n939), .ZN(new_n1150));
  AND3_X1   g0950(.A1(new_n1141), .A2(KEYINPUT116), .A3(new_n854), .ZN(new_n1151));
  AOI21_X1  g0951(.A(KEYINPUT116), .B1(new_n1141), .B2(new_n854), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1150), .B1(new_n1153), .B2(new_n903), .ZN(new_n1154));
  NOR3_X1   g0954(.A1(new_n971), .A2(new_n939), .A3(KEYINPUT39), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(new_n963), .B2(KEYINPUT39), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1154), .B1(new_n1156), .B2(new_n1138), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n967), .A2(G330), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n964), .ZN(new_n1160));
  OAI211_X1 g0960(.A(KEYINPUT117), .B(new_n1149), .C1(new_n1157), .C2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1139), .A2(new_n1147), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT117), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1160), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1161), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1134), .B1(new_n1166), .B2(new_n828), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n903), .B1(new_n766), .B2(new_n856), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n899), .B1(new_n1168), .B2(new_n1164), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1137), .B1(new_n1158), .B2(new_n855), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1148), .A2(new_n1146), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1159), .A2(new_n480), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n668), .B(new_n1173), .C1(new_n748), .C2(new_n669), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1172), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1161), .A2(new_n1165), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n733), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1176), .B1(new_n1161), .B2(new_n1165), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1167), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(KEYINPUT120), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT120), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1167), .B(new_n1182), .C1(new_n1178), .C2(new_n1179), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(G378));
  OAI21_X1  g0985(.A(new_n706), .B1(new_n267), .B2(new_n273), .ZN(new_n1186));
  OR2_X1    g0986(.A1(new_n313), .A2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n313), .B1(new_n274), .B2(new_n707), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1189), .B(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n973), .B2(new_n715), .ZN(new_n1192));
  XOR2_X1   g0992(.A(new_n1189), .B(new_n1190), .Z(new_n1193));
  NAND2_X1  g0993(.A1(new_n968), .A2(new_n969), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n928), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n969), .B1(new_n1140), .B2(new_n968), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1193), .B(G330), .C1(new_n1195), .C2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1192), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n949), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n929), .A2(KEYINPUT104), .B1(new_n943), .B2(new_n945), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1200), .A2(new_n1192), .A3(new_n1197), .A4(new_n948), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1191), .A2(new_n770), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n829), .B1(G50), .B2(new_n863), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n542), .A2(new_n728), .ZN(new_n1205));
  AOI211_X1 g1005(.A(G50), .B(new_n1205), .C1(new_n255), .C2(new_n285), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(G107), .A2(new_n872), .B1(new_n800), .B2(G58), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1207), .B1(new_n482), .B2(new_n792), .C1(new_n484), .C2(new_n776), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1205), .B1(new_n811), .B2(new_n216), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n1023), .A2(new_n865), .B1(new_n323), .B2(new_n780), .ZN(new_n1210));
  OR4_X1    g1010(.A1(new_n1025), .A2(new_n1208), .A3(new_n1209), .A4(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT58), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1206), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n811), .A2(new_n1117), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(G128), .A2(new_n872), .B1(new_n781), .B2(G137), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n1215), .B1(new_n1113), .B2(new_n776), .C1(new_n1115), .C2(new_n792), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1214), .B(new_n1216), .C1(new_n814), .C2(G150), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1218), .A2(KEYINPUT59), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n255), .B(new_n285), .C1(new_n799), .C2(new_n398), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n806), .B2(G124), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT59), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1221), .B1(new_n1217), .B2(new_n1222), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1213), .B1(new_n1212), .B2(new_n1211), .C1(new_n1219), .C2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1204), .B1(new_n1224), .B2(new_n774), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n1202), .A2(new_n828), .B1(new_n1203), .B2(new_n1225), .ZN(new_n1226));
  AOI211_X1 g1026(.A(KEYINPUT117), .B(new_n1160), .C1(new_n1139), .C2(new_n1147), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1163), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1227), .B1(new_n1228), .B2(new_n1149), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1175), .B1(new_n1229), .B2(new_n1176), .ZN(new_n1230));
  AOI21_X1  g1030(.A(KEYINPUT57), .B1(new_n1230), .B2(new_n1202), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1174), .B1(new_n1166), .B2(new_n1172), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1198), .A2(new_n949), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n948), .A2(new_n1200), .B1(new_n1192), .B2(new_n1197), .ZN(new_n1234));
  OAI21_X1  g1034(.A(KEYINPUT57), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n733), .B1(new_n1232), .B2(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1226), .B1(new_n1231), .B2(new_n1236), .ZN(G375));
  NAND3_X1  g1037(.A1(new_n1169), .A2(new_n1174), .A3(new_n1171), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1176), .A2(new_n1013), .A3(new_n1238), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1239), .B(KEYINPUT121), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1172), .A2(new_n828), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n829), .B1(G68), .B2(new_n863), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(G58), .A2(new_n800), .B1(new_n781), .B2(G150), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n542), .B(new_n1243), .C1(new_n1023), .C2(new_n1119), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(G159), .B2(new_n822), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1245), .B1(new_n246), .B2(new_n789), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1246), .B(KEYINPUT122), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n872), .A2(G137), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n1248), .B1(new_n1115), .B2(new_n776), .C1(new_n792), .C2(new_n1117), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n792), .A2(new_n484), .B1(new_n776), .B2(new_n559), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n804), .A2(new_n865), .B1(new_n780), .B2(new_n218), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n414), .B1(new_n799), .B2(new_n216), .ZN(new_n1252));
  NOR3_X1   g1052(.A1(new_n1250), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n1253), .B1(new_n507), .B2(new_n1023), .C1(new_n482), .C2(new_n811), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n1247), .A2(new_n1249), .B1(new_n1054), .B2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1242), .B1(new_n1255), .B2(new_n774), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1256), .B1(new_n903), .B2(new_n771), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1241), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1240), .A2(new_n1259), .ZN(G381));
  OR3_X1    g1060(.A1(G384), .A2(G393), .A3(G396), .ZN(new_n1261));
  NOR4_X1   g1061(.A1(G390), .A2(G387), .A3(G381), .A4(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1180), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n733), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT57), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(new_n1199), .B2(new_n1201), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1264), .B1(new_n1230), .B2(new_n1266), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1230), .A2(new_n1202), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1267), .B1(new_n1268), .B2(KEYINPUT57), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1262), .A2(new_n1263), .A3(new_n1269), .A4(new_n1226), .ZN(G407));
  NAND2_X1  g1070(.A1(new_n708), .A2(G213), .ZN(new_n1271));
  OR3_X1    g1071(.A1(G375), .A2(new_n1180), .A3(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(G407), .A2(G213), .A3(new_n1272), .ZN(G409));
  NAND4_X1  g1073(.A1(new_n1169), .A2(new_n1174), .A3(KEYINPUT60), .A4(new_n1171), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n733), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1176), .A2(KEYINPUT60), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1275), .B1(new_n1276), .B2(new_n1238), .ZN(new_n1277));
  OAI21_X1  g1077(.A(G384), .B1(new_n1277), .B2(new_n1258), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1174), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT60), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1238), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1281), .A2(new_n733), .A3(new_n1274), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1282), .A2(new_n889), .A3(new_n1259), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1278), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT124), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n708), .A2(G213), .A3(G2897), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1278), .A2(KEYINPUT124), .A3(new_n1283), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1286), .A2(new_n1287), .A3(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(KEYINPUT125), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT125), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1286), .A2(new_n1291), .A3(new_n1287), .A4(new_n1288), .ZN(new_n1292));
  OR2_X1    g1092(.A1(new_n1284), .A2(new_n1287), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1290), .A2(new_n1292), .A3(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT123), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1202), .A2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1199), .A2(KEYINPUT123), .A3(new_n1201), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1297), .A2(new_n828), .A3(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1203), .A2(new_n1225), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n1013), .B(new_n1202), .C1(new_n1179), .C2(new_n1174), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1299), .A2(new_n1300), .A3(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1263), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1303), .B1(new_n1184), .B2(G375), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1271), .ZN(new_n1305));
  AOI21_X1  g1105(.A(KEYINPUT61), .B1(new_n1295), .B2(new_n1305), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(G393), .B(new_n845), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1084), .A2(new_n1108), .A3(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1308), .B1(new_n1084), .B2(new_n1108), .ZN(new_n1310));
  NOR3_X1   g1110(.A1(new_n1309), .A2(new_n1310), .A3(G387), .ZN(new_n1311));
  INV_X1    g1111(.A(G387), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(G390), .A2(new_n1307), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1084), .A2(new_n1108), .A3(new_n1308), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1312), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1311), .A2(new_n1315), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1269), .A2(new_n1181), .A3(new_n1183), .A4(new_n1226), .ZN(new_n1317));
  AOI22_X1  g1117(.A1(new_n1317), .A2(new_n1303), .B1(G213), .B2(new_n708), .ZN(new_n1318));
  AND2_X1   g1118(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1318), .A2(KEYINPUT63), .A3(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1304), .A2(new_n1271), .A3(new_n1319), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT63), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1306), .A2(new_n1316), .A3(new_n1320), .A4(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT61), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1325), .B1(new_n1318), .B2(new_n1294), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT127), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1304), .A2(KEYINPUT62), .A3(new_n1271), .A4(new_n1319), .ZN(new_n1328));
  XOR2_X1   g1128(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1329));
  AOI22_X1  g1129(.A1(new_n1327), .A2(new_n1328), .B1(new_n1321), .B2(new_n1329), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1318), .A2(KEYINPUT127), .A3(KEYINPUT62), .A4(new_n1319), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1326), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1324), .B1(new_n1332), .B2(new_n1316), .ZN(G405));
  NAND2_X1  g1133(.A1(G375), .A2(new_n1263), .ZN(new_n1334));
  AND3_X1   g1134(.A1(new_n1317), .A2(new_n1284), .A3(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1319), .B1(new_n1317), .B2(new_n1334), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  XOR2_X1   g1137(.A(new_n1316), .B(new_n1337), .Z(G402));
endmodule


