//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 1 1 1 1 1 1 0 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1279,
    new_n1280, new_n1281, new_n1282, new_n1283, new_n1284, new_n1285,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(new_n207));
  INV_X1    g0007(.A(G13), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  OR2_X1    g0013(.A1(new_n213), .A2(KEYINPUT65), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(KEYINPUT65), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  AND4_X1   g0019(.A1(new_n216), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n220), .A2(new_n207), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT1), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(new_n201), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n225), .A2(G50), .A3(new_n226), .ZN(new_n227));
  NAND4_X1  g0027(.A1(new_n214), .A2(new_n215), .A3(new_n222), .A4(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT66), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G97), .B(G107), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G87), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n202), .A2(G68), .ZN(new_n241));
  INV_X1    g0041(.A(G68), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n240), .B(new_n246), .Z(G351));
  AND2_X1   g0047(.A1(G33), .A2(G41), .ZN(new_n248));
  OAI21_X1  g0048(.A(KEYINPUT67), .B1(new_n248), .B2(new_n223), .ZN(new_n249));
  INV_X1    g0049(.A(G1), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n250), .B1(G41), .B2(G45), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT67), .ZN(new_n254));
  NAND4_X1  g0054(.A1(new_n253), .A2(new_n254), .A3(G1), .A4(G13), .ZN(new_n255));
  NAND4_X1  g0055(.A1(new_n249), .A2(new_n252), .A3(G274), .A4(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  AND2_X1   g0057(.A1(new_n249), .A2(new_n255), .ZN(new_n258));
  AND2_X1   g0058(.A1(new_n258), .A2(new_n251), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n257), .B1(new_n259), .B2(G226), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n248), .A2(new_n223), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT3), .B(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G1698), .ZN(new_n264));
  INV_X1    g0064(.A(G223), .ZN(new_n265));
  INV_X1    g0065(.A(G77), .ZN(new_n266));
  OAI22_X1  g0066(.A1(new_n264), .A2(new_n265), .B1(new_n266), .B2(new_n263), .ZN(new_n267));
  OR2_X1    g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  AOI21_X1  g0069(.A(G1698), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n267), .B1(G222), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n260), .B1(new_n262), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G190), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n274), .B1(G200), .B2(new_n272), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n203), .A2(G20), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G20), .A2(G33), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n277), .A2(KEYINPUT69), .B1(G150), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT68), .ZN(new_n280));
  INV_X1    g0080(.A(G58), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(KEYINPUT8), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT8), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G58), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n280), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT8), .B(G58), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n280), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n224), .A2(G33), .ZN(new_n290));
  OAI221_X1 g0090(.A(new_n279), .B1(KEYINPUT69), .B2(new_n277), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n223), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n292), .B(new_n223), .C1(G1), .C2(new_n224), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G50), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n208), .A2(G1), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G20), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n294), .B(new_n297), .C1(G50), .C2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT9), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n300), .B(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT10), .B1(new_n276), .B2(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n300), .B(KEYINPUT9), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT10), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n304), .A2(new_n305), .A3(new_n275), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  OR2_X1    g0107(.A1(new_n272), .A2(G179), .ZN(new_n308));
  INV_X1    g0108(.A(G169), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n272), .A2(new_n309), .ZN(new_n310));
  AND3_X1   g0110(.A1(new_n308), .A2(new_n300), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT77), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n249), .A2(G232), .A3(new_n255), .A4(new_n251), .ZN(new_n315));
  NOR2_X1   g0115(.A1(G223), .A2(G1698), .ZN(new_n316));
  INV_X1    g0116(.A(G226), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n316), .B1(new_n317), .B2(G1698), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n318), .A2(new_n263), .B1(G33), .B2(G87), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n256), .B(new_n315), .C1(new_n319), .C2(new_n262), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT75), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n317), .A2(G1698), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(G223), .B2(G1698), .ZN(new_n324));
  AND2_X1   g0124(.A1(KEYINPUT3), .A2(G33), .ZN(new_n325));
  NOR2_X1   g0125(.A1(KEYINPUT3), .A2(G33), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G33), .ZN(new_n328));
  INV_X1    g0128(.A(G87), .ZN(new_n329));
  OAI22_X1  g0129(.A1(new_n324), .A2(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n261), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n331), .A2(KEYINPUT75), .A3(new_n256), .A4(new_n315), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n322), .A2(new_n332), .ZN(new_n333));
  AND2_X1   g0133(.A1(KEYINPUT76), .A2(G190), .ZN(new_n334));
  NOR2_X1   g0134(.A1(KEYINPUT76), .A2(G190), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  OAI22_X1  g0137(.A1(new_n333), .A2(G200), .B1(new_n320), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n282), .A2(new_n284), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n339), .A2(KEYINPUT68), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n299), .B1(new_n340), .B2(new_n285), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT74), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n286), .A2(new_n288), .A3(new_n295), .ZN(new_n343));
  AND3_X1   g0143(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n342), .B1(new_n341), .B2(new_n343), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT7), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(new_n263), .B2(G20), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n327), .A2(KEYINPUT7), .A3(new_n224), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(new_n349), .A3(KEYINPUT73), .ZN(new_n350));
  NOR4_X1   g0150(.A1(new_n325), .A2(new_n326), .A3(new_n347), .A4(G20), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT73), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n350), .A2(G68), .A3(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n281), .A2(new_n242), .ZN(new_n355));
  OR2_X1    g0155(.A1(new_n355), .A2(new_n201), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n356), .A2(G20), .B1(G159), .B2(new_n278), .ZN(new_n357));
  AOI21_X1  g0157(.A(KEYINPUT16), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(KEYINPUT7), .B1(new_n327), .B2(new_n224), .ZN(new_n360));
  OAI21_X1  g0160(.A(G68), .B1(new_n360), .B2(new_n351), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n361), .A2(KEYINPUT16), .A3(new_n357), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n293), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n346), .B1(new_n359), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(KEYINPUT17), .B1(new_n338), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n322), .A2(new_n332), .ZN(new_n367));
  INV_X1    g0167(.A(G200), .ZN(new_n368));
  INV_X1    g0168(.A(new_n320), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n367), .A2(new_n368), .B1(new_n369), .B2(new_n336), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n341), .A2(new_n343), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(KEYINPUT74), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n341), .A2(new_n343), .A3(new_n342), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n358), .B2(new_n363), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT17), .ZN(new_n376));
  NOR3_X1   g0176(.A1(new_n370), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n314), .B1(new_n366), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G179), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n367), .A2(new_n309), .B1(new_n379), .B2(new_n369), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT18), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(new_n375), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n381), .B1(new_n380), .B2(new_n375), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n338), .A2(new_n365), .A3(KEYINPUT17), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n376), .B1(new_n370), .B2(new_n375), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n386), .A2(new_n387), .A3(KEYINPUT77), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n378), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n278), .A2(G50), .B1(G20), .B2(new_n242), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(new_n266), .B2(new_n290), .ZN(new_n391));
  AND2_X1   g0191(.A1(new_n391), .A2(new_n293), .ZN(new_n392));
  OR2_X1    g0192(.A1(new_n392), .A2(KEYINPUT11), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n391), .A2(KEYINPUT11), .A3(new_n293), .ZN(new_n394));
  OR3_X1    g0194(.A1(new_n299), .A2(KEYINPUT12), .A3(G68), .ZN(new_n395));
  OAI21_X1  g0195(.A(KEYINPUT12), .B1(new_n299), .B2(G68), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n395), .A2(new_n396), .B1(G68), .B2(new_n296), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n393), .A2(new_n394), .A3(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G97), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n328), .A2(new_n400), .ZN(new_n401));
  MUX2_X1   g0201(.A(G226), .B(G232), .S(G1698), .Z(new_n402));
  AOI21_X1  g0202(.A(new_n401), .B1(new_n402), .B2(new_n263), .ZN(new_n403));
  OR2_X1    g0203(.A1(new_n403), .A2(new_n262), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n258), .A2(G238), .A3(new_n251), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(new_n256), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT13), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT13), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n404), .A2(new_n408), .A3(new_n256), .A4(new_n405), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n410), .A2(KEYINPUT71), .A3(G200), .ZN(new_n411));
  AOI21_X1  g0211(.A(KEYINPUT71), .B1(new_n410), .B2(G200), .ZN(new_n412));
  OAI221_X1 g0212(.A(new_n399), .B1(new_n273), .B2(new_n410), .C1(new_n411), .C2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT72), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT14), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n410), .A2(G169), .A3(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n416), .B1(new_n379), .B2(new_n410), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n415), .B1(new_n410), .B2(G169), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n398), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n413), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n293), .ZN(new_n421));
  XNOR2_X1  g0221(.A(KEYINPUT15), .B(G87), .ZN(new_n422));
  OR2_X1    g0222(.A1(new_n422), .A2(new_n290), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n339), .A2(new_n278), .B1(G20), .B2(G77), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n421), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NOR3_X1   g0225(.A1(new_n208), .A2(new_n224), .A3(G1), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n266), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(new_n266), .B2(new_n295), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n257), .B1(new_n259), .B2(G244), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n270), .A2(G232), .ZN(new_n431));
  INV_X1    g0231(.A(G107), .ZN(new_n432));
  INV_X1    g0232(.A(G238), .ZN(new_n433));
  OAI221_X1 g0233(.A(new_n431), .B1(new_n432), .B2(new_n263), .C1(new_n433), .C2(new_n264), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n261), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n430), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT70), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n430), .A2(new_n435), .A3(KEYINPUT70), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n429), .B1(new_n440), .B2(new_n379), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n438), .A2(new_n309), .A3(new_n439), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n273), .B1(new_n438), .B2(new_n439), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n429), .B1(new_n440), .B2(new_n368), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NOR4_X1   g0246(.A1(new_n313), .A2(new_n389), .A3(new_n420), .A4(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(G1698), .ZN(new_n448));
  OAI211_X1 g0248(.A(G244), .B(new_n448), .C1(new_n325), .C2(new_n326), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT4), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n263), .A2(KEYINPUT4), .A3(G244), .A4(new_n448), .ZN(new_n452));
  NAND2_X1  g0252(.A1(G33), .A2(G283), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n263), .A2(G250), .A3(G1698), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n451), .A2(new_n452), .A3(new_n453), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n261), .ZN(new_n456));
  INV_X1    g0256(.A(G45), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(G1), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT5), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(G41), .ZN(new_n460));
  INV_X1    g0260(.A(G41), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT5), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n458), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  AND4_X1   g0263(.A1(G257), .A2(new_n463), .A3(new_n249), .A4(new_n255), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n250), .B(G45), .C1(new_n461), .C2(KEYINPUT5), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT78), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n458), .A2(KEYINPUT78), .A3(new_n460), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n468), .A2(new_n462), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n249), .A2(G274), .A3(new_n255), .ZN(new_n471));
  OR2_X1    g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AND4_X1   g0272(.A1(G179), .A2(new_n456), .A3(new_n465), .A4(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n464), .B1(new_n455), .B2(new_n261), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n309), .B1(new_n474), .B2(new_n472), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n350), .A2(G107), .A3(new_n353), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n432), .A2(KEYINPUT6), .A3(G97), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n400), .A2(new_n432), .ZN(new_n478));
  NOR2_X1   g0278(.A1(G97), .A2(G107), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n477), .B1(new_n480), .B2(KEYINPUT6), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n481), .A2(G20), .B1(G77), .B2(new_n278), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n421), .B1(new_n476), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n426), .A2(new_n400), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n328), .A2(G1), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n421), .A2(new_n299), .A3(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n484), .B1(new_n487), .B2(new_n400), .ZN(new_n488));
  OAI22_X1  g0288(.A1(new_n473), .A2(new_n475), .B1(new_n483), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n476), .A2(new_n482), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n488), .B1(new_n490), .B2(new_n293), .ZN(new_n491));
  AND4_X1   g0291(.A1(new_n273), .A2(new_n456), .A3(new_n465), .A4(new_n472), .ZN(new_n492));
  AOI21_X1  g0292(.A(G200), .B1(new_n474), .B2(new_n472), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(G20), .B1(new_n401), .B2(KEYINPUT19), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  AND2_X1   g0297(.A1(KEYINPUT79), .A2(G87), .ZN(new_n498));
  NOR2_X1   g0298(.A1(KEYINPUT79), .A2(G87), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(KEYINPUT80), .B1(new_n500), .B2(new_n479), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT79), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n329), .ZN(new_n503));
  NAND2_X1  g0303(.A1(KEYINPUT79), .A2(G87), .ZN(new_n504));
  AND4_X1   g0304(.A1(KEYINPUT80), .A2(new_n503), .A3(new_n479), .A4(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n497), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n263), .A2(new_n224), .A3(G68), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT19), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(new_n290), .B2(new_n400), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n511), .A2(new_n293), .B1(new_n426), .B2(new_n422), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n426), .A2(new_n293), .A3(new_n485), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G87), .ZN(new_n514));
  OAI211_X1 g0314(.A(G238), .B(new_n448), .C1(new_n325), .C2(new_n326), .ZN(new_n515));
  OAI211_X1 g0315(.A(G244), .B(G1698), .C1(new_n325), .C2(new_n326), .ZN(new_n516));
  NAND2_X1  g0316(.A1(G33), .A2(G116), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n261), .ZN(new_n519));
  AOI21_X1  g0319(.A(G250), .B1(new_n250), .B2(G45), .ZN(new_n520));
  INV_X1    g0320(.A(G274), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n520), .B1(new_n521), .B2(new_n458), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n258), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(G200), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n519), .A2(new_n523), .A3(G190), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n512), .A2(new_n514), .A3(new_n525), .A4(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n503), .A2(new_n479), .A3(new_n504), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT80), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n500), .A2(KEYINPUT80), .A3(new_n479), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n496), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n507), .A2(new_n509), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n293), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n422), .A2(new_n426), .ZN(new_n535));
  OR2_X1    g0335(.A1(new_n487), .A2(new_n422), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n261), .A2(new_n518), .B1(new_n258), .B2(new_n522), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n379), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n524), .A2(new_n309), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n537), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT81), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n527), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n542), .B1(new_n527), .B2(new_n541), .ZN(new_n544));
  NOR3_X1   g0344(.A1(new_n495), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT21), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n463), .A2(new_n249), .A3(G270), .A4(new_n255), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(new_n470), .B2(new_n471), .ZN(new_n548));
  OAI211_X1 g0348(.A(G264), .B(G1698), .C1(new_n325), .C2(new_n326), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT82), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n263), .A2(KEYINPUT82), .A3(G264), .A4(G1698), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n327), .A2(G303), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n263), .A2(G257), .A3(new_n448), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n551), .A2(new_n552), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n548), .B1(new_n261), .B2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(G116), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n292), .A2(new_n223), .B1(G20), .B2(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n453), .B(new_n224), .C1(G33), .C2(new_n400), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n558), .A2(KEYINPUT20), .A3(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(KEYINPUT20), .B1(new_n558), .B2(new_n559), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n426), .A2(new_n557), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n487), .B2(new_n557), .ZN(new_n565));
  OAI21_X1  g0365(.A(G169), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n546), .B1(new_n556), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n562), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n560), .ZN(new_n569));
  INV_X1    g0369(.A(new_n564), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n570), .B1(new_n513), .B2(G116), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n556), .A2(G179), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n548), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n555), .A2(new_n261), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n309), .B1(new_n569), .B2(new_n571), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n576), .A2(new_n577), .A3(KEYINPUT21), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n567), .A2(new_n573), .A3(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n572), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(new_n576), .B2(new_n336), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n368), .B1(new_n574), .B2(new_n575), .ZN(new_n582));
  NOR3_X1   g0382(.A1(new_n581), .A2(KEYINPUT83), .A3(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT83), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n572), .B1(new_n556), .B2(new_n337), .ZN(new_n585));
  INV_X1    g0385(.A(new_n582), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n579), .B1(new_n583), .B2(new_n587), .ZN(new_n588));
  OAI211_X1 g0388(.A(G250), .B(new_n448), .C1(new_n325), .C2(new_n326), .ZN(new_n589));
  NAND2_X1  g0389(.A1(G33), .A2(G294), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n263), .A2(G257), .A3(G1698), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n262), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n463), .A2(new_n249), .A3(G264), .A4(new_n255), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n470), .B2(new_n471), .ZN(new_n595));
  OAI211_X1 g0395(.A(KEYINPUT86), .B(G169), .C1(new_n593), .C2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n592), .A2(new_n590), .A3(new_n589), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n261), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n472), .A2(new_n598), .A3(new_n594), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n596), .B1(new_n379), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(KEYINPUT86), .B1(new_n599), .B2(G169), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n224), .B(G87), .C1(new_n325), .C2(new_n326), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT84), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n602), .A2(new_n603), .A3(KEYINPUT22), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(KEYINPUT22), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n263), .A2(new_n224), .A3(G87), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n517), .A2(G20), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n224), .A2(G107), .ZN(new_n609));
  OR2_X1    g0409(.A1(new_n609), .A2(KEYINPUT23), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(KEYINPUT23), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n608), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT24), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT24), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n607), .A2(new_n615), .A3(new_n612), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n421), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n298), .A2(new_n609), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n618), .A2(KEYINPUT85), .A3(KEYINPUT25), .ZN(new_n619));
  OR2_X1    g0419(.A1(KEYINPUT85), .A2(KEYINPUT25), .ZN(new_n620));
  NAND2_X1  g0420(.A1(KEYINPUT85), .A2(KEYINPUT25), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n298), .A2(new_n609), .A3(new_n620), .A4(new_n621), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n619), .B(new_n622), .C1(new_n487), .C2(new_n432), .ZN(new_n623));
  OAI22_X1  g0423(.A1(new_n600), .A2(new_n601), .B1(new_n617), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n368), .B1(new_n593), .B2(new_n595), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n625), .B1(new_n599), .B2(G190), .ZN(new_n626));
  INV_X1    g0426(.A(new_n616), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n615), .B1(new_n607), .B2(new_n612), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n293), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n623), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n626), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n624), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n588), .A2(new_n632), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n447), .A2(new_n545), .A3(new_n633), .ZN(G372));
  NAND2_X1  g0434(.A1(new_n380), .A2(new_n375), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(KEYINPUT18), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n382), .ZN(new_n637));
  INV_X1    g0437(.A(new_n443), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n413), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n419), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n386), .A2(KEYINPUT77), .A3(new_n387), .ZN(new_n641));
  AOI21_X1  g0441(.A(KEYINPUT77), .B1(new_n386), .B2(new_n387), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n637), .B1(new_n640), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n307), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n312), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n540), .A2(new_n539), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n526), .B1(new_n538), .B2(new_n368), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n534), .A2(new_n535), .A3(new_n514), .ZN(new_n651));
  OAI22_X1  g0451(.A1(new_n648), .A2(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(KEYINPUT81), .ZN(new_n653));
  INV_X1    g0453(.A(new_n489), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n527), .A2(new_n541), .A3(new_n542), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(KEYINPUT26), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n512), .A2(new_n514), .A3(new_n526), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT87), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(new_n538), .B2(new_n368), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n524), .A2(KEYINPUT87), .A3(G200), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n541), .B1(new_n658), .B2(new_n662), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n626), .A2(new_n629), .A3(new_n630), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n579), .A2(new_n624), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n489), .A2(new_n494), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n475), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n474), .A2(G179), .A3(new_n472), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT88), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n491), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n663), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT26), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n669), .A2(KEYINPUT88), .A3(new_n670), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n673), .A2(new_n674), .A3(new_n675), .A4(new_n676), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n657), .A2(new_n668), .A3(new_n677), .A4(new_n541), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n447), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n647), .A2(new_n679), .ZN(G369));
  NAND2_X1  g0480(.A1(new_n298), .A2(new_n224), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT89), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT89), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n681), .B(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT27), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n683), .A2(new_n687), .A3(G213), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(G343), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(new_n580), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n567), .A2(new_n578), .A3(new_n573), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n693), .A2(KEYINPUT90), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(KEYINPUT90), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n694), .B(new_n695), .C1(new_n588), .C2(new_n691), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n690), .B1(new_n629), .B2(new_n630), .ZN(new_n698));
  OAI22_X1  g0498(.A1(new_n632), .A2(new_n698), .B1(new_n624), .B2(new_n690), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n692), .A2(new_n690), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n702), .A2(new_n624), .A3(new_n631), .ZN(new_n703));
  INV_X1    g0503(.A(new_n690), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n624), .A2(new_n704), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n700), .A2(new_n706), .ZN(G399));
  NOR2_X1   g0507(.A1(new_n501), .A2(new_n505), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n557), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n209), .A2(G41), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n710), .A2(new_n712), .A3(G1), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n226), .A2(G50), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n713), .B1(new_n714), .B2(new_n712), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT28), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT29), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n678), .A2(new_n717), .A3(new_n690), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT93), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n666), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n579), .A2(new_n624), .A3(KEYINPUT93), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n720), .A2(new_n667), .A3(new_n665), .A4(new_n721), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n722), .A2(new_n541), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n656), .A2(new_n675), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(KEYINPUT92), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n673), .A2(new_n674), .A3(KEYINPUT26), .A4(new_n676), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT92), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n656), .A2(new_n727), .A3(new_n675), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n725), .A2(new_n726), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n704), .B1(new_n723), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n718), .B1(new_n730), .B2(new_n717), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT30), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n556), .A2(G179), .ZN(new_n733));
  INV_X1    g0533(.A(new_n595), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n474), .A2(new_n538), .A3(new_n598), .A4(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n732), .B1(new_n733), .B2(new_n735), .ZN(new_n736));
  AND3_X1   g0536(.A1(new_n574), .A2(new_n575), .A3(G179), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n524), .A2(new_n593), .A3(new_n595), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n737), .A2(new_n738), .A3(KEYINPUT30), .A4(new_n474), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n474), .A2(new_n472), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n538), .A2(G179), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n740), .A2(new_n599), .A3(new_n576), .A4(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n736), .A2(new_n739), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n704), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT31), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n743), .A2(KEYINPUT31), .A3(new_n704), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AND4_X1   g0549(.A1(new_n667), .A2(new_n655), .A3(new_n653), .A4(new_n690), .ZN(new_n750));
  AOI21_X1  g0550(.A(KEYINPUT91), .B1(new_n750), .B2(new_n633), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n667), .A2(new_n655), .A3(new_n653), .A4(new_n690), .ZN(new_n752));
  OAI21_X1  g0552(.A(KEYINPUT83), .B1(new_n581), .B2(new_n582), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n585), .A2(new_n586), .A3(new_n584), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n755), .A2(new_n624), .A3(new_n631), .A4(new_n579), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT91), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n752), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n749), .B1(new_n751), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n731), .B1(G330), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n716), .B1(new_n760), .B2(G1), .ZN(G364));
  NOR2_X1   g0561(.A1(new_n208), .A2(G20), .ZN(new_n762));
  AOI21_X1  g0562(.A(KEYINPUT94), .B1(new_n762), .B2(G45), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n250), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n762), .A2(KEYINPUT94), .A3(G45), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n711), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n697), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(G330), .B2(new_n696), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G13), .A2(G33), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n223), .B1(G20), .B2(new_n309), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n209), .A2(new_n327), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT95), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n776), .A2(G355), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n209), .A2(new_n263), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(G45), .B2(new_n714), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n246), .A2(new_n457), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n779), .A2(new_n780), .B1(G116), .B2(new_n210), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n774), .B1(new_n777), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(new_n767), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G179), .A2(G200), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(G20), .B1(new_n785), .B2(new_n273), .ZN(new_n786));
  INV_X1    g0586(.A(KEYINPUT96), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT98), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n224), .A2(G179), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n793), .A2(G190), .A3(G200), .ZN(new_n794));
  INV_X1    g0594(.A(G303), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n327), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n791), .A2(G294), .B1(new_n792), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(new_n792), .B2(new_n796), .ZN(new_n798));
  NOR3_X1   g0598(.A1(new_n785), .A2(new_n224), .A3(G190), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G329), .ZN(new_n800));
  NAND3_X1  g0600(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n336), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  XOR2_X1   g0603(.A(KEYINPUT97), .B(G326), .Z(new_n804));
  OAI21_X1  g0604(.A(new_n800), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n793), .A2(new_n273), .A3(G200), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n801), .A2(G190), .ZN(new_n808));
  XNOR2_X1  g0608(.A(KEYINPUT33), .B(G317), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n807), .A2(G283), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(G311), .ZN(new_n811));
  NOR3_X1   g0611(.A1(new_n224), .A2(new_n379), .A3(G200), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n273), .ZN(new_n813));
  INV_X1    g0613(.A(G322), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n337), .A2(new_n812), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n810), .B1(new_n811), .B2(new_n813), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  NOR3_X1   g0616(.A1(new_n798), .A2(new_n805), .A3(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n818), .A2(KEYINPUT99), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(KEYINPUT99), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT32), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(new_n799), .B2(G159), .ZN(new_n822));
  INV_X1    g0622(.A(new_n799), .ZN(new_n823));
  INV_X1    g0623(.A(G159), .ZN(new_n824));
  NOR3_X1   g0624(.A1(new_n823), .A2(KEYINPUT32), .A3(new_n824), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n822), .B(new_n825), .C1(G107), .C2(new_n807), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n327), .B1(new_n802), .B2(G50), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n815), .A2(new_n281), .B1(new_n266), .B2(new_n813), .ZN(new_n828));
  INV_X1    g0628(.A(new_n808), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n829), .A2(new_n242), .B1(new_n794), .B2(new_n500), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n791), .A2(G97), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n826), .A2(new_n827), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n819), .A2(new_n820), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n783), .B1(new_n834), .B2(new_n773), .ZN(new_n835));
  INV_X1    g0635(.A(new_n772), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n835), .B1(new_n696), .B2(new_n836), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n769), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(G396));
  NOR2_X1   g0639(.A1(new_n773), .A2(new_n770), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n815), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n842), .A2(G143), .B1(G150), .B2(new_n808), .ZN(new_n843));
  INV_X1    g0643(.A(new_n813), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n844), .A2(G159), .B1(new_n802), .B2(G137), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n846), .A2(KEYINPUT34), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(KEYINPUT34), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n327), .B1(new_n799), .B2(G132), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n849), .B1(new_n202), .B2(new_n794), .C1(new_n242), .C2(new_n806), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(G58), .B2(new_n791), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n847), .A2(new_n848), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n327), .B1(new_n823), .B2(new_n811), .ZN(new_n853));
  INV_X1    g0653(.A(G283), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n803), .A2(new_n795), .B1(new_n854), .B2(new_n829), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n853), .B(new_n855), .C1(G116), .C2(new_n844), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n806), .A2(new_n329), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n794), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n842), .A2(G294), .B1(G107), .B2(new_n859), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n856), .A2(new_n832), .A3(new_n858), .A4(new_n860), .ZN(new_n861));
  AND2_X1   g0661(.A1(new_n852), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n773), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n767), .B1(G77), .B2(new_n841), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n429), .ZN(new_n865));
  INV_X1    g0665(.A(new_n439), .ZN(new_n866));
  AOI21_X1  g0666(.A(KEYINPUT70), .B1(new_n430), .B2(new_n435), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n379), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AND4_X1   g0668(.A1(new_n865), .A2(new_n868), .A3(new_n442), .A4(new_n690), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n704), .A2(new_n865), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n445), .B2(new_n444), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n869), .B1(new_n871), .B2(new_n443), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n864), .B1(new_n873), .B2(new_n770), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n678), .A2(new_n690), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n873), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n678), .A2(new_n872), .A3(new_n690), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n759), .A2(G330), .ZN(new_n879));
  OR2_X1    g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n767), .B1(new_n878), .B2(new_n879), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n874), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(G384));
  INV_X1    g0683(.A(KEYINPUT40), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n759), .A2(KEYINPUT100), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n399), .A2(new_n690), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n413), .A2(new_n419), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n887), .B1(new_n413), .B2(new_n419), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n872), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n633), .A2(new_n545), .A3(KEYINPUT91), .A4(new_n690), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n757), .B1(new_n752), .B2(new_n756), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n748), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT100), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n885), .A2(new_n891), .A3(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT38), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n338), .A2(new_n365), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT37), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n375), .A2(new_n689), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n899), .A2(new_n900), .A3(new_n635), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n361), .A2(new_n357), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT16), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n346), .B1(new_n364), .B2(new_n905), .ZN(new_n906));
  OAI22_X1  g0706(.A1(new_n906), .A2(new_n688), .B1(new_n370), .B2(new_n375), .ZN(new_n907));
  OAI22_X1  g0707(.A1(new_n333), .A2(G169), .B1(G179), .B2(new_n320), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n908), .A2(new_n906), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT37), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n906), .A2(new_n688), .ZN(new_n911));
  AOI221_X4 g0711(.A(new_n898), .B1(new_n902), .B2(new_n910), .C1(new_n389), .C2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n389), .A2(new_n911), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n910), .A2(new_n902), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT38), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n884), .B1(new_n897), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n913), .A2(KEYINPUT38), .A3(new_n914), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n899), .A2(new_n635), .A3(new_n901), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(KEYINPUT37), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n902), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n636), .A2(new_n386), .A3(new_n382), .A4(new_n387), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n922), .A2(new_n375), .A3(new_n689), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n898), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n884), .B1(new_n918), .B2(new_n925), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n926), .A2(new_n891), .A3(new_n885), .A4(new_n896), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n917), .A2(new_n927), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n447), .A2(new_n885), .A3(new_n896), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n928), .A2(new_n929), .ZN(new_n931));
  INV_X1    g0731(.A(G330), .ZN(new_n932));
  NOR3_X1   g0732(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n869), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n877), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n888), .A2(new_n889), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n916), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n637), .B2(new_n688), .ZN(new_n940));
  INV_X1    g0740(.A(new_n915), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n941), .A2(KEYINPUT39), .A3(new_n918), .ZN(new_n942));
  AOI21_X1  g0742(.A(KEYINPUT39), .B1(new_n918), .B2(new_n925), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n419), .A2(new_n704), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n942), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n940), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n646), .B1(new_n731), .B2(new_n447), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n948), .B(new_n949), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n933), .A2(new_n950), .B1(new_n250), .B2(new_n762), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(new_n950), .B2(new_n933), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n481), .A2(KEYINPUT35), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n481), .A2(KEYINPUT35), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n953), .A2(new_n954), .A3(G116), .A4(new_n225), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT36), .Z(new_n956));
  OR3_X1    g0756(.A1(new_n714), .A2(new_n266), .A3(new_n355), .ZN(new_n957));
  AOI211_X1 g0757(.A(new_n250), .B(G13), .C1(new_n957), .C2(new_n241), .ZN(new_n958));
  OR3_X1    g0758(.A1(new_n952), .A2(new_n956), .A3(new_n958), .ZN(G367));
  NOR3_X1   g0759(.A1(new_n236), .A2(new_n209), .A3(new_n263), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n774), .B1(new_n210), .B2(new_n422), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n767), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n799), .A2(G137), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n327), .B(new_n963), .C1(G143), .C2(new_n802), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n791), .A2(G68), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n829), .A2(new_n824), .B1(new_n806), .B2(new_n266), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(G50), .B2(new_n844), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n842), .A2(G150), .B1(G58), .B2(new_n859), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n964), .A2(new_n965), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(G317), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n327), .B1(new_n400), .B2(new_n806), .C1(new_n823), .C2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(KEYINPUT105), .B1(new_n794), .B2(new_n557), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n971), .A2(KEYINPUT106), .B1(KEYINPUT46), .B2(new_n972), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n973), .B1(KEYINPUT106), .B2(new_n971), .C1(new_n432), .C2(new_n790), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n842), .A2(G303), .B1(G294), .B2(new_n808), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n844), .A2(G283), .B1(new_n802), .B2(G311), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n975), .B(new_n976), .C1(KEYINPUT46), .C2(new_n972), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n969), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT47), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n962), .B1(new_n979), .B2(new_n773), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n704), .A2(new_n651), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n981), .A2(new_n541), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n674), .A2(new_n981), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n772), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n980), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n703), .B1(new_n699), .B2(new_n702), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n697), .B(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n760), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT44), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n667), .B1(new_n491), .B2(new_n690), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n673), .A2(new_n676), .A3(new_n704), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n991), .B1(new_n706), .B2(new_n994), .ZN(new_n995));
  AND2_X1   g0795(.A1(new_n992), .A2(new_n993), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n703), .A2(new_n705), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n996), .A2(KEYINPUT44), .A3(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT45), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n996), .B2(new_n997), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n706), .A2(KEYINPUT45), .A3(new_n994), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n995), .A2(new_n998), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(KEYINPUT103), .B1(new_n1002), .B2(new_n700), .ZN(new_n1003));
  AND2_X1   g0803(.A1(new_n697), .A2(new_n699), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n995), .A2(new_n998), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT103), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1004), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1002), .A2(new_n700), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1003), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n760), .B1(new_n990), .B2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n711), .B(KEYINPUT41), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(KEYINPUT104), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT104), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1012), .A2(new_n1016), .A3(new_n1013), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n766), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n996), .A2(new_n703), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(KEYINPUT42), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n489), .B1(new_n996), .B2(new_n624), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n690), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n1023), .A2(KEYINPUT101), .B1(KEYINPUT42), .B2(new_n1019), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT101), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT43), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1027), .A2(new_n1028), .A3(new_n985), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n985), .A2(new_n1028), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1030), .B(new_n1031), .C1(new_n1024), .C2(new_n1026), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n700), .A2(new_n996), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1029), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(KEYINPUT102), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT102), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1029), .A2(new_n1032), .A3(new_n1036), .A4(new_n1033), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1033), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1035), .A2(new_n1037), .A3(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n987), .B1(new_n1018), .B2(new_n1041), .ZN(G387));
  NOR2_X1   g0842(.A1(new_n287), .A2(G50), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT50), .ZN(new_n1044));
  AOI21_X1  g0844(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n710), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1046), .B(new_n778), .C1(new_n233), .C2(new_n457), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n776), .A2(new_n709), .B1(new_n432), .B2(new_n209), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1049), .A2(KEYINPUT107), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(KEYINPUT107), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n774), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n844), .A2(G68), .B1(new_n859), .B2(G77), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1053), .B1(new_n202), .B2(new_n815), .C1(new_n824), .C2(new_n803), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n790), .A2(new_n422), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n327), .B1(new_n799), .B2(G150), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1056), .B1(new_n400), .B2(new_n806), .C1(new_n289), .C2(new_n829), .ZN(new_n1057));
  NOR3_X1   g0857(.A1(new_n1054), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n802), .A2(G322), .B1(G311), .B2(new_n808), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1059), .B1(new_n795), .B2(new_n813), .C1(new_n970), .C2(new_n815), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT48), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n791), .A2(G283), .B1(G294), .B2(new_n859), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT49), .Z(new_n1066));
  OR2_X1    g0866(.A1(new_n1066), .A2(KEYINPUT108), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n327), .B1(new_n557), .B2(new_n806), .C1(new_n823), .C2(new_n804), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n1066), .B2(KEYINPUT108), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1058), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n767), .B1(new_n1050), .B2(new_n1052), .C1(new_n1070), .C2(new_n863), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1071), .A2(KEYINPUT109), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n699), .A2(new_n836), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1071), .A2(KEYINPUT109), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n1074), .A2(new_n1075), .B1(new_n766), .B2(new_n989), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n760), .A2(new_n989), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n990), .A2(new_n711), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1076), .B1(new_n1077), .B2(new_n1078), .ZN(G393));
  INV_X1    g0879(.A(new_n767), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n774), .B1(new_n210), .B2(new_n400), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n240), .B2(new_n778), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n823), .A2(new_n814), .B1(new_n794), .B2(new_n854), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n791), .A2(G116), .B1(KEYINPUT110), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(G294), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n813), .A2(new_n1085), .B1(new_n829), .B2(new_n795), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n263), .B(new_n1086), .C1(G107), .C2(new_n807), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1084), .B(new_n1087), .C1(KEYINPUT110), .C2(new_n1083), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n842), .A2(G311), .B1(G317), .B2(new_n802), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT52), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n842), .A2(G159), .B1(G150), .B2(new_n802), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT51), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n791), .A2(G77), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n327), .B(new_n857), .C1(G143), .C2(new_n799), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n808), .A2(G50), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n844), .A2(new_n339), .B1(new_n859), .B2(G68), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n1088), .A2(new_n1090), .B1(new_n1092), .B2(new_n1097), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n1080), .B(new_n1082), .C1(new_n1098), .C2(new_n773), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n1099), .B(KEYINPUT111), .Z(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n836), .B2(new_n994), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n1010), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n766), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1101), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n990), .A2(new_n1011), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1106), .A2(new_n712), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n990), .A2(new_n1103), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1105), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(G390));
  AOI21_X1  g0910(.A(new_n946), .B1(new_n935), .B2(new_n937), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n944), .B2(new_n942), .ZN(new_n1112));
  AOI21_X1  g0912(.A(KEYINPUT38), .B1(new_n921), .B2(new_n923), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n945), .B1(new_n912), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n728), .A2(new_n726), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n727), .B1(new_n656), .B2(new_n675), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n541), .B(new_n722), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n871), .A2(new_n443), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1117), .A2(new_n690), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n934), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1114), .B1(new_n1120), .B2(new_n937), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n759), .A2(G330), .A3(new_n872), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1122), .A2(new_n936), .ZN(new_n1123));
  NOR3_X1   g0923(.A1(new_n1112), .A2(new_n1121), .A3(new_n1123), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n885), .A2(new_n891), .A3(G330), .A4(new_n896), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n938), .A2(new_n945), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT39), .ZN(new_n1127));
  NOR3_X1   g0927(.A1(new_n912), .A2(new_n915), .A3(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1126), .B1(new_n1128), .B2(new_n943), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n946), .B1(new_n918), .B2(new_n925), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n869), .B1(new_n730), .B2(new_n1118), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1130), .B1(new_n1131), .B2(new_n936), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1125), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1124), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n770), .B1(new_n1128), .B2(new_n943), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n841), .B1(new_n286), .B2(new_n288), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n803), .A2(new_n854), .B1(new_n329), .B2(new_n794), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(G116), .B2(new_n842), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n327), .B1(new_n823), .B2(new_n1085), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(G68), .B2(new_n807), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n844), .A2(G97), .B1(G107), .B2(new_n808), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1138), .A2(new_n1093), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n859), .A2(G150), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1143), .B(KEYINPUT53), .Z(new_n1144));
  OAI21_X1  g0944(.A(new_n1144), .B1(new_n824), .B2(new_n790), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n806), .A2(new_n202), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n327), .B(new_n1146), .C1(G125), .C2(new_n799), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n842), .A2(G132), .B1(G137), .B2(new_n808), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n802), .A2(G128), .ZN(new_n1149));
  XOR2_X1   g0949(.A(KEYINPUT54), .B(G143), .Z(new_n1150));
  XNOR2_X1  g0950(.A(new_n1150), .B(KEYINPUT114), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n844), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .A4(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1142), .B1(new_n1145), .B2(new_n1153), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n1080), .B(new_n1136), .C1(new_n1154), .C2(new_n773), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n1134), .A2(new_n766), .B1(new_n1135), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT113), .ZN(new_n1157));
  NOR3_X1   g0957(.A1(new_n894), .A2(new_n932), .A3(new_n873), .ZN(new_n1158));
  OAI21_X1  g0958(.A(KEYINPUT112), .B1(new_n1158), .B2(new_n937), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT112), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1122), .A2(new_n1160), .A3(new_n936), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1159), .A2(new_n1125), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n935), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n885), .A2(G330), .A3(new_n896), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n936), .B1(new_n1164), .B2(new_n873), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1123), .A2(new_n1120), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1163), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n731), .A2(new_n447), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n447), .A2(new_n885), .A3(G330), .A4(new_n896), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1169), .A2(new_n647), .A3(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1168), .A2(new_n1172), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1129), .B(new_n1132), .C1(new_n936), .C2(new_n1122), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1164), .A2(new_n890), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(new_n1112), .B2(new_n1121), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n712), .B1(new_n1173), .B2(new_n1177), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1168), .A2(new_n1174), .A3(new_n1176), .A4(new_n1172), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1157), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n935), .A2(new_n1162), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n1181), .A2(new_n1171), .B1(new_n1124), .B2(new_n1133), .ZN(new_n1182));
  AND4_X1   g0982(.A1(new_n1157), .A2(new_n1182), .A3(new_n1179), .A4(new_n711), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1156), .B1(new_n1180), .B2(new_n1183), .ZN(G378));
  INV_X1    g0984(.A(KEYINPUT115), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n894), .A2(new_n895), .ZN(new_n1186));
  AOI211_X1 g0986(.A(KEYINPUT100), .B(new_n748), .C1(new_n892), .C2(new_n893), .ZN(new_n1187));
  NOR3_X1   g0987(.A1(new_n1186), .A2(new_n1187), .A3(new_n890), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n916), .ZN(new_n1189));
  AOI21_X1  g0989(.A(KEYINPUT40), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n927), .A2(G330), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1185), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n932), .B1(new_n1188), .B2(new_n926), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1193), .A2(KEYINPUT115), .A3(new_n917), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n300), .A2(new_n689), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n313), .B(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1196), .B(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1192), .A2(new_n1194), .A3(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n948), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1198), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1201), .A2(KEYINPUT115), .A3(new_n1193), .A4(new_n917), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n1199), .A2(new_n1200), .A3(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1200), .B1(new_n1199), .B2(new_n1202), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1201), .A2(new_n770), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n767), .B1(G50), .B2(new_n841), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n263), .A2(G41), .ZN(new_n1208));
  AOI211_X1 g1008(.A(G50), .B(new_n1208), .C1(new_n328), .C2(new_n461), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n806), .A2(new_n281), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1208), .B1(new_n266), .B2(new_n794), .C1(new_n823), .C2(new_n854), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1210), .B(new_n1211), .C1(G97), .C2(new_n808), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n803), .A2(new_n557), .B1(new_n422), .B2(new_n813), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G107), .B2(new_n842), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1212), .A2(new_n965), .A3(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT58), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1209), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n791), .A2(G150), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1151), .A2(new_n859), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n844), .A2(G137), .B1(new_n802), .B2(G125), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n842), .A2(G128), .B1(G132), .B2(new_n808), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1222), .A2(KEYINPUT59), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(KEYINPUT59), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n807), .A2(G159), .ZN(new_n1225));
  AOI211_X1 g1025(.A(G33), .B(G41), .C1(new_n799), .C2(G124), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1217), .B1(new_n1216), .B2(new_n1215), .C1(new_n1223), .C2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1207), .B1(new_n1228), .B2(new_n773), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1205), .A2(new_n766), .B1(new_n1206), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT116), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1171), .A2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n949), .A2(KEYINPUT116), .A3(new_n1170), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1171), .B1(new_n1163), .B2(new_n1167), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1234), .B1(new_n1134), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(KEYINPUT57), .B1(new_n1205), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT57), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1234), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1239), .B1(new_n1179), .B2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1199), .A2(new_n1202), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n948), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1199), .A2(new_n1200), .A3(new_n1202), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1241), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n711), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1230), .B1(new_n1238), .B2(new_n1246), .ZN(G375));
  XNOR2_X1  g1047(.A(new_n766), .B(KEYINPUT117), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1168), .A2(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n767), .B1(G68), .B2(new_n841), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1250), .B(KEYINPUT118), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n813), .A2(new_n432), .B1(new_n794), .B2(new_n400), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n327), .B1(new_n823), .B2(new_n795), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n1252), .B(new_n1253), .C1(G77), .C2(new_n807), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n802), .A2(G294), .B1(G116), .B2(new_n808), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1254), .B(new_n1255), .C1(new_n854), .C2(new_n815), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n790), .A2(new_n202), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n327), .B(new_n1210), .C1(G128), .C2(new_n799), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n842), .A2(G137), .B1(G132), .B2(new_n802), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n844), .A2(G150), .B1(new_n859), .B2(G159), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1151), .A2(new_n808), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1258), .A2(new_n1259), .A3(new_n1260), .A4(new_n1261), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n1256), .A2(new_n1055), .B1(new_n1257), .B2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1251), .B1(new_n1263), .B2(new_n773), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n937), .B2(new_n771), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1249), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1173), .A2(new_n1013), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1168), .A2(new_n1172), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1267), .B1(new_n1268), .B2(new_n1269), .ZN(G381));
  INV_X1    g1070(.A(KEYINPUT119), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(G375), .B(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1109), .A2(new_n882), .ZN(new_n1273));
  OR3_X1    g1073(.A1(new_n1273), .A2(G396), .A3(G393), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1156), .ZN(new_n1276));
  OR4_X1    g1076(.A1(G387), .A2(new_n1274), .A3(G381), .A4(new_n1276), .ZN(new_n1277));
  OR2_X1    g1077(.A1(new_n1272), .A2(new_n1277), .ZN(G407));
  INV_X1    g1078(.A(G343), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(G213), .ZN(new_n1280));
  OR3_X1    g1080(.A1(new_n1272), .A2(new_n1276), .A3(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1281), .A2(G213), .A3(G407), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT120), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1281), .A2(KEYINPUT120), .A3(G213), .A4(G407), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(G409));
  AOI21_X1  g1086(.A(KEYINPUT123), .B1(G387), .B2(new_n1109), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(G393), .B(new_n838), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n987), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n1035), .A2(new_n1037), .A3(new_n1040), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1012), .A2(new_n1016), .A3(new_n1013), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1016), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1104), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1290), .B1(new_n1291), .B2(new_n1294), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1295), .A2(G390), .ZN(new_n1296));
  AOI211_X1 g1096(.A(new_n1290), .B(new_n1109), .C1(new_n1291), .C2(new_n1294), .ZN(new_n1297));
  OAI22_X1  g1097(.A1(new_n1287), .A2(new_n1289), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT61), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(G387), .A2(new_n1109), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1295), .A2(G390), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1300), .A2(new_n1301), .A3(KEYINPUT123), .A4(new_n1288), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1298), .A2(new_n1299), .A3(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1280), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1205), .A2(new_n1013), .A3(new_n1237), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1206), .A2(new_n1229), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1205), .A2(new_n1248), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1305), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1276), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  OAI211_X1 g1110(.A(G378), .B(new_n1230), .C1(new_n1238), .C2(new_n1246), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1304), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1173), .A2(KEYINPUT60), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1313), .B1(new_n1172), .B2(new_n1168), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1181), .A2(KEYINPUT60), .A3(new_n1171), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1314), .A2(new_n711), .A3(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n1267), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n882), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1316), .A2(G384), .A3(new_n1267), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1312), .A2(KEYINPUT63), .A3(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1303), .A2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(KEYINPUT121), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT121), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1310), .A2(new_n1311), .A3(new_n1326), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1325), .A2(new_n1280), .A3(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1304), .A2(G2897), .ZN(new_n1329));
  AND2_X1   g1129(.A1(new_n1320), .A2(new_n1329), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1320), .A2(new_n1329), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1323), .B1(new_n1328), .B2(new_n1333), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1325), .A2(new_n1280), .A3(new_n1321), .A4(new_n1327), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT63), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT122), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1335), .A2(KEYINPUT122), .A3(new_n1336), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1334), .A2(new_n1339), .A3(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1298), .A2(new_n1302), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT62), .ZN(new_n1343));
  NOR2_X1   g1143(.A1(new_n1320), .A2(new_n1343), .ZN(new_n1344));
  AOI22_X1  g1144(.A1(new_n1335), .A2(new_n1343), .B1(new_n1312), .B2(new_n1344), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1299), .B1(new_n1332), .B2(new_n1312), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1342), .B1(new_n1345), .B2(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1341), .A2(new_n1347), .ZN(G405));
  INV_X1    g1148(.A(KEYINPUT125), .ZN(new_n1349));
  NOR3_X1   g1149(.A1(new_n1203), .A2(new_n1204), .A3(new_n1236), .ZN(new_n1350));
  OAI211_X1 g1150(.A(new_n711), .B(new_n1245), .C1(new_n1350), .C2(KEYINPUT57), .ZN(new_n1351));
  AND3_X1   g1151(.A1(new_n1351), .A2(G378), .A3(new_n1230), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1276), .B1(new_n1351), .B2(new_n1230), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT124), .ZN(new_n1354));
  NOR3_X1   g1154(.A1(new_n1352), .A2(new_n1353), .A3(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(G375), .A2(new_n1309), .ZN(new_n1356));
  AOI21_X1  g1156(.A(KEYINPUT124), .B1(new_n1356), .B2(new_n1311), .ZN(new_n1357));
  OAI211_X1 g1157(.A(new_n1349), .B(new_n1321), .C1(new_n1355), .C2(new_n1357), .ZN(new_n1358));
  NOR3_X1   g1158(.A1(new_n1321), .A2(new_n1352), .A3(new_n1353), .ZN(new_n1359));
  INV_X1    g1159(.A(new_n1359), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1358), .A2(new_n1360), .ZN(new_n1361));
  OAI21_X1  g1161(.A(new_n1354), .B1(new_n1352), .B2(new_n1353), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1356), .A2(KEYINPUT124), .A3(new_n1311), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1362), .A2(new_n1363), .ZN(new_n1364));
  AOI21_X1  g1164(.A(new_n1349), .B1(new_n1364), .B2(new_n1321), .ZN(new_n1365));
  INV_X1    g1165(.A(KEYINPUT126), .ZN(new_n1366));
  AND3_X1   g1166(.A1(new_n1298), .A2(new_n1366), .A3(new_n1302), .ZN(new_n1367));
  AOI21_X1  g1167(.A(new_n1366), .B1(new_n1298), .B2(new_n1302), .ZN(new_n1368));
  OR2_X1    g1168(.A1(new_n1367), .A2(new_n1368), .ZN(new_n1369));
  NOR3_X1   g1169(.A1(new_n1361), .A2(new_n1365), .A3(new_n1369), .ZN(new_n1370));
  NOR2_X1   g1170(.A1(new_n1367), .A2(new_n1368), .ZN(new_n1371));
  AOI21_X1  g1171(.A(new_n1320), .B1(new_n1362), .B2(new_n1363), .ZN(new_n1372));
  AOI21_X1  g1172(.A(new_n1359), .B1(new_n1372), .B2(new_n1349), .ZN(new_n1373));
  OAI21_X1  g1173(.A(new_n1321), .B1(new_n1355), .B2(new_n1357), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1374), .A2(KEYINPUT125), .ZN(new_n1375));
  AOI21_X1  g1175(.A(new_n1371), .B1(new_n1373), .B2(new_n1375), .ZN(new_n1376));
  NOR2_X1   g1176(.A1(new_n1370), .A2(new_n1376), .ZN(G402));
endmodule


