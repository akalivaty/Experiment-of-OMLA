//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 1 0 1 1 1 0 0 0 1 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 0 0 1 0 0 0 1 0 1 0 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n803, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1016, new_n1017, new_n1018, new_n1019;
  INV_X1    g000(.A(KEYINPUT33), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(KEYINPUT32), .ZN(new_n203));
  INV_X1    g002(.A(G183gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT27), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT27), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G183gat), .ZN(new_n207));
  INV_X1    g006(.A(G190gat), .ZN(new_n208));
  AND4_X1   g007(.A1(KEYINPUT28), .A2(new_n205), .A3(new_n207), .A4(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT67), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n205), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT27), .B(G183gat), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n208), .B(new_n211), .C1(new_n212), .C2(new_n210), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT28), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n209), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT26), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NOR3_X1   g019(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n216), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT68), .B1(new_n215), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n222), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT68), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n205), .A2(new_n207), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT67), .ZN(new_n227));
  AOI21_X1  g026(.A(G190gat), .B1(new_n205), .B2(new_n210), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT28), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n224), .B(new_n225), .C1(new_n229), .C2(new_n209), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n218), .A2(KEYINPUT23), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT23), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(G169gat), .B2(G176gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n231), .A2(new_n217), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT64), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT24), .ZN(new_n236));
  AND3_X1   g035(.A1(new_n216), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n235), .B1(new_n216), .B2(new_n236), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n204), .A2(new_n208), .A3(KEYINPUT65), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT65), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(G183gat), .B2(G190gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n243));
  AND3_X1   g042(.A1(new_n240), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n234), .B1(new_n239), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n204), .A2(new_n208), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n236), .A2(KEYINPUT66), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n246), .A2(new_n247), .A3(new_n216), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n248), .B(KEYINPUT25), .C1(new_n216), .C2(new_n247), .ZN(new_n249));
  OAI22_X1  g048(.A1(new_n245), .A2(KEYINPUT25), .B1(new_n234), .B2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n223), .A2(new_n230), .A3(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G127gat), .B(G134gat), .ZN(new_n252));
  INV_X1    g051(.A(G113gat), .ZN(new_n253));
  INV_X1    g052(.A(G120gat), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT1), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n252), .B(new_n255), .C1(new_n253), .C2(new_n254), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n253), .A2(new_n254), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT1), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n258), .B1(G113gat), .B2(G120gat), .ZN(new_n259));
  INV_X1    g058(.A(G134gat), .ZN(new_n260));
  AND2_X1   g059(.A1(new_n260), .A2(G127gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(G127gat), .ZN(new_n262));
  OAI22_X1  g061(.A1(new_n257), .A2(new_n259), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n256), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n251), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT69), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n251), .A2(new_n267), .A3(new_n264), .ZN(new_n268));
  INV_X1    g067(.A(new_n264), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n223), .A2(new_n250), .A3(new_n230), .A4(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n266), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(G227gat), .A2(G233gat), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n203), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G15gat), .B(G43gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(G71gat), .B(G99gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n270), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n278), .B1(KEYINPUT69), .B2(new_n265), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n272), .B1(new_n279), .B2(new_n268), .ZN(new_n280));
  OAI21_X1  g079(.A(KEYINPUT32), .B1(new_n277), .B2(new_n202), .ZN(new_n281));
  OAI22_X1  g080(.A1(new_n274), .A2(new_n277), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n266), .A2(new_n272), .A3(new_n268), .A4(new_n270), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT34), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n279), .A2(KEYINPUT34), .A3(new_n272), .A4(new_n268), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(KEYINPUT71), .B1(new_n282), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n277), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n289), .B1(new_n280), .B2(new_n203), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n285), .A2(new_n286), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n271), .A2(new_n273), .ZN(new_n293));
  INV_X1    g092(.A(new_n281), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n290), .A2(new_n291), .A3(new_n292), .A4(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT70), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n291), .B1(new_n282), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n290), .A2(KEYINPUT70), .A3(new_n295), .ZN(new_n299));
  AOI22_X1  g098(.A1(new_n288), .A2(new_n296), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT30), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n224), .B1(new_n229), .B2(new_n209), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n250), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G226gat), .A2(G233gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n305), .B1(new_n251), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(G211gat), .A2(G218gat), .ZN(new_n308));
  INV_X1    g107(.A(G211gat), .ZN(new_n309));
  INV_X1    g108(.A(G218gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AND2_X1   g110(.A1(G197gat), .A2(G204gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(G197gat), .A2(G204gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT22), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n308), .B(new_n311), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n311), .A2(new_n308), .ZN(new_n317));
  XNOR2_X1  g116(.A(G197gat), .B(G204gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n308), .A2(new_n315), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  AND2_X1   g119(.A1(new_n316), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n322), .ZN(new_n323));
  OR2_X1    g122(.A1(new_n303), .A2(new_n306), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n251), .A2(new_n304), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n324), .A2(new_n321), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G8gat), .B(G36gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(G64gat), .ZN(new_n329));
  INV_X1    g128(.A(G92gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n329), .B(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n301), .B1(new_n327), .B2(new_n332), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n323), .A2(new_n326), .A3(KEYINPUT30), .A4(new_n331), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT72), .B1(new_n327), .B2(new_n332), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT72), .ZN(new_n336));
  AOI211_X1 g135(.A(new_n336), .B(new_n331), .C1(new_n323), .C2(new_n326), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n333), .B(new_n334), .C1(new_n335), .C2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT77), .ZN(new_n339));
  XOR2_X1   g138(.A(G141gat), .B(G148gat), .Z(new_n340));
  INV_X1    g139(.A(G155gat), .ZN(new_n341));
  INV_X1    g140(.A(G162gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(G155gat), .A2(G162gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(KEYINPUT2), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n340), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G141gat), .B(G148gat), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n344), .B(new_n343), .C1(new_n348), .C2(KEYINPUT2), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n350), .A2(new_n264), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT4), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n339), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n349), .A2(new_n347), .A3(new_n256), .A4(new_n263), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT4), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n354), .A2(new_n339), .A3(KEYINPUT4), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT3), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n347), .A2(new_n349), .A3(new_n359), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n360), .A2(new_n264), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT73), .B1(new_n350), .B2(KEYINPUT3), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT73), .ZN(new_n363));
  AOI211_X1 g162(.A(new_n363), .B(new_n359), .C1(new_n347), .C2(new_n349), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n361), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(G225gat), .A2(G233gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NOR3_X1   g166(.A1(new_n358), .A2(new_n367), .A3(KEYINPUT5), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT75), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n350), .A2(new_n264), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(new_n354), .ZN(new_n371));
  INV_X1    g170(.A(new_n366), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT74), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT74), .ZN(new_n374));
  AOI211_X1 g173(.A(new_n374), .B(new_n366), .C1(new_n370), .C2(new_n354), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT5), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n354), .B(KEYINPUT4), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n365), .A2(new_n377), .A3(new_n366), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n369), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT5), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n349), .A2(new_n347), .B1(new_n256), .B2(new_n263), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n372), .B1(new_n351), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n374), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n371), .A2(KEYINPUT74), .A3(new_n372), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n380), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n365), .A2(new_n377), .A3(new_n366), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n385), .A2(KEYINPUT75), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n368), .B1(new_n379), .B2(new_n387), .ZN(new_n388));
  XOR2_X1   g187(.A(KEYINPUT76), .B(KEYINPUT0), .Z(new_n389));
  XNOR2_X1  g188(.A(G1gat), .B(G29gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n389), .B(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(G57gat), .B(G85gat), .ZN(new_n392));
  XOR2_X1   g191(.A(new_n391), .B(new_n392), .Z(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT78), .B1(new_n388), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT6), .B1(new_n388), .B2(new_n394), .ZN(new_n396));
  OR3_X1    g195(.A1(new_n358), .A2(KEYINPUT5), .A3(new_n367), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n383), .A2(new_n384), .ZN(new_n398));
  AND4_X1   g197(.A1(KEYINPUT75), .A2(new_n398), .A3(KEYINPUT5), .A4(new_n386), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT75), .B1(new_n385), .B2(new_n386), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n397), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT78), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(new_n402), .A3(new_n393), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n395), .A2(new_n396), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n401), .A2(KEYINPUT6), .A3(new_n393), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n338), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT81), .ZN(new_n407));
  INV_X1    g206(.A(G228gat), .ZN(new_n408));
  INV_X1    g207(.A(G233gat), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT29), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n360), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(new_n321), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT3), .B1(new_n322), .B2(new_n411), .ZN(new_n414));
  INV_X1    g213(.A(new_n350), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n410), .B(new_n413), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n413), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT80), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n316), .A2(KEYINPUT79), .A3(new_n320), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT79), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n317), .A2(new_n318), .A3(new_n420), .A4(new_n319), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n411), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n418), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n316), .A2(KEYINPUT79), .A3(new_n320), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n424), .A2(KEYINPUT80), .A3(new_n411), .A4(new_n421), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n423), .A2(new_n359), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n417), .B1(new_n426), .B2(new_n350), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n416), .B1(new_n427), .B2(new_n410), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n407), .B1(new_n428), .B2(G22gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(G78gat), .B(G106gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(KEYINPUT31), .ZN(new_n431));
  INV_X1    g230(.A(G50gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(KEYINPUT82), .B1(new_n429), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT82), .ZN(new_n436));
  INV_X1    g235(.A(G22gat), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n424), .A2(new_n411), .A3(new_n421), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT3), .B1(new_n438), .B2(new_n418), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n415), .B1(new_n439), .B2(new_n425), .ZN(new_n440));
  OAI22_X1  g239(.A1(new_n440), .A2(new_n417), .B1(new_n408), .B2(new_n409), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n437), .B1(new_n441), .B2(new_n416), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n436), .B(new_n433), .C1(new_n442), .C2(new_n407), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n428), .B(new_n437), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n435), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n444), .B1(new_n435), .B2(new_n443), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n300), .A2(new_n406), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT35), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n288), .A2(new_n296), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n291), .B1(new_n290), .B2(new_n295), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT83), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n338), .A2(KEYINPUT35), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n435), .A2(new_n443), .ZN(new_n457));
  INV_X1    g256(.A(new_n444), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT6), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n460), .B1(new_n401), .B2(new_n393), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n388), .A2(new_n394), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n405), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AND4_X1   g262(.A1(new_n445), .A2(new_n456), .A3(new_n459), .A4(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT83), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n451), .A2(new_n465), .A3(new_n453), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n455), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT36), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n282), .A2(new_n297), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n470), .A2(new_n299), .A3(new_n287), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n469), .B1(new_n451), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n404), .A2(new_n405), .ZN(new_n474));
  INV_X1    g273(.A(new_n338), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n445), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n451), .A2(new_n469), .A3(new_n453), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n307), .A2(new_n321), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n324), .A2(new_n322), .A3(new_n325), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(KEYINPUT37), .A3(new_n481), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n482), .B(new_n332), .C1(new_n327), .C2(KEYINPUT37), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT38), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n323), .A2(new_n326), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT37), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n327), .A2(KEYINPUT37), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(KEYINPUT38), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n401), .A2(new_n393), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n396), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n331), .B1(new_n486), .B2(KEYINPUT38), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n491), .A2(new_n493), .A3(new_n405), .A4(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n356), .A2(new_n365), .A3(new_n357), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT39), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(new_n497), .A3(new_n372), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n496), .A2(new_n372), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT39), .B1(new_n371), .B2(new_n372), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n394), .B(new_n498), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT40), .ZN(new_n502));
  OR2_X1    g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n501), .A2(new_n502), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n338), .A2(new_n503), .A3(new_n492), .A4(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n448), .A2(new_n495), .A3(new_n505), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n473), .A2(new_n478), .A3(new_n479), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n468), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(G15gat), .B(G22gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT87), .ZN(new_n510));
  INV_X1    g309(.A(G1gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT16), .ZN(new_n512));
  AOI22_X1  g311(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n509), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n509), .A2(KEYINPUT87), .A3(G1gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(G8gat), .ZN(new_n516));
  INV_X1    g315(.A(G8gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n513), .A2(new_n517), .A3(new_n514), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT17), .ZN(new_n520));
  INV_X1    g319(.A(G29gat), .ZN(new_n521));
  INV_X1    g320(.A(G36gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT14), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT14), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n524), .B1(G29gat), .B2(G36gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(G29gat), .A2(G36gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G43gat), .B(G50gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(KEYINPUT15), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT85), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT85), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n527), .A2(new_n532), .A3(KEYINPUT15), .A4(new_n529), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n528), .A2(new_n530), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT86), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n536), .B1(new_n529), .B2(KEYINPUT15), .ZN(new_n537));
  OR3_X1    g336(.A1(new_n529), .A2(new_n536), .A3(KEYINPUT15), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n520), .B1(new_n534), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n537), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n541), .A2(new_n530), .A3(new_n528), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n531), .A2(new_n533), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n542), .A2(KEYINPUT17), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n519), .A2(new_n540), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n516), .A2(new_n518), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n542), .A2(new_n543), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(G229gat), .A2(G233gat), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT88), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT18), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT18), .ZN(new_n554));
  OAI211_X1 g353(.A(KEYINPUT88), .B(new_n554), .C1(new_n549), .C2(new_n551), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n546), .B(new_n547), .ZN(new_n556));
  XOR2_X1   g355(.A(new_n550), .B(KEYINPUT13), .Z(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G169gat), .B(G197gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(G113gat), .B(G141gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(KEYINPUT12), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n553), .A2(new_n555), .A3(new_n558), .A4(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT89), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n552), .A2(KEYINPUT18), .B1(new_n556), .B2(new_n557), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT89), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n567), .A2(new_n568), .A3(new_n555), .A4(new_n564), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n567), .A2(new_n555), .ZN(new_n571));
  INV_X1    g370(.A(new_n564), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G190gat), .B(G218gat), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT41), .ZN(new_n577));
  INV_X1    g376(.A(G232gat), .ZN(new_n578));
  NOR3_X1   g377(.A1(new_n577), .A2(new_n578), .A3(new_n409), .ZN(new_n579));
  NAND2_X1  g378(.A1(G85gat), .A2(G92gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT7), .ZN(new_n581));
  XNOR2_X1  g380(.A(G99gat), .B(G106gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(G99gat), .A2(G106gat), .ZN(new_n583));
  INV_X1    g382(.A(G85gat), .ZN(new_n584));
  AOI22_X1  g383(.A1(KEYINPUT8), .A2(new_n583), .B1(new_n584), .B2(new_n330), .ZN(new_n585));
  AND3_X1   g384(.A1(new_n581), .A2(new_n582), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n582), .B1(new_n581), .B2(new_n585), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n579), .B1(new_n547), .B2(new_n588), .ZN(new_n589));
  OR2_X1    g388(.A1(new_n588), .A2(KEYINPUT93), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(KEYINPUT93), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n540), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n544), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n576), .B(new_n589), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(KEYINPUT94), .ZN(new_n595));
  XNOR2_X1  g394(.A(KEYINPUT92), .B(G134gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(G162gat), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n577), .B1(new_n578), .B2(new_n409), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n589), .B1(new_n592), .B2(new_n593), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(new_n575), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(new_n594), .ZN(new_n603));
  OR2_X1    g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(G64gat), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n605), .A2(G57gat), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n605), .A2(G57gat), .ZN(new_n607));
  INV_X1    g406(.A(G71gat), .ZN(new_n608));
  INV_X1    g407(.A(G78gat), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI22_X1  g409(.A1(new_n606), .A2(new_n607), .B1(new_n610), .B2(KEYINPUT9), .ZN(new_n611));
  XOR2_X1   g410(.A(G71gat), .B(G78gat), .Z(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT21), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g414(.A(KEYINPUT91), .B1(new_n546), .B2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT91), .ZN(new_n617));
  INV_X1    g416(.A(new_n615), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n519), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n613), .A2(new_n614), .ZN(new_n620));
  INV_X1    g419(.A(G231gat), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n621), .A2(new_n409), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G127gat), .B(G155gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT20), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  OAI211_X1 g425(.A(new_n613), .B(new_n614), .C1(new_n621), .C2(new_n409), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n623), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n626), .B1(new_n623), .B2(new_n627), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n616), .B(new_n619), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n619), .A2(new_n616), .ZN(new_n632));
  INV_X1    g431(.A(new_n630), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n632), .A2(new_n633), .A3(new_n628), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G183gat), .B(G211gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n631), .A2(new_n634), .A3(new_n638), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n613), .B1(new_n586), .B2(new_n587), .ZN(new_n643));
  INV_X1    g442(.A(new_n612), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n611), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(new_n588), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(G230gat), .A2(G233gat), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n648), .B(KEYINPUT95), .Z(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT96), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT10), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n643), .A2(new_n653), .A3(new_n646), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n645), .A2(new_n588), .A3(KEYINPUT10), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n649), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(G120gat), .B(G148gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(G176gat), .ZN(new_n660));
  INV_X1    g459(.A(G204gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n652), .A2(new_n658), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n662), .ZN(new_n664));
  INV_X1    g463(.A(new_n650), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n649), .B1(new_n654), .B2(new_n655), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n600), .A2(new_n603), .ZN(new_n669));
  AND4_X1   g468(.A1(new_n604), .A2(new_n642), .A3(new_n668), .A4(new_n669), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n574), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n508), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n672), .A2(new_n474), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(new_n511), .ZN(G1324gat));
  XOR2_X1   g473(.A(KEYINPUT16), .B(G8gat), .Z(new_n675));
  NAND4_X1  g474(.A1(new_n508), .A2(new_n338), .A3(new_n671), .A4(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT42), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT97), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n676), .A2(new_n677), .ZN(new_n681));
  OAI21_X1  g480(.A(G8gat), .B1(new_n672), .B2(new_n475), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT98), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n680), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT99), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1325gat));
  AOI211_X1 g485(.A(KEYINPUT36), .B(new_n452), .C1(new_n288), .C2(new_n296), .ZN(new_n687));
  OAI21_X1  g486(.A(KEYINPUT100), .B1(new_n472), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT100), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n479), .B(new_n689), .C1(new_n300), .C2(new_n469), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT101), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(G15gat), .B1(new_n693), .B2(new_n672), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n465), .B1(new_n451), .B2(new_n453), .ZN(new_n695));
  AOI211_X1 g494(.A(KEYINPUT83), .B(new_n452), .C1(new_n288), .C2(new_n296), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n698), .A2(G15gat), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n694), .B1(new_n672), .B2(new_n699), .ZN(G1326gat));
  NOR2_X1   g499(.A1(new_n672), .A2(new_n448), .ZN(new_n701));
  XOR2_X1   g500(.A(KEYINPUT43), .B(G22gat), .Z(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1327gat));
  NAND2_X1  g502(.A1(new_n604), .A2(new_n669), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n508), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n574), .ZN(new_n706));
  INV_X1    g505(.A(new_n668), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n706), .A2(new_n642), .A3(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n474), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(new_n521), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT45), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n505), .A2(new_n445), .A3(new_n459), .ZN(new_n714));
  OAI211_X1 g513(.A(new_n405), .B(new_n494), .C1(new_n461), .C2(new_n462), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n485), .A2(new_n490), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OAI22_X1  g516(.A1(new_n714), .A2(new_n717), .B1(new_n448), .B2(new_n406), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n691), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT102), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n720), .A2(new_n721), .A3(new_n468), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n718), .B1(new_n688), .B2(new_n690), .ZN(new_n723));
  AOI22_X1  g522(.A1(new_n697), .A2(new_n464), .B1(new_n449), .B2(KEYINPUT35), .ZN(new_n724));
  OAI21_X1  g523(.A(KEYINPUT102), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n704), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n726), .A2(KEYINPUT44), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n722), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n705), .A2(KEYINPUT44), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n708), .ZN(new_n731));
  OAI21_X1  g530(.A(G29gat), .B1(new_n731), .B2(new_n474), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n713), .A2(new_n732), .ZN(G1328gat));
  NAND3_X1  g532(.A1(new_n710), .A2(new_n522), .A3(new_n338), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n734), .B(KEYINPUT46), .Z(new_n735));
  OAI21_X1  g534(.A(G36gat), .B1(new_n731), .B2(new_n475), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(G1329gat));
  NOR2_X1   g536(.A1(new_n698), .A2(G43gat), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n508), .A2(new_n704), .A3(new_n708), .A4(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(KEYINPUT103), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n726), .B1(new_n468), .B2(new_n507), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT103), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n741), .A2(new_n742), .A3(new_n708), .A4(new_n738), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT47), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  AOI211_X1 g543(.A(new_n693), .B(new_n709), .C1(new_n728), .C2(new_n729), .ZN(new_n745));
  INV_X1    g544(.A(G43gat), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n744), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT104), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n740), .A2(new_n743), .ZN(new_n749));
  INV_X1    g548(.A(new_n691), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n730), .A2(new_n750), .A3(new_n708), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n749), .B1(new_n751), .B2(G43gat), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT47), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n747), .B(new_n748), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n709), .B1(new_n728), .B2(new_n729), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n746), .B1(new_n756), .B2(new_n750), .ZN(new_n757));
  OAI21_X1  g556(.A(KEYINPUT47), .B1(new_n757), .B2(new_n749), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n748), .B1(new_n758), .B2(new_n747), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n755), .A2(new_n759), .ZN(G1330gat));
  INV_X1    g559(.A(KEYINPUT48), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT105), .ZN(new_n762));
  OAI21_X1  g561(.A(G50gat), .B1(new_n731), .B2(new_n448), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n710), .A2(new_n432), .A3(new_n477), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n432), .B1(new_n756), .B2(new_n477), .ZN(new_n766));
  INV_X1    g565(.A(new_n764), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n766), .A2(KEYINPUT105), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n761), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n763), .A2(new_n762), .A3(new_n764), .ZN(new_n770));
  OAI21_X1  g569(.A(KEYINPUT105), .B1(new_n766), .B2(new_n767), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n770), .A2(KEYINPUT48), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n769), .A2(new_n772), .ZN(G1331gat));
  INV_X1    g572(.A(new_n642), .ZN(new_n774));
  NOR4_X1   g573(.A1(new_n574), .A2(new_n704), .A3(new_n774), .A4(new_n668), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n722), .A2(new_n725), .A3(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT106), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n722), .A2(new_n725), .A3(KEYINPUT106), .A4(new_n775), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n778), .A2(new_n711), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(G57gat), .ZN(G1332gat));
  INV_X1    g580(.A(KEYINPUT49), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n475), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n778), .A2(new_n779), .A3(new_n783), .ZN(new_n784));
  OR2_X1    g583(.A1(new_n784), .A2(KEYINPUT107), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(KEYINPUT107), .ZN(new_n786));
  AND4_X1   g585(.A1(new_n782), .A2(new_n785), .A3(new_n605), .A4(new_n786), .ZN(new_n787));
  AOI22_X1  g586(.A1(new_n785), .A2(new_n786), .B1(new_n782), .B2(new_n605), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n787), .A2(new_n788), .ZN(G1333gat));
  NOR2_X1   g588(.A1(new_n693), .A2(new_n608), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n778), .A2(new_n779), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT108), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n778), .A2(KEYINPUT108), .A3(new_n779), .A4(new_n790), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n778), .A2(new_n697), .A3(new_n779), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n608), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT50), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT50), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n795), .A2(new_n800), .A3(new_n797), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(G1334gat));
  NAND3_X1  g601(.A1(new_n778), .A2(new_n477), .A3(new_n779), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g603(.A1(new_n574), .A2(new_n642), .A3(new_n668), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n730), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(G85gat), .B1(new_n806), .B2(new_n474), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT51), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n720), .A2(new_n468), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n809), .A2(KEYINPUT109), .A3(new_n704), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n574), .A2(new_n642), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT109), .B1(new_n809), .B2(new_n704), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n808), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n809), .A2(new_n704), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT109), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n817), .A2(KEYINPUT51), .A3(new_n810), .A4(new_n811), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n707), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n711), .A2(new_n584), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n807), .B1(new_n820), .B2(new_n821), .ZN(G1336gat));
  NOR2_X1   g621(.A1(new_n475), .A2(G92gat), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n819), .A2(new_n707), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(G92gat), .B1(new_n806), .B2(new_n475), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g625(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n824), .A2(new_n827), .A3(new_n825), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(G1337gat));
  OAI21_X1  g630(.A(G99gat), .B1(new_n806), .B2(new_n693), .ZN(new_n832));
  INV_X1    g631(.A(new_n819), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n698), .A2(G99gat), .A3(new_n668), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(KEYINPUT111), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n832), .B1(new_n833), .B2(new_n835), .ZN(G1338gat));
  OAI21_X1  g635(.A(G106gat), .B1(new_n806), .B2(new_n448), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  OR3_X1    g637(.A1(new_n448), .A2(G106gat), .A3(new_n668), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT112), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n840), .B1(new_n814), .B2(new_n818), .ZN(new_n841));
  OAI21_X1  g640(.A(KEYINPUT53), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT53), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n837), .B(new_n843), .C1(new_n833), .C2(new_n839), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n844), .ZN(G1339gat));
  NAND3_X1  g644(.A1(new_n654), .A2(new_n649), .A3(new_n655), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n658), .A2(KEYINPUT54), .A3(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n662), .B1(new_n666), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n847), .A2(KEYINPUT55), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n663), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT55), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n847), .A2(new_n849), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n854), .A2(new_n704), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n549), .A2(new_n551), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n856), .B1(new_n556), .B2(new_n557), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n857), .A2(new_n563), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n858), .B1(new_n566), .B2(new_n569), .ZN(new_n859));
  AOI21_X1  g658(.A(KEYINPUT113), .B1(new_n855), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n855), .A2(KEYINPUT113), .A3(new_n859), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n574), .A2(new_n854), .ZN(new_n864));
  AOI211_X1 g663(.A(new_n668), .B(new_n858), .C1(new_n566), .C2(new_n569), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n726), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n642), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n670), .A2(new_n573), .A3(new_n570), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n448), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT114), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI211_X1 g671(.A(KEYINPUT114), .B(new_n448), .C1(new_n867), .C2(new_n869), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n474), .A2(new_n338), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n872), .A2(new_n873), .A3(new_n697), .A4(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT115), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n698), .B1(new_n870), .B2(new_n871), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n878), .A2(KEYINPUT115), .A3(new_n874), .A4(new_n873), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n877), .A2(new_n879), .A3(G113gat), .A4(new_n574), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n863), .A2(new_n866), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n869), .B1(new_n881), .B2(new_n774), .ZN(new_n882));
  INV_X1    g681(.A(new_n874), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n300), .A2(new_n448), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n253), .B1(new_n887), .B2(new_n706), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n880), .A2(new_n888), .ZN(G1340gat));
  NAND3_X1  g688(.A1(new_n877), .A2(new_n879), .A3(new_n707), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT116), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n890), .A2(new_n891), .A3(G120gat), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n891), .B1(new_n890), .B2(G120gat), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n707), .A2(new_n254), .ZN(new_n894));
  OAI22_X1  g693(.A1(new_n892), .A2(new_n893), .B1(new_n887), .B2(new_n894), .ZN(G1341gat));
  NAND3_X1  g694(.A1(new_n877), .A2(new_n879), .A3(new_n642), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(G127gat), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n774), .A2(G127gat), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n897), .B1(new_n887), .B2(new_n898), .ZN(G1342gat));
  NAND2_X1  g698(.A1(new_n704), .A2(new_n260), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT56), .B1(new_n887), .B2(new_n900), .ZN(new_n901));
  OR3_X1    g700(.A1(new_n887), .A2(KEYINPUT56), .A3(new_n900), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n877), .A2(new_n879), .A3(new_n704), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n901), .B(new_n902), .C1(new_n903), .C2(new_n260), .ZN(G1343gat));
  NAND3_X1  g703(.A1(new_n884), .A2(new_n477), .A3(new_n693), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(G141gat), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n906), .A2(new_n907), .A3(new_n574), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n750), .A2(new_n883), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT57), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n911), .B1(new_n882), .B2(new_n448), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n448), .A2(new_n911), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n853), .A2(KEYINPUT117), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT117), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n847), .A2(new_n915), .A3(new_n849), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n914), .A2(new_n852), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n917), .A2(new_n663), .A3(new_n850), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n918), .B1(new_n570), .B2(new_n573), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n726), .B1(new_n919), .B2(new_n865), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n642), .B1(new_n863), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n913), .B1(new_n921), .B2(new_n869), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n910), .B1(new_n912), .B2(new_n922), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n923), .A2(new_n574), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n908), .B1(new_n924), .B2(new_n907), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT58), .ZN(G1344gat));
  NAND2_X1  g725(.A1(new_n923), .A2(new_n707), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT59), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n927), .A2(new_n928), .A3(G148gat), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n750), .A2(KEYINPUT118), .A3(new_n883), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT118), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n931), .B1(new_n691), .B2(new_n874), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n868), .A2(KEYINPUT119), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT119), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n670), .A2(new_n935), .A3(new_n573), .A4(new_n570), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n855), .A2(new_n859), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n920), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n937), .B1(new_n939), .B2(new_n774), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n448), .B1(new_n940), .B2(KEYINPUT120), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT120), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n642), .B1(new_n920), .B2(new_n938), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n942), .B1(new_n943), .B2(new_n937), .ZN(new_n944));
  AOI21_X1  g743(.A(KEYINPUT57), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(new_n913), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n882), .A2(new_n946), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n707), .B(new_n933), .C1(new_n945), .C2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(G148gat), .ZN(new_n949));
  AOI21_X1  g748(.A(KEYINPUT121), .B1(new_n949), .B2(KEYINPUT59), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT121), .ZN(new_n951));
  AOI211_X1 g750(.A(new_n951), .B(new_n928), .C1(new_n948), .C2(G148gat), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n929), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  OR3_X1    g752(.A1(new_n905), .A2(G148gat), .A3(new_n668), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(G1345gat));
  NAND3_X1  g754(.A1(new_n906), .A2(new_n341), .A3(new_n642), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n923), .A2(new_n642), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n956), .B1(new_n957), .B2(new_n341), .ZN(G1346gat));
  NAND3_X1  g757(.A1(new_n906), .A2(new_n342), .A3(new_n704), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n923), .A2(new_n704), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n959), .B1(new_n960), .B2(new_n342), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT122), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n961), .B(new_n962), .ZN(G1347gat));
  NOR4_X1   g762(.A1(new_n882), .A2(new_n711), .A3(new_n475), .A4(new_n885), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(new_n574), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n711), .A2(new_n475), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n878), .A2(new_n873), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n574), .A2(G169gat), .ZN(new_n969));
  OAI22_X1  g768(.A1(new_n966), .A2(G169gat), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  XNOR2_X1  g769(.A(new_n970), .B(KEYINPUT123), .ZN(G1348gat));
  OAI21_X1  g770(.A(G176gat), .B1(new_n968), .B2(new_n668), .ZN(new_n972));
  INV_X1    g771(.A(G176gat), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n964), .A2(new_n973), .A3(new_n707), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n972), .A2(new_n974), .ZN(G1349gat));
  OAI21_X1  g774(.A(G183gat), .B1(new_n968), .B2(new_n774), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n774), .A2(new_n226), .ZN(new_n977));
  AOI21_X1  g776(.A(KEYINPUT124), .B1(new_n964), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g778(.A(new_n979), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g779(.A(KEYINPUT125), .ZN(new_n981));
  NAND4_X1  g780(.A1(new_n878), .A2(new_n704), .A3(new_n873), .A4(new_n967), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n981), .B1(new_n982), .B2(G190gat), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT61), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n982), .A2(new_n981), .A3(G190gat), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n964), .A2(new_n208), .A3(new_n704), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n983), .A2(new_n984), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(G1351gat));
  NAND2_X1  g789(.A1(new_n693), .A2(new_n967), .ZN(new_n991));
  INV_X1    g790(.A(new_n991), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n882), .A2(new_n448), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g793(.A(new_n994), .ZN(new_n995));
  INV_X1    g794(.A(G197gat), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n995), .A2(new_n996), .A3(new_n574), .ZN(new_n997));
  NOR2_X1   g796(.A1(new_n945), .A2(new_n947), .ZN(new_n998));
  NOR3_X1   g797(.A1(new_n998), .A2(new_n706), .A3(new_n991), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n997), .B1(new_n999), .B2(new_n996), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n1000), .A2(KEYINPUT126), .ZN(new_n1001));
  INV_X1    g800(.A(KEYINPUT126), .ZN(new_n1002));
  OAI211_X1 g801(.A(new_n997), .B(new_n1002), .C1(new_n999), .C2(new_n996), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1001), .A2(new_n1003), .ZN(G1352gat));
  NAND2_X1  g803(.A1(new_n707), .A2(new_n661), .ZN(new_n1005));
  OR3_X1    g804(.A1(new_n994), .A2(KEYINPUT62), .A3(new_n1005), .ZN(new_n1006));
  OAI21_X1  g805(.A(KEYINPUT62), .B1(new_n994), .B2(new_n1005), .ZN(new_n1007));
  NOR3_X1   g806(.A1(new_n998), .A2(new_n668), .A3(new_n991), .ZN(new_n1008));
  OAI211_X1 g807(.A(new_n1006), .B(new_n1007), .C1(new_n661), .C2(new_n1008), .ZN(G1353gat));
  NAND3_X1  g808(.A1(new_n995), .A2(new_n309), .A3(new_n642), .ZN(new_n1010));
  NOR2_X1   g809(.A1(new_n998), .A2(new_n991), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1011), .A2(new_n642), .ZN(new_n1012));
  AND3_X1   g811(.A1(new_n1012), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1013));
  AOI21_X1  g812(.A(KEYINPUT63), .B1(new_n1012), .B2(G211gat), .ZN(new_n1014));
  OAI21_X1  g813(.A(new_n1010), .B1(new_n1013), .B2(new_n1014), .ZN(G1354gat));
  AOI21_X1  g814(.A(G218gat), .B1(new_n995), .B2(new_n704), .ZN(new_n1016));
  OR2_X1    g815(.A1(new_n1016), .A2(KEYINPUT127), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n1016), .A2(KEYINPUT127), .ZN(new_n1018));
  NOR2_X1   g817(.A1(new_n726), .A2(new_n310), .ZN(new_n1019));
  AOI22_X1  g818(.A1(new_n1017), .A2(new_n1018), .B1(new_n1011), .B2(new_n1019), .ZN(G1355gat));
endmodule


