

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U548 ( .A1(n542), .A2(n541), .ZN(G160) );
  OR2_X4 U549 ( .A1(n678), .A2(n677), .ZN(n723) );
  NOR2_X1 U550 ( .A1(n721), .A2(n720), .ZN(n722) );
  INV_X1 U551 ( .A(KEYINPUT99), .ZN(n747) );
  NOR2_X1 U552 ( .A1(n746), .A2(KEYINPUT33), .ZN(n748) );
  XNOR2_X1 U553 ( .A(KEYINPUT101), .B(n786), .ZN(n511) );
  XNOR2_X1 U554 ( .A(KEYINPUT93), .B(KEYINPUT26), .ZN(n679) );
  XNOR2_X1 U555 ( .A(n680), .B(n679), .ZN(n681) );
  INV_X1 U556 ( .A(KEYINPUT94), .ZN(n684) );
  NAND2_X1 U557 ( .A1(n787), .A2(n511), .ZN(n788) );
  NOR2_X1 U558 ( .A1(G2105), .A2(G2104), .ZN(n538) );
  XOR2_X1 U559 ( .A(G543), .B(KEYINPUT0), .Z(n646) );
  INV_X1 U560 ( .A(G651), .ZN(n519) );
  NOR2_X1 U561 ( .A1(n646), .A2(n519), .ZN(n635) );
  NAND2_X1 U562 ( .A1(G76), .A2(n635), .ZN(n516) );
  XOR2_X1 U563 ( .A(KEYINPUT4), .B(KEYINPUT73), .Z(n513) );
  NOR2_X1 U564 ( .A1(G543), .A2(G651), .ZN(n632) );
  NAND2_X1 U565 ( .A1(G89), .A2(n632), .ZN(n512) );
  XNOR2_X1 U566 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U567 ( .A(KEYINPUT72), .B(n514), .ZN(n515) );
  NAND2_X1 U568 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U569 ( .A(n517), .B(KEYINPUT74), .ZN(n518) );
  XNOR2_X1 U570 ( .A(KEYINPUT5), .B(n518), .ZN(n527) );
  XNOR2_X1 U571 ( .A(KEYINPUT75), .B(KEYINPUT6), .ZN(n525) );
  NOR2_X1 U572 ( .A1(G543), .A2(n519), .ZN(n521) );
  XNOR2_X1 U573 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n520) );
  XNOR2_X1 U574 ( .A(n521), .B(n520), .ZN(n645) );
  NAND2_X1 U575 ( .A1(G63), .A2(n645), .ZN(n523) );
  NOR2_X2 U576 ( .A1(n646), .A2(G651), .ZN(n641) );
  NAND2_X1 U577 ( .A1(G51), .A2(n641), .ZN(n522) );
  NAND2_X1 U578 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U579 ( .A(n525), .B(n524), .ZN(n526) );
  NAND2_X1 U580 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U581 ( .A(n528), .B(KEYINPUT76), .ZN(n529) );
  XNOR2_X1 U582 ( .A(KEYINPUT7), .B(n529), .ZN(G168) );
  XNOR2_X1 U583 ( .A(KEYINPUT77), .B(KEYINPUT8), .ZN(n530) );
  XNOR2_X1 U584 ( .A(n530), .B(G168), .ZN(G286) );
  XOR2_X1 U585 ( .A(KEYINPUT66), .B(KEYINPUT23), .Z(n533) );
  INV_X1 U586 ( .A(G2105), .ZN(n545) );
  AND2_X1 U587 ( .A1(n545), .A2(G101), .ZN(n531) );
  NAND2_X1 U588 ( .A1(G2104), .A2(n531), .ZN(n532) );
  XNOR2_X1 U589 ( .A(n533), .B(n532), .ZN(n537) );
  INV_X1 U590 ( .A(G2104), .ZN(n534) );
  AND2_X4 U591 ( .A1(n534), .A2(G2105), .ZN(n882) );
  NAND2_X1 U592 ( .A1(G125), .A2(n882), .ZN(n535) );
  XOR2_X1 U593 ( .A(KEYINPUT65), .B(n535), .Z(n536) );
  NAND2_X1 U594 ( .A1(n537), .A2(n536), .ZN(n542) );
  XOR2_X1 U595 ( .A(KEYINPUT17), .B(n538), .Z(n601) );
  NAND2_X1 U596 ( .A1(G137), .A2(n601), .ZN(n540) );
  AND2_X1 U597 ( .A1(G2105), .A2(G2104), .ZN(n883) );
  NAND2_X1 U598 ( .A1(G113), .A2(n883), .ZN(n539) );
  NAND2_X1 U599 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U600 ( .A1(G126), .A2(n882), .ZN(n544) );
  NAND2_X1 U601 ( .A1(G138), .A2(n601), .ZN(n543) );
  NAND2_X1 U602 ( .A1(n544), .A2(n543), .ZN(n549) );
  NAND2_X1 U603 ( .A1(G114), .A2(n883), .ZN(n547) );
  AND2_X1 U604 ( .A1(n545), .A2(G2104), .ZN(n887) );
  NAND2_X1 U605 ( .A1(G102), .A2(n887), .ZN(n546) );
  NAND2_X1 U606 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U607 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U608 ( .A(KEYINPUT85), .B(n550), .Z(n677) );
  BUF_X1 U609 ( .A(n677), .Z(G164) );
  AND2_X1 U610 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U611 ( .A(G132), .ZN(G219) );
  INV_X1 U612 ( .A(G82), .ZN(G220) );
  INV_X1 U613 ( .A(G57), .ZN(G237) );
  INV_X1 U614 ( .A(G120), .ZN(G236) );
  INV_X1 U615 ( .A(G108), .ZN(G238) );
  NAND2_X1 U616 ( .A1(G64), .A2(n645), .ZN(n552) );
  NAND2_X1 U617 ( .A1(G52), .A2(n641), .ZN(n551) );
  NAND2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n557) );
  NAND2_X1 U619 ( .A1(G90), .A2(n632), .ZN(n554) );
  NAND2_X1 U620 ( .A1(G77), .A2(n635), .ZN(n553) );
  NAND2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U622 ( .A(KEYINPUT9), .B(n555), .Z(n556) );
  NOR2_X1 U623 ( .A1(n557), .A2(n556), .ZN(G171) );
  NAND2_X1 U624 ( .A1(G7), .A2(G661), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n558), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U626 ( .A(KEYINPUT11), .B(KEYINPUT68), .Z(n560) );
  INV_X1 U627 ( .A(G223), .ZN(n834) );
  NAND2_X1 U628 ( .A1(G567), .A2(n834), .ZN(n559) );
  XNOR2_X1 U629 ( .A(n560), .B(n559), .ZN(G234) );
  NAND2_X1 U630 ( .A1(n645), .A2(G56), .ZN(n561) );
  XNOR2_X1 U631 ( .A(KEYINPUT14), .B(n561), .ZN(n567) );
  NAND2_X1 U632 ( .A1(n632), .A2(G81), .ZN(n562) );
  XNOR2_X1 U633 ( .A(n562), .B(KEYINPUT12), .ZN(n564) );
  NAND2_X1 U634 ( .A1(G68), .A2(n635), .ZN(n563) );
  NAND2_X1 U635 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U636 ( .A(KEYINPUT13), .B(n565), .ZN(n566) );
  NAND2_X1 U637 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U638 ( .A(n568), .B(KEYINPUT69), .ZN(n570) );
  NAND2_X1 U639 ( .A1(n641), .A2(G43), .ZN(n569) );
  NAND2_X1 U640 ( .A1(n570), .A2(n569), .ZN(n970) );
  INV_X1 U641 ( .A(n970), .ZN(n571) );
  XNOR2_X1 U642 ( .A(G860), .B(KEYINPUT70), .ZN(n590) );
  NAND2_X1 U643 ( .A1(n571), .A2(n590), .ZN(G153) );
  INV_X1 U644 ( .A(G171), .ZN(G301) );
  NAND2_X1 U645 ( .A1(G868), .A2(G301), .ZN(n581) );
  NAND2_X1 U646 ( .A1(n635), .A2(G79), .ZN(n578) );
  NAND2_X1 U647 ( .A1(G66), .A2(n645), .ZN(n573) );
  NAND2_X1 U648 ( .A1(G92), .A2(n632), .ZN(n572) );
  NAND2_X1 U649 ( .A1(n573), .A2(n572), .ZN(n576) );
  NAND2_X1 U650 ( .A1(G54), .A2(n641), .ZN(n574) );
  XNOR2_X1 U651 ( .A(KEYINPUT71), .B(n574), .ZN(n575) );
  NOR2_X1 U652 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U653 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U654 ( .A(KEYINPUT15), .B(n579), .Z(n965) );
  INV_X1 U655 ( .A(G868), .ZN(n657) );
  NAND2_X1 U656 ( .A1(n965), .A2(n657), .ZN(n580) );
  NAND2_X1 U657 ( .A1(n581), .A2(n580), .ZN(G284) );
  NAND2_X1 U658 ( .A1(G65), .A2(n645), .ZN(n583) );
  NAND2_X1 U659 ( .A1(G53), .A2(n641), .ZN(n582) );
  NAND2_X1 U660 ( .A1(n583), .A2(n582), .ZN(n587) );
  NAND2_X1 U661 ( .A1(G91), .A2(n632), .ZN(n585) );
  NAND2_X1 U662 ( .A1(G78), .A2(n635), .ZN(n584) );
  NAND2_X1 U663 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U664 ( .A1(n587), .A2(n586), .ZN(n973) );
  INV_X1 U665 ( .A(n973), .ZN(G299) );
  NAND2_X1 U666 ( .A1(G868), .A2(G286), .ZN(n589) );
  NAND2_X1 U667 ( .A1(G299), .A2(n657), .ZN(n588) );
  NAND2_X1 U668 ( .A1(n589), .A2(n588), .ZN(G297) );
  INV_X1 U669 ( .A(G559), .ZN(n591) );
  NOR2_X1 U670 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U671 ( .A1(n965), .A2(n592), .ZN(n593) );
  XOR2_X1 U672 ( .A(KEYINPUT16), .B(n593), .Z(G148) );
  NOR2_X1 U673 ( .A1(G868), .A2(n970), .ZN(n596) );
  INV_X1 U674 ( .A(n965), .ZN(n616) );
  NAND2_X1 U675 ( .A1(G868), .A2(n616), .ZN(n594) );
  NOR2_X1 U676 ( .A1(G559), .A2(n594), .ZN(n595) );
  NOR2_X1 U677 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U678 ( .A(KEYINPUT78), .B(n597), .ZN(G282) );
  NAND2_X1 U679 ( .A1(n882), .A2(G123), .ZN(n598) );
  XNOR2_X1 U680 ( .A(n598), .B(KEYINPUT18), .ZN(n600) );
  NAND2_X1 U681 ( .A1(G111), .A2(n883), .ZN(n599) );
  NAND2_X1 U682 ( .A1(n600), .A2(n599), .ZN(n605) );
  BUF_X1 U683 ( .A(n601), .Z(n886) );
  NAND2_X1 U684 ( .A1(G135), .A2(n886), .ZN(n603) );
  NAND2_X1 U685 ( .A1(G99), .A2(n887), .ZN(n602) );
  NAND2_X1 U686 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U687 ( .A1(n605), .A2(n604), .ZN(n915) );
  XNOR2_X1 U688 ( .A(n915), .B(G2096), .ZN(n607) );
  INV_X1 U689 ( .A(G2100), .ZN(n606) );
  NAND2_X1 U690 ( .A1(n607), .A2(n606), .ZN(G156) );
  NAND2_X1 U691 ( .A1(G55), .A2(n641), .ZN(n608) );
  XNOR2_X1 U692 ( .A(n608), .B(KEYINPUT80), .ZN(n615) );
  NAND2_X1 U693 ( .A1(G93), .A2(n632), .ZN(n610) );
  NAND2_X1 U694 ( .A1(G80), .A2(n635), .ZN(n609) );
  NAND2_X1 U695 ( .A1(n610), .A2(n609), .ZN(n613) );
  NAND2_X1 U696 ( .A1(G67), .A2(n645), .ZN(n611) );
  XNOR2_X1 U697 ( .A(KEYINPUT79), .B(n611), .ZN(n612) );
  NOR2_X1 U698 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U699 ( .A1(n615), .A2(n614), .ZN(n658) );
  NAND2_X1 U700 ( .A1(G559), .A2(n616), .ZN(n617) );
  XNOR2_X1 U701 ( .A(n970), .B(n617), .ZN(n655) );
  NOR2_X1 U702 ( .A1(G860), .A2(n655), .ZN(n618) );
  XOR2_X1 U703 ( .A(n658), .B(n618), .Z(G145) );
  NAND2_X1 U704 ( .A1(n635), .A2(G75), .ZN(n621) );
  NAND2_X1 U705 ( .A1(G88), .A2(n632), .ZN(n619) );
  XOR2_X1 U706 ( .A(KEYINPUT81), .B(n619), .Z(n620) );
  NAND2_X1 U707 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U708 ( .A1(G62), .A2(n645), .ZN(n623) );
  NAND2_X1 U709 ( .A1(G50), .A2(n641), .ZN(n622) );
  NAND2_X1 U710 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U711 ( .A1(n625), .A2(n624), .ZN(G166) );
  AND2_X1 U712 ( .A1(n645), .A2(G60), .ZN(n629) );
  NAND2_X1 U713 ( .A1(G85), .A2(n632), .ZN(n627) );
  NAND2_X1 U714 ( .A1(G72), .A2(n635), .ZN(n626) );
  NAND2_X1 U715 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U716 ( .A1(n629), .A2(n628), .ZN(n631) );
  NAND2_X1 U717 ( .A1(n641), .A2(G47), .ZN(n630) );
  NAND2_X1 U718 ( .A1(n631), .A2(n630), .ZN(G290) );
  NAND2_X1 U719 ( .A1(G61), .A2(n645), .ZN(n634) );
  NAND2_X1 U720 ( .A1(G86), .A2(n632), .ZN(n633) );
  NAND2_X1 U721 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U722 ( .A1(n635), .A2(G73), .ZN(n636) );
  XOR2_X1 U723 ( .A(KEYINPUT2), .B(n636), .Z(n637) );
  NOR2_X1 U724 ( .A1(n638), .A2(n637), .ZN(n640) );
  NAND2_X1 U725 ( .A1(n641), .A2(G48), .ZN(n639) );
  NAND2_X1 U726 ( .A1(n640), .A2(n639), .ZN(G305) );
  NAND2_X1 U727 ( .A1(G49), .A2(n641), .ZN(n643) );
  NAND2_X1 U728 ( .A1(G74), .A2(G651), .ZN(n642) );
  NAND2_X1 U729 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U730 ( .A1(n645), .A2(n644), .ZN(n648) );
  NAND2_X1 U731 ( .A1(n646), .A2(G87), .ZN(n647) );
  NAND2_X1 U732 ( .A1(n648), .A2(n647), .ZN(G288) );
  XNOR2_X1 U733 ( .A(n973), .B(G166), .ZN(n654) );
  XOR2_X1 U734 ( .A(G290), .B(G305), .Z(n649) );
  XNOR2_X1 U735 ( .A(n658), .B(n649), .ZN(n650) );
  XNOR2_X1 U736 ( .A(KEYINPUT19), .B(n650), .ZN(n652) );
  XNOR2_X1 U737 ( .A(G288), .B(KEYINPUT82), .ZN(n651) );
  XNOR2_X1 U738 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U739 ( .A(n654), .B(n653), .ZN(n904) );
  XNOR2_X1 U740 ( .A(n904), .B(n655), .ZN(n656) );
  NOR2_X1 U741 ( .A1(n657), .A2(n656), .ZN(n660) );
  NOR2_X1 U742 ( .A1(G868), .A2(n658), .ZN(n659) );
  NOR2_X1 U743 ( .A1(n660), .A2(n659), .ZN(G295) );
  NAND2_X1 U744 ( .A1(G2084), .A2(G2078), .ZN(n661) );
  XOR2_X1 U745 ( .A(KEYINPUT20), .B(n661), .Z(n662) );
  NAND2_X1 U746 ( .A1(G2090), .A2(n662), .ZN(n663) );
  XNOR2_X1 U747 ( .A(KEYINPUT21), .B(n663), .ZN(n664) );
  NAND2_X1 U748 ( .A1(n664), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U749 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U750 ( .A1(G661), .A2(G483), .ZN(n673) );
  NOR2_X1 U751 ( .A1(G238), .A2(G236), .ZN(n665) );
  NAND2_X1 U752 ( .A1(G69), .A2(n665), .ZN(n666) );
  NOR2_X1 U753 ( .A1(n666), .A2(G237), .ZN(n667) );
  XNOR2_X1 U754 ( .A(n667), .B(KEYINPUT83), .ZN(n839) );
  NAND2_X1 U755 ( .A1(G567), .A2(n839), .ZN(n672) );
  NOR2_X1 U756 ( .A1(G220), .A2(G219), .ZN(n668) );
  XOR2_X1 U757 ( .A(KEYINPUT22), .B(n668), .Z(n669) );
  NOR2_X1 U758 ( .A1(G218), .A2(n669), .ZN(n670) );
  NAND2_X1 U759 ( .A1(G96), .A2(n670), .ZN(n840) );
  NAND2_X1 U760 ( .A1(G2106), .A2(n840), .ZN(n671) );
  NAND2_X1 U761 ( .A1(n672), .A2(n671), .ZN(n841) );
  NOR2_X1 U762 ( .A1(n673), .A2(n841), .ZN(n674) );
  XNOR2_X1 U763 ( .A(n674), .B(KEYINPUT84), .ZN(n838) );
  NAND2_X1 U764 ( .A1(G36), .A2(n838), .ZN(G176) );
  XOR2_X1 U765 ( .A(KEYINPUT86), .B(G166), .Z(G303) );
  NAND2_X1 U766 ( .A1(G160), .A2(G40), .ZN(n749) );
  INV_X1 U767 ( .A(n749), .ZN(n676) );
  INV_X1 U768 ( .A(G1384), .ZN(n675) );
  NAND2_X1 U769 ( .A1(n676), .A2(n675), .ZN(n678) );
  INV_X1 U770 ( .A(n723), .ZN(n707) );
  NAND2_X1 U771 ( .A1(n707), .A2(G1996), .ZN(n680) );
  NOR2_X1 U772 ( .A1(n681), .A2(n970), .ZN(n683) );
  NAND2_X1 U773 ( .A1(G1341), .A2(n723), .ZN(n682) );
  NAND2_X1 U774 ( .A1(n683), .A2(n682), .ZN(n691) );
  NOR2_X1 U775 ( .A1(n691), .A2(n965), .ZN(n685) );
  XNOR2_X1 U776 ( .A(n685), .B(n684), .ZN(n690) );
  AND2_X1 U777 ( .A1(n723), .A2(G1348), .ZN(n686) );
  XNOR2_X1 U778 ( .A(n686), .B(KEYINPUT95), .ZN(n688) );
  NAND2_X1 U779 ( .A1(n707), .A2(G2067), .ZN(n687) );
  NAND2_X1 U780 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U781 ( .A1(n690), .A2(n689), .ZN(n700) );
  NAND2_X1 U782 ( .A1(n691), .A2(n965), .ZN(n698) );
  NAND2_X1 U783 ( .A1(n707), .A2(G2072), .ZN(n692) );
  XNOR2_X1 U784 ( .A(KEYINPUT27), .B(n692), .ZN(n695) );
  NAND2_X1 U785 ( .A1(G1956), .A2(n723), .ZN(n693) );
  XOR2_X1 U786 ( .A(KEYINPUT92), .B(n693), .Z(n694) );
  NOR2_X1 U787 ( .A1(n695), .A2(n694), .ZN(n701) );
  NOR2_X1 U788 ( .A1(n973), .A2(n701), .ZN(n696) );
  XNOR2_X1 U789 ( .A(n696), .B(KEYINPUT28), .ZN(n703) );
  INV_X1 U790 ( .A(n703), .ZN(n697) );
  AND2_X1 U791 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U792 ( .A1(n700), .A2(n699), .ZN(n705) );
  NAND2_X1 U793 ( .A1(n973), .A2(n701), .ZN(n702) );
  OR2_X1 U794 ( .A1(n703), .A2(n702), .ZN(n704) );
  AND2_X1 U795 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U796 ( .A(n706), .B(KEYINPUT29), .ZN(n711) );
  NAND2_X1 U797 ( .A1(G1961), .A2(n723), .ZN(n709) );
  XOR2_X1 U798 ( .A(G2078), .B(KEYINPUT25), .Z(n948) );
  NAND2_X1 U799 ( .A1(n707), .A2(n948), .ZN(n708) );
  NAND2_X1 U800 ( .A1(n709), .A2(n708), .ZN(n716) );
  NOR2_X1 U801 ( .A1(G301), .A2(n716), .ZN(n710) );
  NOR2_X1 U802 ( .A1(n711), .A2(n710), .ZN(n721) );
  NOR2_X1 U803 ( .A1(G2084), .A2(n723), .ZN(n737) );
  NAND2_X1 U804 ( .A1(G8), .A2(n723), .ZN(n798) );
  NOR2_X1 U805 ( .A1(G1966), .A2(n798), .ZN(n734) );
  NOR2_X1 U806 ( .A1(n737), .A2(n734), .ZN(n712) );
  NAND2_X1 U807 ( .A1(G8), .A2(n712), .ZN(n713) );
  XNOR2_X1 U808 ( .A(KEYINPUT96), .B(n713), .ZN(n714) );
  XNOR2_X1 U809 ( .A(KEYINPUT30), .B(n714), .ZN(n715) );
  NOR2_X1 U810 ( .A1(G168), .A2(n715), .ZN(n718) );
  AND2_X1 U811 ( .A1(G301), .A2(n716), .ZN(n717) );
  NOR2_X1 U812 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U813 ( .A(n719), .B(KEYINPUT31), .ZN(n720) );
  XNOR2_X1 U814 ( .A(n722), .B(KEYINPUT97), .ZN(n733) );
  NAND2_X1 U815 ( .A1(n733), .A2(G286), .ZN(n728) );
  NOR2_X1 U816 ( .A1(G1971), .A2(n798), .ZN(n725) );
  NOR2_X1 U817 ( .A1(G2090), .A2(n723), .ZN(n724) );
  NOR2_X1 U818 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U819 ( .A1(n726), .A2(G303), .ZN(n727) );
  NAND2_X1 U820 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U821 ( .A1(n729), .A2(G8), .ZN(n730) );
  XNOR2_X1 U822 ( .A(n730), .B(KEYINPUT32), .ZN(n791) );
  NAND2_X1 U823 ( .A1(G1976), .A2(G288), .ZN(n974) );
  INV_X1 U824 ( .A(n798), .ZN(n731) );
  NAND2_X1 U825 ( .A1(n974), .A2(n731), .ZN(n742) );
  INV_X1 U826 ( .A(n742), .ZN(n732) );
  AND2_X1 U827 ( .A1(n791), .A2(n732), .ZN(n740) );
  INV_X1 U828 ( .A(n733), .ZN(n735) );
  NOR2_X1 U829 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U830 ( .A(n736), .B(KEYINPUT98), .ZN(n739) );
  NAND2_X1 U831 ( .A1(n737), .A2(G8), .ZN(n738) );
  NAND2_X1 U832 ( .A1(n739), .A2(n738), .ZN(n790) );
  NAND2_X1 U833 ( .A1(n740), .A2(n790), .ZN(n744) );
  NOR2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n783) );
  NOR2_X1 U835 ( .A1(G303), .A2(G1971), .ZN(n741) );
  NOR2_X1 U836 ( .A1(n783), .A2(n741), .ZN(n979) );
  OR2_X1 U837 ( .A1(n742), .A2(n979), .ZN(n743) );
  NAND2_X1 U838 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U839 ( .A(n745), .B(KEYINPUT64), .ZN(n746) );
  XNOR2_X1 U840 ( .A(n748), .B(n747), .ZN(n789) );
  XOR2_X1 U841 ( .A(G1981), .B(G305), .Z(n962) );
  XNOR2_X1 U842 ( .A(G1986), .B(G290), .ZN(n981) );
  NOR2_X1 U843 ( .A1(G164), .A2(G1384), .ZN(n750) );
  NOR2_X1 U844 ( .A1(n750), .A2(n749), .ZN(n818) );
  AND2_X1 U845 ( .A1(n981), .A2(n818), .ZN(n782) );
  NAND2_X1 U846 ( .A1(n886), .A2(G141), .ZN(n751) );
  XNOR2_X1 U847 ( .A(KEYINPUT90), .B(n751), .ZN(n759) );
  NAND2_X1 U848 ( .A1(G129), .A2(n882), .ZN(n753) );
  NAND2_X1 U849 ( .A1(G117), .A2(n883), .ZN(n752) );
  NAND2_X1 U850 ( .A1(n753), .A2(n752), .ZN(n756) );
  NAND2_X1 U851 ( .A1(n887), .A2(G105), .ZN(n754) );
  XOR2_X1 U852 ( .A(KEYINPUT38), .B(n754), .Z(n755) );
  NOR2_X1 U853 ( .A1(n756), .A2(n755), .ZN(n757) );
  XOR2_X1 U854 ( .A(KEYINPUT89), .B(n757), .Z(n758) );
  NAND2_X1 U855 ( .A1(n759), .A2(n758), .ZN(n870) );
  NAND2_X1 U856 ( .A1(n870), .A2(G1996), .ZN(n767) );
  NAND2_X1 U857 ( .A1(G119), .A2(n882), .ZN(n761) );
  NAND2_X1 U858 ( .A1(G131), .A2(n886), .ZN(n760) );
  NAND2_X1 U859 ( .A1(n761), .A2(n760), .ZN(n765) );
  NAND2_X1 U860 ( .A1(G107), .A2(n883), .ZN(n763) );
  NAND2_X1 U861 ( .A1(G95), .A2(n887), .ZN(n762) );
  NAND2_X1 U862 ( .A1(n763), .A2(n762), .ZN(n764) );
  OR2_X1 U863 ( .A1(n765), .A2(n764), .ZN(n895) );
  NAND2_X1 U864 ( .A1(G1991), .A2(n895), .ZN(n766) );
  NAND2_X1 U865 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U866 ( .A(n768), .B(KEYINPUT91), .ZN(n918) );
  INV_X1 U867 ( .A(n918), .ZN(n769) );
  NAND2_X1 U868 ( .A1(n769), .A2(n818), .ZN(n805) );
  NAND2_X1 U869 ( .A1(G140), .A2(n886), .ZN(n771) );
  NAND2_X1 U870 ( .A1(G104), .A2(n887), .ZN(n770) );
  NAND2_X1 U871 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U872 ( .A(KEYINPUT34), .B(n772), .ZN(n778) );
  NAND2_X1 U873 ( .A1(G128), .A2(n882), .ZN(n774) );
  NAND2_X1 U874 ( .A1(G116), .A2(n883), .ZN(n773) );
  NAND2_X1 U875 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U876 ( .A(KEYINPUT35), .B(n775), .ZN(n776) );
  XNOR2_X1 U877 ( .A(KEYINPUT87), .B(n776), .ZN(n777) );
  NOR2_X1 U878 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U879 ( .A(KEYINPUT36), .B(n779), .ZN(n899) );
  XNOR2_X1 U880 ( .A(KEYINPUT37), .B(G2067), .ZN(n815) );
  NOR2_X1 U881 ( .A1(n899), .A2(n815), .ZN(n780) );
  XNOR2_X1 U882 ( .A(n780), .B(KEYINPUT88), .ZN(n935) );
  NAND2_X1 U883 ( .A1(n818), .A2(n935), .ZN(n813) );
  NAND2_X1 U884 ( .A1(n805), .A2(n813), .ZN(n781) );
  NOR2_X1 U885 ( .A1(n782), .A2(n781), .ZN(n802) );
  AND2_X1 U886 ( .A1(n962), .A2(n802), .ZN(n787) );
  NAND2_X1 U887 ( .A1(n783), .A2(KEYINPUT33), .ZN(n784) );
  XNOR2_X1 U888 ( .A(KEYINPUT100), .B(n784), .ZN(n785) );
  NOR2_X1 U889 ( .A1(n798), .A2(n785), .ZN(n786) );
  NOR2_X1 U890 ( .A1(n789), .A2(n788), .ZN(n804) );
  NAND2_X1 U891 ( .A1(n791), .A2(n790), .ZN(n794) );
  NOR2_X1 U892 ( .A1(G2090), .A2(G303), .ZN(n792) );
  NAND2_X1 U893 ( .A1(G8), .A2(n792), .ZN(n793) );
  NAND2_X1 U894 ( .A1(n794), .A2(n793), .ZN(n795) );
  NAND2_X1 U895 ( .A1(n795), .A2(n798), .ZN(n800) );
  NOR2_X1 U896 ( .A1(G1981), .A2(G305), .ZN(n796) );
  XOR2_X1 U897 ( .A(n796), .B(KEYINPUT24), .Z(n797) );
  OR2_X1 U898 ( .A1(n798), .A2(n797), .ZN(n799) );
  NAND2_X1 U899 ( .A1(n800), .A2(n799), .ZN(n801) );
  AND2_X1 U900 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U901 ( .A1(n804), .A2(n803), .ZN(n821) );
  XOR2_X1 U902 ( .A(KEYINPUT103), .B(KEYINPUT39), .Z(n812) );
  NOR2_X1 U903 ( .A1(G1996), .A2(n870), .ZN(n925) );
  INV_X1 U904 ( .A(n805), .ZN(n808) );
  NOR2_X1 U905 ( .A1(G1991), .A2(n895), .ZN(n916) );
  NOR2_X1 U906 ( .A1(G1986), .A2(G290), .ZN(n806) );
  NOR2_X1 U907 ( .A1(n916), .A2(n806), .ZN(n807) );
  NOR2_X1 U908 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U909 ( .A(n809), .B(KEYINPUT102), .ZN(n810) );
  NOR2_X1 U910 ( .A1(n925), .A2(n810), .ZN(n811) );
  XNOR2_X1 U911 ( .A(n812), .B(n811), .ZN(n814) );
  NAND2_X1 U912 ( .A1(n814), .A2(n813), .ZN(n816) );
  NAND2_X1 U913 ( .A1(n815), .A2(n899), .ZN(n921) );
  NAND2_X1 U914 ( .A1(n816), .A2(n921), .ZN(n817) );
  XNOR2_X1 U915 ( .A(KEYINPUT104), .B(n817), .ZN(n819) );
  NAND2_X1 U916 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U917 ( .A1(n821), .A2(n820), .ZN(n824) );
  XOR2_X1 U918 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n822) );
  XNOR2_X1 U919 ( .A(KEYINPUT40), .B(n822), .ZN(n823) );
  XNOR2_X1 U920 ( .A(n824), .B(n823), .ZN(G329) );
  XNOR2_X1 U921 ( .A(G1348), .B(G2451), .ZN(n825) );
  XNOR2_X1 U922 ( .A(n825), .B(G2435), .ZN(n826) );
  XNOR2_X1 U923 ( .A(n826), .B(G1341), .ZN(n832) );
  XOR2_X1 U924 ( .A(G2446), .B(G2427), .Z(n828) );
  XNOR2_X1 U925 ( .A(G2454), .B(G2443), .ZN(n827) );
  XNOR2_X1 U926 ( .A(n828), .B(n827), .ZN(n830) );
  XOR2_X1 U927 ( .A(G2438), .B(G2430), .Z(n829) );
  XNOR2_X1 U928 ( .A(n830), .B(n829), .ZN(n831) );
  XNOR2_X1 U929 ( .A(n832), .B(n831), .ZN(n833) );
  NAND2_X1 U930 ( .A1(n833), .A2(G14), .ZN(n908) );
  XNOR2_X1 U931 ( .A(KEYINPUT107), .B(n908), .ZN(G401) );
  NAND2_X1 U932 ( .A1(n834), .A2(G2106), .ZN(n835) );
  XNOR2_X1 U933 ( .A(n835), .B(KEYINPUT108), .ZN(G217) );
  AND2_X1 U934 ( .A1(G15), .A2(G2), .ZN(n836) );
  NAND2_X1 U935 ( .A1(G661), .A2(n836), .ZN(G259) );
  NAND2_X1 U936 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U937 ( .A1(n838), .A2(n837), .ZN(G188) );
  XNOR2_X1 U938 ( .A(G69), .B(KEYINPUT109), .ZN(G235) );
  NOR2_X1 U939 ( .A1(n840), .A2(n839), .ZN(G325) );
  XOR2_X1 U940 ( .A(KEYINPUT110), .B(G325), .Z(G261) );
  INV_X1 U942 ( .A(G96), .ZN(G221) );
  XNOR2_X1 U943 ( .A(KEYINPUT111), .B(n841), .ZN(G319) );
  XNOR2_X1 U944 ( .A(G1961), .B(KEYINPUT114), .ZN(n851) );
  XOR2_X1 U945 ( .A(G1981), .B(G1956), .Z(n843) );
  XNOR2_X1 U946 ( .A(G1986), .B(G1966), .ZN(n842) );
  XNOR2_X1 U947 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U948 ( .A(G1976), .B(G1971), .Z(n845) );
  XNOR2_X1 U949 ( .A(G1996), .B(G1991), .ZN(n844) );
  XNOR2_X1 U950 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U951 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U952 ( .A(G2474), .B(KEYINPUT41), .ZN(n848) );
  XNOR2_X1 U953 ( .A(n849), .B(n848), .ZN(n850) );
  XNOR2_X1 U954 ( .A(n851), .B(n850), .ZN(G229) );
  XOR2_X1 U955 ( .A(G2100), .B(KEYINPUT43), .Z(n853) );
  XNOR2_X1 U956 ( .A(KEYINPUT113), .B(KEYINPUT112), .ZN(n852) );
  XNOR2_X1 U957 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U958 ( .A(KEYINPUT42), .B(G2090), .Z(n855) );
  XNOR2_X1 U959 ( .A(G2067), .B(G2072), .ZN(n854) );
  XNOR2_X1 U960 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U961 ( .A(n857), .B(n856), .Z(n859) );
  XNOR2_X1 U962 ( .A(G2678), .B(G2096), .ZN(n858) );
  XNOR2_X1 U963 ( .A(n859), .B(n858), .ZN(n861) );
  XOR2_X1 U964 ( .A(G2084), .B(G2078), .Z(n860) );
  XNOR2_X1 U965 ( .A(n861), .B(n860), .ZN(G227) );
  NAND2_X1 U966 ( .A1(n882), .A2(G124), .ZN(n862) );
  XNOR2_X1 U967 ( .A(n862), .B(KEYINPUT44), .ZN(n864) );
  NAND2_X1 U968 ( .A1(G112), .A2(n883), .ZN(n863) );
  NAND2_X1 U969 ( .A1(n864), .A2(n863), .ZN(n868) );
  NAND2_X1 U970 ( .A1(G136), .A2(n886), .ZN(n866) );
  NAND2_X1 U971 ( .A1(G100), .A2(n887), .ZN(n865) );
  NAND2_X1 U972 ( .A1(n866), .A2(n865), .ZN(n867) );
  NOR2_X1 U973 ( .A1(n868), .A2(n867), .ZN(G162) );
  XOR2_X1 U974 ( .A(G164), .B(n915), .Z(n869) );
  XNOR2_X1 U975 ( .A(n870), .B(n869), .ZN(n879) );
  NAND2_X1 U976 ( .A1(G139), .A2(n886), .ZN(n872) );
  NAND2_X1 U977 ( .A1(G103), .A2(n887), .ZN(n871) );
  NAND2_X1 U978 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U979 ( .A(KEYINPUT116), .B(n873), .ZN(n878) );
  NAND2_X1 U980 ( .A1(G127), .A2(n882), .ZN(n875) );
  NAND2_X1 U981 ( .A1(G115), .A2(n883), .ZN(n874) );
  NAND2_X1 U982 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U983 ( .A(KEYINPUT47), .B(n876), .Z(n877) );
  NOR2_X1 U984 ( .A1(n878), .A2(n877), .ZN(n929) );
  XOR2_X1 U985 ( .A(n879), .B(n929), .Z(n881) );
  XNOR2_X1 U986 ( .A(G160), .B(G162), .ZN(n880) );
  XNOR2_X1 U987 ( .A(n881), .B(n880), .ZN(n901) );
  XNOR2_X1 U988 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n897) );
  NAND2_X1 U989 ( .A1(G130), .A2(n882), .ZN(n885) );
  NAND2_X1 U990 ( .A1(G118), .A2(n883), .ZN(n884) );
  NAND2_X1 U991 ( .A1(n885), .A2(n884), .ZN(n893) );
  NAND2_X1 U992 ( .A1(G142), .A2(n886), .ZN(n889) );
  NAND2_X1 U993 ( .A1(G106), .A2(n887), .ZN(n888) );
  NAND2_X1 U994 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U995 ( .A(KEYINPUT45), .B(n890), .ZN(n891) );
  XNOR2_X1 U996 ( .A(KEYINPUT115), .B(n891), .ZN(n892) );
  NOR2_X1 U997 ( .A1(n893), .A2(n892), .ZN(n894) );
  XNOR2_X1 U998 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U999 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U1000 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U1001 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n902), .ZN(G395) );
  XNOR2_X1 U1003 ( .A(G171), .B(n965), .ZN(n903) );
  XNOR2_X1 U1004 ( .A(n903), .B(G286), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(n970), .B(n904), .ZN(n905) );
  XNOR2_X1 U1006 ( .A(n906), .B(n905), .ZN(n907) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n907), .ZN(G397) );
  NAND2_X1 U1008 ( .A1(G319), .A2(n908), .ZN(n911) );
  NOR2_X1 U1009 ( .A1(G229), .A2(G227), .ZN(n909) );
  XNOR2_X1 U1010 ( .A(n909), .B(KEYINPUT49), .ZN(n910) );
  NOR2_X1 U1011 ( .A1(n911), .A2(n910), .ZN(n912) );
  XOR2_X1 U1012 ( .A(KEYINPUT117), .B(n912), .Z(n914) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n913) );
  NAND2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  NOR2_X1 U1016 ( .A1(n916), .A2(n915), .ZN(n917) );
  NAND2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n920) );
  XOR2_X1 U1018 ( .A(G160), .B(G2084), .Z(n919) );
  NOR2_X1 U1019 ( .A1(n920), .A2(n919), .ZN(n922) );
  NAND2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n928) );
  XOR2_X1 U1021 ( .A(G2090), .B(G162), .Z(n923) );
  XNOR2_X1 U1022 ( .A(KEYINPUT118), .B(n923), .ZN(n924) );
  NOR2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1024 ( .A(KEYINPUT51), .B(n926), .ZN(n927) );
  NOR2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n937) );
  XOR2_X1 U1026 ( .A(G2072), .B(n929), .Z(n931) );
  XOR2_X1 U1027 ( .A(G164), .B(G2078), .Z(n930) );
  NOR2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1029 ( .A(n932), .B(KEYINPUT119), .ZN(n933) );
  XNOR2_X1 U1030 ( .A(KEYINPUT50), .B(n933), .ZN(n934) );
  NOR2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1033 ( .A(KEYINPUT52), .B(n938), .ZN(n939) );
  NAND2_X1 U1034 ( .A1(n939), .A2(G29), .ZN(n1018) );
  XNOR2_X1 U1035 ( .A(G1991), .B(G25), .ZN(n941) );
  XNOR2_X1 U1036 ( .A(G33), .B(G2072), .ZN(n940) );
  NOR2_X1 U1037 ( .A1(n941), .A2(n940), .ZN(n947) );
  XOR2_X1 U1038 ( .A(G1996), .B(G32), .Z(n942) );
  NAND2_X1 U1039 ( .A1(n942), .A2(G28), .ZN(n945) );
  XNOR2_X1 U1040 ( .A(KEYINPUT120), .B(G2067), .ZN(n943) );
  XNOR2_X1 U1041 ( .A(G26), .B(n943), .ZN(n944) );
  NOR2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n951) );
  XOR2_X1 U1044 ( .A(G27), .B(n948), .Z(n949) );
  XNOR2_X1 U1045 ( .A(KEYINPUT121), .B(n949), .ZN(n950) );
  NOR2_X1 U1046 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1047 ( .A(KEYINPUT53), .B(n952), .Z(n955) );
  XOR2_X1 U1048 ( .A(KEYINPUT54), .B(G34), .Z(n953) );
  XNOR2_X1 U1049 ( .A(G2084), .B(n953), .ZN(n954) );
  NAND2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(G35), .B(G2090), .ZN(n956) );
  NOR2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(n958), .B(KEYINPUT122), .ZN(n959) );
  NOR2_X1 U1054 ( .A1(G29), .A2(n959), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(KEYINPUT55), .B(n960), .ZN(n961) );
  NAND2_X1 U1056 ( .A1(n961), .A2(G11), .ZN(n1016) );
  XNOR2_X1 U1057 ( .A(G16), .B(KEYINPUT56), .ZN(n986) );
  XNOR2_X1 U1058 ( .A(G1966), .B(G168), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1060 ( .A(KEYINPUT57), .B(n964), .ZN(n969) );
  XNOR2_X1 U1061 ( .A(G301), .B(G1961), .ZN(n967) );
  XNOR2_X1 U1062 ( .A(n965), .B(G1348), .ZN(n966) );
  NOR2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(G1341), .B(n970), .ZN(n971) );
  NOR2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n984) );
  XNOR2_X1 U1067 ( .A(n973), .B(G1956), .ZN(n975) );
  NAND2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n977) );
  AND2_X1 U1069 ( .A1(G303), .A2(G1971), .ZN(n976) );
  NOR2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1073 ( .A(KEYINPUT123), .B(n982), .Z(n983) );
  NAND2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n1014) );
  INV_X1 U1076 ( .A(G16), .ZN(n1012) );
  XNOR2_X1 U1077 ( .A(KEYINPUT127), .B(KEYINPUT61), .ZN(n1010) );
  XNOR2_X1 U1078 ( .A(KEYINPUT125), .B(G1966), .ZN(n987) );
  XNOR2_X1 U1079 ( .A(n987), .B(G21), .ZN(n1008) );
  XOR2_X1 U1080 ( .A(G1961), .B(G5), .Z(n998) );
  XOR2_X1 U1081 ( .A(G1956), .B(G20), .Z(n992) );
  XNOR2_X1 U1082 ( .A(G1341), .B(G19), .ZN(n989) );
  XNOR2_X1 U1083 ( .A(G6), .B(G1981), .ZN(n988) );
  NOR2_X1 U1084 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1085 ( .A(KEYINPUT124), .B(n990), .ZN(n991) );
  NAND2_X1 U1086 ( .A1(n992), .A2(n991), .ZN(n995) );
  XOR2_X1 U1087 ( .A(G4), .B(G1348), .Z(n993) );
  XNOR2_X1 U1088 ( .A(KEYINPUT59), .B(n993), .ZN(n994) );
  NOR2_X1 U1089 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1090 ( .A(KEYINPUT60), .B(n996), .ZN(n997) );
  NAND2_X1 U1091 ( .A1(n998), .A2(n997), .ZN(n1006) );
  XNOR2_X1 U1092 ( .A(G1986), .B(G24), .ZN(n1000) );
  XNOR2_X1 U1093 ( .A(G23), .B(G1976), .ZN(n999) );
  NOR2_X1 U1094 ( .A1(n1000), .A2(n999), .ZN(n1003) );
  XOR2_X1 U1095 ( .A(G1971), .B(KEYINPUT126), .Z(n1001) );
  XNOR2_X1 U1096 ( .A(G22), .B(n1001), .ZN(n1002) );
  NAND2_X1 U1097 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1098 ( .A(KEYINPUT58), .B(n1004), .ZN(n1005) );
  NOR2_X1 U1099 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1100 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1101 ( .A(n1010), .B(n1009), .ZN(n1011) );
  NAND2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1106 ( .A(KEYINPUT62), .B(n1019), .Z(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

