//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 0 1 0 0 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1225,
    new_n1226, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G116), .A2(G270), .ZN(new_n206));
  INV_X1    g0006(.A(G77), .ZN(new_n207));
  INV_X1    g0007(.A(G244), .ZN(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n206), .B1(new_n207), .B2(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(G226), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n212), .B1(new_n202), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n211), .B(new_n216), .C1(G97), .C2(G257), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n217), .B1(G1), .B2(G20), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT64), .Z(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n222), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT0), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(G50), .B1(G58), .B2(G68), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  AOI22_X1  g0030(.A1(new_n219), .A2(KEYINPUT1), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n221), .A2(new_n225), .A3(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G264), .ZN(new_n240));
  XOR2_X1   g0040(.A(KEYINPUT65), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n238), .B(new_n242), .Z(G358));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT67), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT66), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G68), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n247), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(G179), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT3), .B(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n235), .A2(G1698), .ZN(new_n255));
  OAI211_X1 g0055(.A(new_n254), .B(new_n255), .C1(G226), .C2(G1698), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G97), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AND2_X1   g0058(.A1(G1), .A2(G13), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT13), .ZN(new_n264));
  OR2_X1    g0064(.A1(KEYINPUT69), .A2(G1), .ZN(new_n265));
  NAND2_X1  g0065(.A1(KEYINPUT69), .A2(G1), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G41), .ZN(new_n268));
  AND2_X1   g0068(.A1(KEYINPUT69), .A2(G1), .ZN(new_n269));
  NOR2_X1   g0069(.A1(KEYINPUT69), .A2(G1), .ZN(new_n270));
  OAI21_X1  g0070(.A(G45), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n268), .A2(G238), .A3(new_n261), .A4(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G1), .ZN(new_n273));
  OR2_X1    g0073(.A1(KEYINPUT68), .A2(G41), .ZN(new_n274));
  NAND2_X1  g0074(.A1(KEYINPUT68), .A2(G41), .ZN(new_n275));
  AND2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n273), .B(G274), .C1(new_n276), .C2(G45), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n263), .A2(new_n264), .A3(new_n272), .A4(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n272), .A2(new_n277), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n261), .B1(new_n256), .B2(new_n257), .ZN(new_n280));
  OAI21_X1  g0080(.A(KEYINPUT13), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n278), .A2(new_n281), .A3(KEYINPUT76), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT76), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n283), .B(KEYINPUT13), .C1(new_n279), .C2(new_n280), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n253), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT14), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n278), .A2(new_n281), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n286), .B1(new_n287), .B2(G169), .ZN(new_n288));
  INV_X1    g0088(.A(G169), .ZN(new_n289));
  AOI211_X1 g0089(.A(KEYINPUT14), .B(new_n289), .C1(new_n278), .C2(new_n281), .ZN(new_n290));
  NOR3_X1   g0090(.A1(new_n285), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G20), .A2(G33), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(new_n202), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n227), .A2(G68), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n227), .A2(G33), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n296), .B(KEYINPUT71), .ZN(new_n297));
  AOI211_X1 g0097(.A(new_n294), .B(new_n295), .C1(new_n297), .C2(G77), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT11), .ZN(new_n299));
  NAND3_X1  g0099(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n226), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  OR3_X1    g0102(.A1(new_n298), .A2(new_n299), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n301), .B1(new_n267), .B2(G20), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G68), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n299), .B1(new_n298), .B2(new_n302), .ZN(new_n306));
  OAI211_X1 g0106(.A(G13), .B(G20), .C1(new_n269), .C2(new_n270), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n214), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n309), .B(KEYINPUT12), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n303), .A2(new_n305), .A3(new_n306), .A4(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n291), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G190), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n315), .B1(new_n282), .B2(new_n284), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G200), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n318), .B1(new_n278), .B2(new_n281), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n317), .A2(new_n312), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n314), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G33), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT3), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT3), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G33), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G1698), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n327), .B1(G222), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G223), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n329), .B1(new_n330), .B2(new_n328), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n331), .B(new_n262), .C1(G77), .C2(new_n254), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n268), .A2(new_n261), .A3(new_n271), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n332), .B(new_n277), .C1(new_n213), .C2(new_n333), .ZN(new_n334));
  OR2_X1    g0134(.A1(new_n334), .A2(new_n315), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(G200), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n307), .A2(G50), .ZN(new_n337));
  INV_X1    g0137(.A(new_n304), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n338), .A2(new_n202), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n203), .A2(G20), .ZN(new_n340));
  INV_X1    g0140(.A(G150), .ZN(new_n341));
  INV_X1    g0141(.A(G58), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(KEYINPUT70), .A3(KEYINPUT8), .ZN(new_n343));
  XOR2_X1   g0143(.A(KEYINPUT8), .B(G58), .Z(new_n344));
  OAI21_X1  g0144(.A(new_n343), .B1(new_n344), .B2(KEYINPUT70), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT71), .ZN(new_n346));
  XNOR2_X1  g0146(.A(new_n296), .B(new_n346), .ZN(new_n347));
  OAI221_X1 g0147(.A(new_n340), .B1(new_n341), .B2(new_n293), .C1(new_n345), .C2(new_n347), .ZN(new_n348));
  AOI211_X1 g0148(.A(new_n337), .B(new_n339), .C1(new_n348), .C2(new_n301), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT9), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n349), .A2(new_n350), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n335), .B(new_n336), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(KEYINPUT75), .A2(KEYINPUT10), .ZN(new_n355));
  OR2_X1    g0155(.A1(KEYINPUT75), .A2(KEYINPUT10), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n337), .B1(new_n348), .B2(new_n301), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(new_n202), .B2(new_n338), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(KEYINPUT9), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n360), .A2(new_n351), .B1(G200), .B2(new_n334), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n361), .A2(KEYINPUT75), .A3(KEYINPUT10), .A4(new_n335), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n334), .A2(new_n289), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n363), .B(new_n359), .C1(G179), .C2(new_n334), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n357), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n322), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n327), .A2(new_n227), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT7), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT77), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n325), .B2(G33), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n323), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(new_n326), .A3(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n368), .A2(G20), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n367), .A2(new_n368), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(KEYINPUT78), .B1(new_n374), .B2(new_n214), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n342), .A2(new_n214), .ZN(new_n376));
  OAI21_X1  g0176(.A(G20), .B1(new_n376), .B2(new_n201), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n292), .A2(G159), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n372), .A2(new_n373), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n368), .B1(new_n254), .B2(G20), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT78), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(new_n384), .A3(G68), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n375), .A2(new_n380), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT16), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n327), .A2(new_n373), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n382), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n379), .B1(new_n390), .B2(G68), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n302), .B1(new_n391), .B2(KEYINPUT16), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n345), .A2(new_n304), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n394), .B1(new_n307), .B2(new_n345), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n277), .B1(new_n333), .B2(new_n235), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n213), .A2(G1698), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n254), .B(new_n398), .C1(G223), .C2(G1698), .ZN(new_n399));
  NAND2_X1  g0199(.A1(G33), .A2(G87), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n261), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G190), .ZN(new_n403));
  OAI21_X1  g0203(.A(G200), .B1(new_n397), .B2(new_n401), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n393), .A2(new_n396), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT17), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n393), .A2(new_n396), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT18), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n402), .A2(G179), .ZN(new_n410));
  OAI21_X1  g0210(.A(G169), .B1(new_n397), .B2(new_n401), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n408), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n395), .B1(new_n388), .B2(new_n392), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n410), .A2(new_n411), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT18), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n414), .A2(KEYINPUT17), .A3(new_n403), .A4(new_n404), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n407), .A2(new_n413), .A3(new_n416), .A4(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n327), .B1(G232), .B2(new_n328), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n215), .B2(new_n328), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n421), .B(new_n262), .C1(G107), .C2(new_n254), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n268), .A2(G244), .A3(new_n261), .A4(new_n271), .ZN(new_n423));
  AND3_X1   g0223(.A1(new_n423), .A2(new_n277), .A3(KEYINPUT72), .ZN(new_n424));
  AOI21_X1  g0224(.A(KEYINPUT72), .B1(new_n423), .B2(new_n277), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n422), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OR2_X1    g0226(.A1(new_n426), .A2(new_n315), .ZN(new_n427));
  NAND2_X1  g0227(.A1(G20), .A2(G77), .ZN(new_n428));
  OR2_X1    g0228(.A1(KEYINPUT15), .A2(G87), .ZN(new_n429));
  NAND2_X1  g0229(.A1(KEYINPUT15), .A2(G87), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT74), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n429), .A2(KEYINPUT74), .A3(new_n430), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g0235(.A(new_n344), .B(KEYINPUT73), .ZN(new_n436));
  OAI221_X1 g0236(.A(new_n428), .B1(new_n435), .B2(new_n296), .C1(new_n436), .C2(new_n293), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n437), .A2(new_n301), .B1(new_n207), .B2(new_n308), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n304), .A2(G77), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n426), .A2(G200), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n427), .A2(new_n438), .A3(new_n439), .A4(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n426), .A2(G169), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n422), .B(G179), .C1(new_n425), .C2(new_n424), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n438), .A2(new_n439), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n441), .A2(new_n446), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n366), .A2(new_n419), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n271), .A2(G250), .A3(new_n261), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT79), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT79), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n271), .A2(new_n451), .A3(G250), .A4(new_n261), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(G45), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n454), .B1(new_n265), .B2(new_n266), .ZN(new_n455));
  INV_X1    g0255(.A(G274), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n456), .B1(new_n259), .B2(new_n260), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(G116), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n323), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(G238), .A2(G1698), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n461), .B1(new_n208), .B2(G1698), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n460), .B1(new_n462), .B2(new_n254), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n458), .B1(new_n463), .B2(new_n261), .ZN(new_n464));
  OAI21_X1  g0264(.A(G169), .B1(new_n453), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n460), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n208), .A2(G1698), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(G238), .B2(G1698), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n466), .B1(new_n468), .B2(new_n327), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n469), .A2(new_n262), .B1(new_n455), .B2(new_n457), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n470), .A2(G179), .A3(new_n450), .A4(new_n452), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT80), .ZN(new_n473));
  OAI21_X1  g0273(.A(G33), .B1(new_n269), .B2(new_n270), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n307), .A2(new_n302), .A3(new_n474), .ZN(new_n475));
  OR3_X1    g0275(.A1(new_n435), .A2(new_n475), .A3(KEYINPUT82), .ZN(new_n476));
  OAI21_X1  g0276(.A(KEYINPUT82), .B1(new_n435), .B2(new_n475), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n227), .ZN(new_n480));
  INV_X1    g0280(.A(G97), .ZN(new_n481));
  INV_X1    g0281(.A(G107), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n209), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT81), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n324), .A2(new_n326), .A3(new_n227), .A4(G68), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT19), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(new_n296), .B2(new_n481), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n480), .A2(KEYINPUT81), .A3(new_n483), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n486), .A2(new_n487), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n491), .A2(new_n301), .B1(new_n308), .B2(new_n435), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n478), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT80), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n465), .A2(new_n471), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n473), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n324), .A2(new_n326), .A3(new_n227), .A4(G87), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT22), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n254), .A2(KEYINPUT22), .A3(new_n227), .A4(G87), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT84), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n502), .A2(KEYINPUT23), .A3(G107), .ZN(new_n503));
  AOI21_X1  g0303(.A(KEYINPUT84), .B1(new_n482), .B2(G20), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n502), .A2(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n505));
  OAI221_X1 g0305(.A(new_n503), .B1(new_n504), .B2(KEYINPUT23), .C1(G20), .C2(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(KEYINPUT24), .B1(new_n501), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n505), .A2(G20), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n482), .A2(G20), .ZN(new_n509));
  AOI21_X1  g0309(.A(KEYINPUT23), .B1(new_n509), .B2(new_n502), .ZN(new_n510));
  INV_X1    g0310(.A(new_n503), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n508), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT24), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n512), .A2(new_n513), .A3(new_n499), .A4(new_n500), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n302), .B1(new_n507), .B2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(KEYINPUT25), .B1(new_n308), .B2(new_n482), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT25), .ZN(new_n517));
  NOR3_X1   g0317(.A1(new_n307), .A2(new_n517), .A3(G107), .ZN(new_n518));
  OAI22_X1  g0318(.A1(new_n516), .A2(new_n518), .B1(new_n482), .B2(new_n475), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n328), .A2(G257), .ZN(new_n521));
  NOR2_X1   g0321(.A1(G250), .A2(G1698), .ZN(new_n522));
  NOR3_X1   g0322(.A1(new_n327), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(G294), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n323), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n262), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT5), .ZN(new_n527));
  OR2_X1    g0327(.A1(new_n527), .A2(G41), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n274), .A2(new_n527), .A3(new_n275), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n455), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n530), .A2(G264), .A3(new_n261), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n455), .A2(new_n529), .A3(new_n457), .A4(new_n528), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n526), .A2(new_n531), .A3(new_n315), .A4(new_n532), .ZN(new_n533));
  AND3_X1   g0333(.A1(new_n526), .A2(new_n531), .A3(new_n532), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n533), .B1(new_n534), .B2(G200), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n520), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n526), .A2(new_n531), .A3(new_n253), .A4(new_n532), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n526), .A2(new_n531), .A3(new_n532), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n289), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n537), .B(new_n539), .C1(new_n515), .C2(new_n519), .ZN(new_n540));
  OAI21_X1  g0340(.A(G200), .B1(new_n453), .B2(new_n464), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n470), .A2(G190), .A3(new_n450), .A4(new_n452), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OR2_X1    g0343(.A1(new_n475), .A2(new_n209), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n435), .A2(new_n308), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n487), .A2(new_n489), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n480), .A2(KEYINPUT81), .A3(new_n483), .ZN(new_n547));
  AOI21_X1  g0347(.A(KEYINPUT81), .B1(new_n480), .B2(new_n483), .ZN(new_n548));
  NOR3_X1   g0348(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n544), .B(new_n545), .C1(new_n549), .C2(new_n302), .ZN(new_n550));
  OR2_X1    g0350(.A1(new_n543), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n496), .A2(new_n536), .A3(new_n540), .A4(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n308), .A2(new_n459), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n307), .A2(new_n302), .A3(new_n474), .A4(G116), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n300), .A2(new_n226), .B1(G20), .B2(new_n459), .ZN(new_n555));
  NAND2_X1  g0355(.A1(G33), .A2(G283), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n556), .B(new_n227), .C1(G33), .C2(new_n481), .ZN(new_n557));
  AND3_X1   g0357(.A1(new_n555), .A2(KEYINPUT20), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(KEYINPUT20), .B1(new_n555), .B2(new_n557), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n553), .B(new_n554), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(G303), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n327), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n328), .A2(G257), .ZN(new_n563));
  NAND2_X1  g0363(.A1(G264), .A2(G1698), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n324), .A2(new_n326), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n562), .A2(new_n262), .A3(new_n565), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n566), .A2(new_n532), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n530), .A2(G270), .A3(new_n261), .ZN(new_n568));
  AND4_X1   g0368(.A1(G179), .A2(new_n560), .A3(new_n567), .A4(new_n568), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n530), .A2(G270), .A3(new_n261), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n566), .A2(new_n532), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n560), .B(G169), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(KEYINPUT21), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n567), .A2(new_n568), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT21), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n574), .A2(new_n575), .A3(G169), .A4(new_n560), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n569), .B1(new_n573), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT83), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n318), .B1(new_n567), .B2(new_n568), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n578), .B1(new_n579), .B2(new_n560), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n570), .A2(new_n571), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G190), .ZN(new_n582));
  INV_X1    g0382(.A(new_n560), .ZN(new_n583));
  OAI211_X1 g0383(.A(KEYINPUT83), .B(new_n583), .C1(new_n581), .C2(new_n318), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n580), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n324), .A2(new_n326), .A3(G244), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT4), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n587), .A2(G1698), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n254), .A2(G244), .A3(new_n589), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n588), .A2(new_n590), .A3(new_n556), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n254), .A2(G250), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT4), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(G1698), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n261), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n530), .A2(G257), .A3(new_n261), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n532), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n289), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT6), .ZN(new_n599));
  AND2_X1   g0399(.A1(G97), .A2(G107), .ZN(new_n600));
  NOR2_X1   g0400(.A1(G97), .A2(G107), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n482), .A2(KEYINPUT6), .A3(G97), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI22_X1  g0404(.A1(new_n604), .A2(new_n227), .B1(new_n207), .B2(new_n293), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n482), .B1(new_n381), .B2(new_n382), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n301), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n307), .A2(G97), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(new_n475), .B2(new_n481), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n596), .A2(new_n532), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n588), .A2(new_n590), .A3(new_n556), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n328), .B1(new_n592), .B2(KEYINPUT4), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n262), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n613), .A2(new_n253), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n598), .A2(new_n612), .A3(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(G200), .B1(new_n595), .B2(new_n597), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n602), .A2(new_n603), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n620), .A2(G20), .B1(G77), .B2(new_n292), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n374), .B2(new_n482), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n610), .B1(new_n622), .B2(new_n301), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n613), .A2(G190), .A3(new_n616), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n619), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n577), .A2(new_n585), .A3(new_n618), .A4(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n552), .A2(new_n626), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n448), .A2(new_n627), .ZN(G372));
  NOR3_X1   g0428(.A1(new_n316), .A2(new_n311), .A3(new_n319), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n314), .B1(new_n629), .B2(new_n446), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n630), .A2(new_n407), .A3(new_n417), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n413), .A2(new_n416), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n357), .B(new_n362), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n633), .A2(new_n364), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n598), .A2(new_n612), .A3(new_n617), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n496), .A2(new_n635), .A3(new_n551), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT26), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n550), .A2(KEYINPUT85), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT85), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n492), .A2(new_n639), .A3(new_n544), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n543), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n478), .A2(new_n492), .B1(new_n465), .B2(new_n471), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n641), .A2(new_n618), .A3(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT26), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n618), .A2(new_n625), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n573), .A2(new_n576), .ZN(new_n647));
  INV_X1    g0447(.A(new_n569), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(new_n648), .A3(new_n540), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n638), .A2(new_n640), .ZN(new_n650));
  INV_X1    g0450(.A(new_n543), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n650), .A2(new_n651), .B1(new_n520), .B2(new_n535), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n646), .A2(new_n649), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n642), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n637), .A2(new_n645), .A3(new_n653), .A4(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n448), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n634), .A2(new_n656), .ZN(G369));
  INV_X1    g0457(.A(G13), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n658), .A2(G20), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n267), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT27), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT86), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n660), .A2(new_n663), .A3(new_n661), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n663), .B1(new_n660), .B2(new_n661), .ZN(new_n665));
  OAI211_X1 g0465(.A(G213), .B(new_n662), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(G343), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n560), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n577), .A2(new_n585), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(new_n577), .B2(new_n669), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(G330), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n536), .A2(new_n540), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n668), .B1(new_n515), .B2(new_n519), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n668), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n676), .B1(new_n540), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n673), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n676), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n577), .A2(new_n668), .ZN(new_n681));
  INV_X1    g0481(.A(new_n540), .ZN(new_n682));
  AOI22_X1  g0482(.A1(new_n680), .A2(new_n681), .B1(new_n682), .B2(new_n677), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n679), .A2(new_n683), .ZN(G399));
  INV_X1    g0484(.A(new_n223), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n276), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n483), .A2(G116), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G1), .A3(new_n688), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n689), .A2(KEYINPUT87), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(KEYINPUT87), .ZN(new_n691));
  OAI211_X1 g0491(.A(new_n690), .B(new_n691), .C1(new_n229), .C2(new_n687), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT28), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n655), .A2(new_n677), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(KEYINPUT29), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n650), .A2(new_n651), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n696), .A2(new_n635), .A3(new_n654), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(KEYINPUT26), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n496), .A2(new_n644), .A3(new_n635), .A4(new_n551), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n698), .A2(new_n653), .A3(new_n654), .A4(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT89), .ZN(new_n701));
  AND3_X1   g0501(.A1(new_n700), .A2(new_n701), .A3(new_n677), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n701), .B1(new_n700), .B2(new_n677), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n695), .B1(new_n704), .B2(KEYINPUT29), .ZN(new_n705));
  AND4_X1   g0505(.A1(new_n577), .A2(new_n585), .A3(new_n618), .A4(new_n625), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n496), .A2(new_n551), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n706), .A2(new_n674), .A3(new_n707), .A4(new_n677), .ZN(new_n708));
  AND4_X1   g0508(.A1(new_n568), .A2(new_n567), .A3(new_n526), .A4(new_n531), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n595), .A2(new_n597), .ZN(new_n710));
  INV_X1    g0510(.A(new_n471), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT30), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(KEYINPUT88), .A3(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n710), .A2(new_n534), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n470), .A2(new_n450), .A3(new_n452), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n715), .A2(new_n253), .A3(new_n574), .A4(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n713), .A2(KEYINPUT88), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n709), .A2(new_n710), .A3(new_n711), .A4(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n714), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(new_n668), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n708), .A2(KEYINPUT31), .A3(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT31), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n720), .A2(new_n723), .A3(new_n668), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n722), .A2(G330), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n705), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n693), .B1(new_n727), .B2(G1), .ZN(G364));
  NAND2_X1  g0528(.A1(new_n659), .A2(G45), .ZN(new_n729));
  XOR2_X1   g0529(.A(new_n729), .B(KEYINPUT90), .Z(new_n730));
  NAND3_X1  g0530(.A1(new_n730), .A2(G1), .A3(new_n687), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n673), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(G330), .B2(new_n671), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n226), .B1(G20), .B2(new_n289), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n315), .A2(new_n318), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n227), .A2(G179), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n327), .B1(new_n738), .B2(new_n561), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT94), .ZN(new_n740));
  NAND2_X1  g0540(.A1(G20), .A2(G179), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT93), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(new_n736), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G326), .ZN(new_n745));
  INV_X1    g0545(.A(G322), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n315), .A2(G200), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n742), .A2(new_n747), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n740), .B(new_n745), .C1(new_n746), .C2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n742), .A2(new_n315), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n318), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(G317), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n752), .B1(KEYINPUT33), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n754), .B1(KEYINPUT33), .B2(new_n753), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n227), .B1(new_n747), .B2(new_n253), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n737), .A2(new_n315), .A3(new_n318), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI22_X1  g0559(.A1(G294), .A2(new_n757), .B1(new_n759), .B2(G329), .ZN(new_n760));
  INV_X1    g0560(.A(G311), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n750), .A2(G200), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n755), .B(new_n760), .C1(new_n761), .C2(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n737), .A2(new_n315), .A3(G200), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI211_X1 g0566(.A(new_n749), .B(new_n764), .C1(G283), .C2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(G159), .ZN(new_n768));
  OR3_X1    g0568(.A1(new_n758), .A2(KEYINPUT32), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(KEYINPUT32), .B1(new_n758), .B2(new_n768), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n769), .B(new_n770), .C1(new_n202), .C2(new_n743), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n756), .A2(new_n481), .ZN(new_n772));
  INV_X1    g0572(.A(new_n738), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n327), .B(new_n772), .C1(G87), .C2(new_n773), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n762), .A2(G77), .B1(G107), .B2(new_n766), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n774), .B(new_n775), .C1(new_n214), .C2(new_n752), .ZN(new_n776));
  INV_X1    g0576(.A(new_n748), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n771), .B(new_n776), .C1(G58), .C2(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n735), .B1(new_n767), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G13), .A2(G33), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT91), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(G20), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n779), .B1(new_n671), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n251), .A2(G45), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n685), .A2(new_n254), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n786), .B(new_n787), .C1(G45), .C2(new_n229), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n685), .A2(new_n327), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G355), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n788), .B(new_n790), .C1(G116), .C2(new_n223), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n783), .A2(new_n735), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n731), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n793), .B(KEYINPUT92), .Z(new_n794));
  OAI21_X1  g0594(.A(new_n734), .B1(new_n785), .B2(new_n794), .ZN(G396));
  OAI21_X1  g0595(.A(KEYINPUT97), .B1(new_n446), .B2(new_n677), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n445), .A2(new_n668), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n441), .A2(new_n446), .A3(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT97), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n444), .A2(new_n445), .A3(new_n799), .A4(new_n668), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n796), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n694), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n655), .A2(new_n801), .A3(new_n677), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  AND3_X1   g0605(.A1(new_n722), .A2(G330), .A3(new_n724), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n731), .ZN(new_n808));
  INV_X1    g0608(.A(G132), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n254), .B1(new_n758), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT96), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n757), .A2(G58), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n766), .A2(G68), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n812), .A2(new_n813), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n751), .A2(G150), .B1(new_n777), .B2(G143), .ZN(new_n817));
  INV_X1    g0617(.A(G137), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n817), .B1(new_n818), .B2(new_n743), .C1(new_n768), .C2(new_n763), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT34), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n816), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n821), .B1(new_n820), .B2(new_n819), .C1(new_n202), .C2(new_n738), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n327), .B1(new_n738), .B2(new_n482), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT95), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n524), .A2(new_n748), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(G303), .B2(new_n744), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n758), .A2(new_n761), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n772), .B(new_n827), .C1(new_n751), .C2(G283), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n823), .A2(new_n824), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n762), .A2(G116), .B1(G87), .B2(new_n766), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n826), .A2(new_n828), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n822), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n735), .A2(new_n780), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n832), .A2(new_n735), .B1(new_n207), .B2(new_n833), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n834), .B(new_n732), .C1(new_n782), .C2(new_n801), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n808), .A2(new_n835), .ZN(G384));
  INV_X1    g0636(.A(new_n448), .ZN(new_n837));
  OR2_X1    g0637(.A1(new_n837), .A2(new_n705), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n634), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT39), .ZN(new_n840));
  INV_X1    g0640(.A(new_n666), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n367), .A2(new_n368), .B1(new_n327), .B2(new_n373), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n380), .B1(new_n842), .B2(new_n214), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n387), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n395), .B1(new_n392), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT98), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n845), .A2(new_n846), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n418), .A2(new_n841), .A3(new_n849), .ZN(new_n850));
  AND3_X1   g0650(.A1(new_n410), .A2(new_n666), .A3(new_n411), .ZN(new_n851));
  NOR3_X1   g0651(.A1(new_n847), .A2(new_n848), .A3(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n405), .ZN(new_n853));
  OAI21_X1  g0653(.A(KEYINPUT37), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT37), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n405), .B(new_n855), .C1(new_n414), .C2(new_n851), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  AND3_X1   g0657(.A1(new_n850), .A2(new_n857), .A3(KEYINPUT38), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n418), .A2(new_n408), .A3(new_n841), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n414), .A2(new_n851), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT37), .B1(new_n853), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n856), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT38), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n840), .B1(new_n858), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n850), .A2(new_n857), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT38), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n850), .A2(new_n857), .A3(KEYINPUT38), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n867), .A2(KEYINPUT39), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n314), .A2(new_n668), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n864), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n446), .A2(new_n668), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n804), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n285), .ZN(new_n875));
  INV_X1    g0675(.A(new_n290), .ZN(new_n876));
  INV_X1    g0676(.A(new_n288), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n311), .B(new_n668), .C1(new_n878), .C2(new_n629), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n311), .A2(new_n668), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n321), .B(new_n880), .C1(new_n291), .C2(new_n312), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n874), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n867), .A2(new_n868), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n632), .A2(new_n666), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n871), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n839), .B(new_n889), .ZN(new_n890));
  AND4_X1   g0690(.A1(new_n722), .A2(new_n724), .A3(new_n882), .A4(new_n801), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(new_n858), .B2(new_n863), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n722), .A2(new_n724), .A3(new_n882), .A4(new_n801), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n893), .A2(KEYINPUT40), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n892), .A2(KEYINPUT40), .B1(new_n885), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n724), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n723), .B1(new_n627), .B2(new_n677), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n896), .B1(new_n897), .B2(new_n721), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n448), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n895), .B(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(G330), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n890), .B(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n267), .B2(new_n659), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n459), .B1(new_n620), .B2(KEYINPUT35), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n904), .B(new_n228), .C1(KEYINPUT35), .C2(new_n620), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT36), .ZN(new_n906));
  OAI21_X1  g0706(.A(G77), .B1(new_n342), .B2(new_n214), .ZN(new_n907));
  OAI22_X1  g0707(.A1(new_n907), .A2(new_n229), .B1(G50), .B2(new_n214), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n658), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n903), .B(new_n906), .C1(new_n267), .C2(new_n909), .ZN(G367));
  NAND3_X1  g0710(.A1(new_n668), .A2(new_n638), .A3(new_n640), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n696), .A2(new_n911), .A3(new_n654), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n654), .B2(new_n911), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(KEYINPUT43), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n646), .B1(new_n623), .B2(new_n677), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n618), .B2(new_n677), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT99), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n682), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n668), .B1(new_n918), .B2(new_n618), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n916), .A2(new_n680), .A3(new_n681), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT42), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n914), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n679), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n917), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n913), .A2(KEYINPUT43), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n925), .B(KEYINPUT100), .Z(new_n926));
  XNOR2_X1  g0726(.A(new_n924), .B(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n922), .B(new_n927), .ZN(new_n928));
  XOR2_X1   g0728(.A(KEYINPUT101), .B(KEYINPUT41), .Z(new_n929));
  XNOR2_X1  g0729(.A(new_n686), .B(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n680), .A2(new_n681), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n931), .B(KEYINPUT102), .C1(new_n678), .C2(new_n681), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(KEYINPUT102), .B2(new_n931), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(new_n673), .ZN(new_n934));
  OR3_X1    g0734(.A1(new_n934), .A2(new_n726), .A3(KEYINPUT103), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n683), .A2(new_n916), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n936), .B(KEYINPUT45), .Z(new_n937));
  OAI21_X1  g0737(.A(KEYINPUT44), .B1(new_n683), .B2(new_n916), .ZN(new_n938));
  OR3_X1    g0738(.A1(new_n683), .A2(KEYINPUT44), .A3(new_n916), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n937), .A2(new_n679), .A3(new_n938), .A4(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n936), .B(KEYINPUT45), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n939), .A2(new_n938), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n923), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(KEYINPUT103), .B1(new_n726), .B2(new_n934), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n935), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n930), .B1(new_n946), .B2(new_n727), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n730), .A2(G1), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT104), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n928), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  AOI22_X1  g0750(.A1(G50), .A2(new_n762), .B1(new_n751), .B2(G159), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n756), .A2(new_n214), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n254), .B1(new_n758), .B2(new_n818), .ZN(new_n953));
  AOI211_X1 g0753(.A(new_n952), .B(new_n953), .C1(G77), .C2(new_n766), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n773), .A2(G58), .ZN(new_n955));
  AOI22_X1  g0755(.A1(G143), .A2(new_n744), .B1(new_n777), .B2(G150), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n951), .A2(new_n954), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n773), .A2(KEYINPUT46), .A3(G116), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT46), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n738), .B2(new_n459), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n958), .B(new_n960), .C1(new_n753), .C2(new_n758), .ZN(new_n961));
  AOI211_X1 g0761(.A(new_n254), .B(new_n961), .C1(G107), .C2(new_n757), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n561), .A2(new_n748), .B1(new_n743), .B2(new_n761), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT105), .ZN(new_n964));
  AOI22_X1  g0764(.A1(G283), .A2(new_n762), .B1(new_n751), .B2(G294), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n962), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n765), .A2(new_n481), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n957), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT47), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n731), .B1(new_n969), .B2(new_n735), .ZN(new_n970));
  INV_X1    g0770(.A(new_n787), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n792), .B1(new_n223), .B2(new_n435), .C1(new_n242), .C2(new_n971), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n970), .B(new_n972), .C1(new_n784), .C2(new_n913), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n950), .A2(new_n973), .ZN(G387));
  AOI21_X1  g0774(.A(new_n687), .B1(new_n935), .B2(new_n945), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n933), .B(new_n672), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n975), .B1(new_n727), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n436), .A2(G50), .ZN(new_n978));
  XNOR2_X1  g0778(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n688), .B1(new_n978), .B2(new_n979), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n214), .A2(new_n207), .ZN(new_n982));
  NOR4_X1   g0782(.A1(new_n980), .A2(new_n981), .A3(G45), .A4(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n971), .B1(new_n238), .B2(G45), .ZN(new_n984));
  INV_X1    g0784(.A(new_n688), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n984), .B1(new_n985), .B2(new_n789), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n983), .A2(new_n986), .B1(G107), .B2(new_n223), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n792), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n678), .B2(new_n784), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n967), .B1(G150), .B2(new_n759), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n990), .B1(new_n752), .B2(new_n345), .C1(new_n214), .C2(new_n763), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n435), .A2(new_n756), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(G50), .B2(new_n777), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n768), .B2(new_n743), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n738), .A2(new_n207), .ZN(new_n995));
  NOR4_X1   g0795(.A1(new_n991), .A2(new_n994), .A3(new_n327), .A4(new_n995), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT108), .Z(new_n997));
  AOI22_X1  g0797(.A1(new_n751), .A2(G311), .B1(new_n777), .B2(G317), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(new_n561), .B2(new_n763), .C1(new_n746), .C2(new_n743), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT48), .ZN(new_n1000));
  INV_X1    g0800(.A(G283), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1000), .B1(new_n1001), .B2(new_n756), .C1(new_n524), .C2(new_n738), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT49), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n254), .B1(new_n759), .B2(G326), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n765), .A2(new_n459), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n997), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n731), .B(new_n989), .C1(new_n1009), .C2(new_n735), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n976), .A2(new_n949), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT106), .Z(new_n1013));
  NAND3_X1  g0813(.A1(new_n977), .A2(new_n1011), .A3(new_n1013), .ZN(G393));
  NAND3_X1  g0814(.A1(new_n940), .A2(KEYINPUT109), .A3(new_n943), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n943), .A2(KEYINPUT109), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n949), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n247), .A2(new_n787), .B1(G97), .B2(new_n685), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n792), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n757), .A2(G77), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1021), .B1(new_n752), .B2(new_n202), .C1(new_n436), .C2(new_n763), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT110), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n341), .A2(new_n743), .B1(new_n748), .B2(new_n768), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT51), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n327), .B1(new_n773), .B2(G68), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n766), .A2(G87), .B1(new_n759), .B2(G143), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1023), .A2(new_n1025), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G116), .A2(new_n757), .B1(new_n759), .B2(G322), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n254), .B1(new_n766), .B2(G107), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1029), .B(new_n1030), .C1(new_n752), .C2(new_n561), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(G294), .B2(new_n762), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n761), .A2(new_n748), .B1(new_n743), .B2(new_n753), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT52), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1032), .B(new_n1034), .C1(new_n1001), .C2(new_n738), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1028), .A2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n731), .B1(new_n1036), .B2(new_n735), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1020), .B(new_n1037), .C1(new_n917), .C2(new_n784), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1018), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1017), .B1(new_n945), .B2(new_n935), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n946), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1039), .B1(new_n1042), .B2(new_n686), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(G390));
  INV_X1    g0844(.A(new_n870), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n864), .A2(new_n869), .B1(new_n1045), .B2(new_n883), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n806), .A2(KEYINPUT112), .A3(new_n801), .A4(new_n882), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT112), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n722), .A2(G330), .A3(new_n724), .A4(new_n801), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n882), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1048), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AND2_X1   g0851(.A1(new_n1047), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n653), .A2(new_n654), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n699), .B1(new_n643), .B2(new_n644), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n677), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(KEYINPUT89), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n700), .A2(new_n701), .A3(new_n677), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n802), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(KEYINPUT111), .B1(new_n1058), .B2(new_n872), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n801), .B1(new_n702), .B2(new_n703), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT111), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1060), .A2(new_n1061), .A3(new_n873), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1059), .A2(new_n882), .A3(new_n1062), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n858), .A2(new_n863), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1064), .A2(new_n870), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1046), .B(new_n1052), .C1(new_n1063), .C2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1046), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1066), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT113), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n725), .A2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n722), .A2(KEYINPUT113), .A3(G330), .A4(new_n724), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1073), .A2(new_n801), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n1050), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT114), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1075), .A2(KEYINPUT114), .A3(new_n1050), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1078), .A2(new_n1052), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1049), .B(new_n1050), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n874), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n899), .A2(G330), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n838), .A2(new_n1085), .A3(new_n634), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1071), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1047), .A2(new_n1051), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1068), .A2(new_n1090), .A3(new_n1069), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1046), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1091), .B1(new_n1067), .B2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1093), .A2(new_n1084), .A3(new_n1087), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1089), .A2(new_n1094), .A3(new_n686), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n731), .B1(new_n345), .B2(new_n833), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT115), .Z(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n782), .B1(new_n864), .B2(new_n869), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n459), .A2(new_n748), .B1(new_n743), .B2(new_n1001), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n759), .A2(G294), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1021), .A2(new_n815), .A3(new_n1101), .A4(new_n327), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n1100), .B(new_n1102), .C1(G87), .C2(new_n773), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n1103), .B1(new_n481), .B2(new_n763), .C1(new_n482), .C2(new_n752), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT116), .Z(new_n1105));
  NOR3_X1   g0905(.A1(new_n738), .A2(KEYINPUT53), .A3(new_n341), .ZN(new_n1106));
  INV_X1    g0906(.A(G128), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n254), .B1(new_n743), .B2(new_n1107), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1106), .B(new_n1108), .C1(G132), .C2(new_n777), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(G159), .A2(new_n757), .B1(new_n759), .B2(G125), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n202), .B2(new_n765), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(G137), .B2(new_n751), .ZN(new_n1112));
  OAI21_X1  g0912(.A(KEYINPUT53), .B1(new_n738), .B2(new_n341), .ZN(new_n1113));
  XOR2_X1   g0913(.A(KEYINPUT54), .B(G143), .Z(new_n1114));
  NAND2_X1  g0914(.A1(new_n762), .A2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1109), .A2(new_n1112), .A3(new_n1113), .A4(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1105), .A2(new_n1116), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n1098), .B(new_n1099), .C1(new_n735), .C2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n1093), .B2(new_n949), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1119), .A2(KEYINPUT117), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT117), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1121), .B(new_n1118), .C1(new_n1093), .C2(new_n949), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1095), .B1(new_n1120), .B2(new_n1122), .ZN(G378));
  AND2_X1   g0923(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1090), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n1124), .A2(new_n1125), .B1(new_n874), .B2(new_n1082), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1087), .B1(new_n1071), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n365), .A2(KEYINPUT55), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT55), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n357), .A2(new_n362), .A3(new_n1129), .A4(new_n364), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n349), .A2(new_n666), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT56), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n1128), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1132), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(G330), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1135), .B1(new_n895), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n859), .A2(new_n862), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n866), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n893), .B1(new_n1139), .B2(new_n868), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT40), .ZN(new_n1141));
  AOI21_X1  g0941(.A(KEYINPUT38), .B1(new_n850), .B2(new_n857), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n858), .A2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n898), .A2(new_n1141), .A3(new_n801), .A4(new_n882), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n1140), .A2(new_n1141), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1135), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1145), .A2(G330), .A3(new_n1146), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1137), .A2(new_n889), .A3(KEYINPUT123), .A4(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(KEYINPUT40), .B1(new_n1064), .B2(new_n893), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n885), .A2(new_n894), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1136), .B(new_n1135), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1146), .B1(new_n1145), .B2(G330), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n888), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT123), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1137), .A2(new_n889), .A3(new_n1147), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1127), .A2(KEYINPUT57), .A3(new_n1148), .A4(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT57), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1153), .A2(KEYINPUT122), .A3(new_n1155), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT122), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1160), .B(new_n888), .C1(new_n1151), .C2(new_n1152), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1086), .B1(new_n1093), .B2(new_n1084), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1158), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1157), .A2(new_n1164), .A3(new_n686), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1159), .A2(new_n949), .A3(new_n1161), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(G132), .A2(new_n751), .B1(new_n762), .B2(G137), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n744), .A2(G125), .B1(new_n773), .B2(new_n1114), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1167), .B(new_n1168), .C1(new_n1107), .C2(new_n748), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(G150), .B2(new_n757), .ZN(new_n1170));
  XOR2_X1   g0970(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n1171));
  OR2_X1    g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n759), .A2(G124), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1174));
  AOI211_X1 g0974(.A(G33), .B(G41), .C1(new_n766), .C2(G159), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n202), .B1(G33), .B2(G41), .C1(new_n276), .C2(new_n254), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n765), .A2(new_n342), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT118), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(G97), .B2(new_n751), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n482), .A2(new_n748), .B1(new_n743), .B2(new_n459), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n276), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1183), .B(new_n327), .C1(new_n1001), .C2(new_n758), .ZN(new_n1184));
  NOR4_X1   g0984(.A1(new_n1182), .A2(new_n1184), .A3(new_n952), .A4(new_n995), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1181), .B(new_n1185), .C1(new_n435), .C2(new_n763), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1186), .B(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1176), .A2(new_n1177), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n735), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n1190), .B(KEYINPUT121), .Z(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(new_n202), .B2(new_n833), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1192), .B(new_n732), .C1(new_n782), .C2(new_n1146), .ZN(new_n1193));
  AND2_X1   g0993(.A1(new_n1166), .A2(new_n1193), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n1165), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(G375));
  INV_X1    g0996(.A(new_n930), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1081), .A2(new_n1086), .A3(new_n1083), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1088), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1050), .A2(new_n780), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n763), .A2(new_n341), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n759), .A2(G128), .B1(new_n773), .B2(G159), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1202), .B1(new_n748), .B2(new_n818), .C1(new_n809), .C2(new_n743), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1201), .B(new_n1203), .C1(new_n751), .C2(new_n1114), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1179), .A2(new_n254), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT124), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1204), .B(new_n1206), .C1(new_n202), .C2(new_n756), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n738), .A2(new_n481), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n748), .A2(new_n1001), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n1209), .B(new_n992), .C1(G294), .C2(new_n744), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n327), .B1(new_n765), .B2(new_n207), .C1(new_n561), .C2(new_n758), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n751), .B2(G116), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1210), .B(new_n1212), .C1(new_n482), .C2(new_n763), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1207), .B1(new_n1208), .B2(new_n1213), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n1214), .A2(new_n735), .B1(new_n214), .B2(new_n833), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n1200), .A2(new_n732), .A3(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n1084), .B2(new_n949), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1199), .A2(new_n1217), .ZN(G381));
  AND2_X1   g1018(.A1(new_n1095), .A2(new_n1119), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1195), .A2(new_n1219), .ZN(new_n1220));
  NOR3_X1   g1020(.A1(new_n1220), .A2(G384), .A3(G381), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1043), .A2(new_n973), .A3(new_n950), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n1222), .A2(G396), .A3(G393), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1221), .A2(new_n1223), .ZN(G407));
  NAND2_X1  g1024(.A1(new_n667), .A2(G213), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT125), .Z(new_n1226));
  OAI211_X1 g1026(.A(G407), .B(G213), .C1(new_n1220), .C2(new_n1226), .ZN(G409));
  INV_X1    g1027(.A(KEYINPUT126), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1225), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT60), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1198), .A2(new_n1230), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1081), .A2(new_n1086), .A3(KEYINPUT60), .A4(new_n1083), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1231), .A2(new_n1088), .A3(new_n686), .A4(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n1217), .ZN(new_n1234));
  INV_X1    g1034(.A(G384), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1233), .A2(G384), .A3(new_n1217), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1165), .A2(G378), .A3(new_n1194), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(new_n1162), .A2(new_n1163), .A3(new_n930), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1156), .A2(new_n949), .A3(new_n1148), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1193), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1219), .B1(new_n1240), .B2(new_n1242), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n1229), .B(new_n1238), .C1(new_n1239), .C2(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1228), .B1(new_n1244), .B2(KEYINPUT63), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1239), .A2(new_n1243), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n1225), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1238), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1229), .A2(G2897), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1226), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n1248), .A2(new_n1249), .B1(new_n1250), .B2(G2897), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT61), .B1(new_n1247), .B2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1246), .A2(new_n1225), .A3(new_n1248), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT63), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1253), .A2(KEYINPUT126), .A3(new_n1254), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1246), .A2(KEYINPUT63), .A3(new_n1226), .A4(new_n1248), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1245), .A2(new_n1252), .A3(new_n1255), .A4(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(G390), .A2(G387), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(G393), .B(G396), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1258), .A2(new_n1259), .A3(new_n1222), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1259), .B1(new_n1258), .B2(new_n1222), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT62), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1253), .A2(new_n1263), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1246), .A2(KEYINPUT62), .A3(new_n1226), .A4(new_n1248), .ZN(new_n1265));
  AOI21_X1  g1065(.A(KEYINPUT61), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1246), .A2(new_n1226), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1262), .B1(new_n1251), .B2(new_n1267), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1257), .A2(new_n1262), .B1(new_n1266), .B2(new_n1268), .ZN(G405));
  NAND2_X1  g1069(.A1(new_n1238), .A2(KEYINPUT127), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1262), .A2(new_n1270), .ZN(new_n1271));
  OAI211_X1 g1071(.A(KEYINPUT127), .B(new_n1238), .C1(new_n1260), .C2(new_n1261), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1219), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1239), .B1(new_n1195), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT127), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1275), .B1(new_n1276), .B2(new_n1248), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(new_n1273), .B(new_n1277), .ZN(G402));
endmodule


