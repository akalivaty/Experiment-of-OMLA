//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 1 0 1 0 1 0 0 0 0 0 1 1 0 0 0 0 0 1 1 0 0 1 1 1 0 0 0 1 0 0 0 1 0 0 0 0 0 0 1 1 0 0 0 0 0 1 0 1 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n565, new_n566,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n624, new_n625, new_n626, new_n629, new_n631, new_n632, new_n634,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1173, new_n1174, new_n1176;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT65), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT66), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT68), .Z(G217));
  NOR4_X1   g027(.A1(G221), .A2(G219), .A3(G220), .A4(G218), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G101), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(KEYINPUT69), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT69), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI211_X1 g042(.A(new_n463), .B(new_n465), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n462), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT3), .B(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(KEYINPUT70), .B1(new_n472), .B2(G125), .ZN(new_n473));
  OAI211_X1 g048(.A(KEYINPUT70), .B(G125), .C1(new_n466), .C2(new_n467), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n471), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT69), .B(G2105), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n470), .B1(new_n476), .B2(new_n478), .ZN(G160));
  OAI21_X1  g054(.A(G2104), .B1(new_n477), .B2(G112), .ZN(new_n480));
  NOR2_X1   g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT71), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n466), .A2(new_n467), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n484), .A2(new_n477), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n484), .A2(G2105), .ZN(new_n487));
  AOI211_X1 g062(.A(new_n483), .B(new_n486), .C1(G136), .C2(new_n487), .ZN(G162));
  NAND3_X1  g063(.A1(new_n472), .A2(G126), .A3(G2105), .ZN(new_n489));
  OR2_X1    g064(.A1(G102), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G114), .C2(new_n460), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  OAI21_X1  g068(.A(KEYINPUT4), .B1(new_n468), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n477), .A2(new_n472), .A3(new_n495), .A4(G138), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n492), .B1(new_n494), .B2(new_n496), .ZN(G164));
  INV_X1    g072(.A(KEYINPUT74), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(G543), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n501), .A2(KEYINPUT74), .A3(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n499), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT72), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G651), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n507), .A2(new_n509), .A3(KEYINPUT6), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT73), .B1(new_n506), .B2(KEYINPUT6), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT73), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n507), .A2(new_n509), .A3(new_n514), .A4(KEYINPUT6), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n505), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n501), .B1(new_n513), .B2(new_n515), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n516), .A2(G88), .B1(new_n517), .B2(G50), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n500), .A2(new_n502), .B1(new_n499), .B2(G543), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n519), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT72), .B(G651), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n518), .A2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  NAND2_X1  g099(.A1(new_n513), .A2(new_n515), .ZN(new_n525));
  XOR2_X1   g100(.A(KEYINPUT76), .B(G89), .Z(new_n526));
  NAND3_X1  g101(.A1(new_n525), .A2(new_n519), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(KEYINPUT75), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT75), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n530), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT7), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n529), .A2(new_n534), .A3(new_n531), .ZN(new_n535));
  AND2_X1   g110(.A1(G63), .A2(G651), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n533), .A2(new_n535), .B1(new_n519), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n511), .B1(new_n521), .B2(KEYINPUT6), .ZN(new_n538));
  AND4_X1   g113(.A1(new_n514), .A2(new_n507), .A3(new_n509), .A4(KEYINPUT6), .ZN(new_n539));
  OAI211_X1 g114(.A(G51), .B(G543), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n527), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(KEYINPUT77), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT77), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n527), .A2(new_n537), .A3(new_n540), .A4(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n544), .ZN(G168));
  NAND2_X1  g120(.A1(G77), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G64), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n505), .B2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n521), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n517), .A2(G52), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n525), .A2(G90), .A3(new_n519), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  NAND2_X1  g129(.A1(G68), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G56), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n505), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(new_n549), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n517), .A2(G43), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n525), .A2(G81), .A3(new_n519), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(G188));
  NAND2_X1  g142(.A1(G53), .A2(G543), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n568), .B1(new_n513), .B2(new_n515), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT78), .ZN(new_n570));
  OAI21_X1  g145(.A(KEYINPUT9), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AOI211_X1 g146(.A(KEYINPUT78), .B(new_n568), .C1(new_n513), .C2(new_n515), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT79), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT9), .ZN(new_n574));
  INV_X1    g149(.A(new_n568), .ZN(new_n575));
  OAI211_X1 g150(.A(new_n574), .B(new_n575), .C1(new_n538), .C2(new_n539), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n576), .A2(KEYINPUT80), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT80), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n578), .B1(new_n569), .B2(new_n574), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n538), .A2(new_n539), .ZN(new_n581));
  OAI21_X1  g156(.A(KEYINPUT78), .B1(new_n581), .B2(new_n568), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n569), .A2(new_n570), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .A4(KEYINPUT9), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n573), .A2(new_n580), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(G78), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G65), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n505), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n516), .A2(G91), .B1(new_n589), .B2(G651), .ZN(new_n590));
  AND3_X1   g165(.A1(new_n586), .A2(KEYINPUT81), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(KEYINPUT81), .B1(new_n586), .B2(new_n590), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n591), .A2(new_n592), .ZN(G299));
  INV_X1    g168(.A(G168), .ZN(G286));
  NAND2_X1  g169(.A1(new_n516), .A2(G87), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n517), .A2(G49), .ZN(new_n596));
  OAI21_X1  g171(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(G288));
  NAND3_X1  g173(.A1(new_n525), .A2(G48), .A3(G543), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n599), .B(KEYINPUT82), .ZN(new_n600));
  NAND2_X1  g175(.A1(G73), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G61), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n505), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n516), .A2(G86), .B1(new_n603), .B2(new_n549), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n600), .A2(new_n604), .ZN(G305));
  AOI22_X1  g180(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n606), .A2(new_n521), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n517), .A2(G47), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n516), .A2(G85), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(G290));
  NAND2_X1  g185(.A1(G301), .A2(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n516), .A2(G92), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT10), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n612), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(G79), .A2(G543), .ZN(new_n615));
  INV_X1    g190(.A(G66), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n505), .B2(new_n616), .ZN(new_n617));
  AOI22_X1  g192(.A1(G651), .A2(new_n617), .B1(new_n517), .B2(G54), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n611), .B1(new_n620), .B2(G868), .ZN(G284));
  OAI21_X1  g196(.A(new_n611), .B1(new_n620), .B2(G868), .ZN(G321));
  INV_X1    g197(.A(G868), .ZN(new_n623));
  NOR2_X1   g198(.A1(G168), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT83), .ZN(new_n625));
  INV_X1    g200(.A(G299), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(G868), .ZN(G297));
  OAI21_X1  g202(.A(new_n625), .B1(new_n626), .B2(G868), .ZN(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n620), .B1(new_n629), .B2(G860), .ZN(G148));
  NAND2_X1  g205(.A1(new_n561), .A2(new_n623), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n619), .A2(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(new_n632), .B2(new_n623), .ZN(G323));
  XOR2_X1   g208(.A(KEYINPUT84), .B(KEYINPUT11), .Z(new_n634));
  XNOR2_X1  g209(.A(G323), .B(new_n634), .ZN(G282));
  NAND2_X1  g210(.A1(new_n472), .A2(new_n461), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  INV_X1    g213(.A(G2100), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  AOI22_X1  g216(.A1(G123), .A2(new_n485), .B1(new_n487), .B2(G135), .ZN(new_n642));
  OAI221_X1 g217(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n477), .C2(G111), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(G2096), .Z(new_n645));
  NAND3_X1  g220(.A1(new_n640), .A2(new_n641), .A3(new_n645), .ZN(G156));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT85), .B(G2438), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2427), .B(G2430), .Z(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(KEYINPUT14), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n653), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  AND3_X1   g236(.A1(new_n660), .A2(G14), .A3(new_n661), .ZN(G401));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  NAND3_X1  g241(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT18), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT86), .B(KEYINPUT17), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n663), .B(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n666), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n670), .A2(new_n665), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n671), .B1(new_n664), .B2(new_n665), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n670), .B2(new_n665), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n668), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2096), .B(G2100), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G227));
  XNOR2_X1  g252(.A(G1971), .B(G1976), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1956), .B(G2474), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1961), .B(G1966), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT20), .ZN(new_n685));
  INV_X1    g260(.A(new_n680), .ZN(new_n686));
  INV_X1    g261(.A(new_n683), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n681), .A2(new_n682), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  OAI211_X1 g264(.A(new_n685), .B(new_n689), .C1(new_n686), .C2(new_n688), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1981), .B(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(G229));
  INV_X1    g271(.A(G29), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G25), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n485), .A2(G119), .ZN(new_n699));
  OAI221_X1 g274(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n477), .C2(G107), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n487), .A2(G131), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n698), .B1(new_n703), .B2(new_n697), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT35), .B(G1991), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G24), .ZN(new_n708));
  INV_X1    g283(.A(G290), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(new_n707), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT88), .B(G1986), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  MUX2_X1   g287(.A(G6), .B(G305), .S(G16), .Z(new_n713));
  XOR2_X1   g288(.A(KEYINPUT32), .B(G1981), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n707), .A2(G22), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G166), .B2(new_n707), .ZN(new_n717));
  INV_X1    g292(.A(G1971), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n707), .A2(G23), .ZN(new_n720));
  INV_X1    g295(.A(G288), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(new_n707), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT33), .B(G1976), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n715), .A2(new_n719), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT89), .B(KEYINPUT34), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n706), .B(new_n712), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n726), .B2(new_n725), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT36), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n707), .A2(G20), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT23), .Z(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G299), .B2(G16), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G1956), .ZN(new_n734));
  OAI21_X1  g309(.A(KEYINPUT92), .B1(G16), .B2(G21), .ZN(new_n735));
  NAND2_X1  g310(.A1(G168), .A2(G16), .ZN(new_n736));
  MUX2_X1   g311(.A(KEYINPUT92), .B(new_n735), .S(new_n736), .Z(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G1966), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n707), .A2(G19), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n562), .B2(new_n707), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n707), .A2(G5), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G171), .B2(new_n707), .ZN(new_n742));
  AOI22_X1  g317(.A1(G1341), .A2(new_n740), .B1(new_n742), .B2(G1961), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G1341), .B2(new_n740), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT30), .B(G28), .ZN(new_n745));
  OR2_X1    g320(.A1(KEYINPUT31), .A2(G11), .ZN(new_n746));
  NAND2_X1  g321(.A1(KEYINPUT31), .A2(G11), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n745), .A2(new_n697), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n485), .A2(G129), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n487), .A2(G141), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n461), .A2(G105), .ZN(new_n751));
  NAND3_X1  g326(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT26), .Z(new_n753));
  NAND4_X1  g328(.A1(new_n749), .A2(new_n750), .A3(new_n751), .A4(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n755), .A2(new_n697), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n697), .B2(G32), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT27), .B(G1996), .ZN(new_n758));
  OAI221_X1 g333(.A(new_n748), .B1(new_n697), .B2(new_n644), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n757), .B2(new_n758), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n697), .A2(G26), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  AOI22_X1  g338(.A1(G128), .A2(new_n485), .B1(new_n487), .B2(G140), .ZN(new_n764));
  OAI221_X1 g339(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n477), .C2(G116), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n763), .B1(new_n766), .B2(G29), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G2067), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n697), .A2(G27), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G164), .B2(new_n697), .ZN(new_n770));
  INV_X1    g345(.A(G2078), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n477), .A2(G103), .A3(G2104), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT91), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT25), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n774), .A2(new_n775), .ZN(new_n777));
  NAND2_X1  g352(.A1(G115), .A2(G2104), .ZN(new_n778));
  INV_X1    g353(.A(G127), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n778), .B1(new_n484), .B2(new_n779), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n780), .A2(new_n478), .B1(new_n487), .B2(G139), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n776), .A2(new_n777), .A3(new_n781), .ZN(new_n782));
  MUX2_X1   g357(.A(G33), .B(new_n782), .S(G29), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(G2072), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n760), .A2(new_n768), .A3(new_n772), .A4(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(G29), .A2(G35), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G162), .B2(G29), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT29), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G2090), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n742), .A2(G1961), .ZN(new_n790));
  OR4_X1    g365(.A1(new_n744), .A2(new_n785), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(G4), .A2(G16), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n620), .B2(G16), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n793), .A2(G1348), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n793), .A2(G1348), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n783), .A2(G2072), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT24), .ZN(new_n797));
  INV_X1    g372(.A(G34), .ZN(new_n798));
  AOI21_X1  g373(.A(G29), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n797), .B2(new_n798), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G160), .B2(new_n697), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n796), .B1(G2084), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G2084), .B2(new_n801), .ZN(new_n803));
  NOR4_X1   g378(.A1(new_n791), .A2(new_n794), .A3(new_n795), .A4(new_n803), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n730), .A2(new_n734), .A3(new_n738), .A4(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT93), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(G311));
  XNOR2_X1  g382(.A(new_n805), .B(KEYINPUT94), .ZN(G150));
  NAND2_X1  g383(.A1(G80), .A2(G543), .ZN(new_n809));
  INV_X1    g384(.A(G67), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n505), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(new_n549), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT95), .B(G55), .Z(new_n813));
  NAND2_X1  g388(.A1(new_n517), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n525), .A2(G93), .A3(new_n519), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n812), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(G860), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT37), .Z(new_n818));
  NOR2_X1   g393(.A1(new_n619), .A2(new_n629), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT38), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n516), .A2(G93), .B1(new_n811), .B2(new_n549), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n516), .A2(G81), .B1(new_n517), .B2(G43), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n821), .A2(new_n822), .A3(new_n558), .A4(new_n814), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n561), .A2(new_n816), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n820), .B(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT39), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT96), .ZN(new_n829));
  INV_X1    g404(.A(G860), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n826), .B2(new_n827), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n818), .B1(new_n829), .B2(new_n831), .ZN(G145));
  XNOR2_X1  g407(.A(G162), .B(G160), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT97), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(new_n644), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n702), .B(KEYINPUT99), .Z(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n637), .ZN(new_n838));
  AOI22_X1  g413(.A1(G130), .A2(new_n485), .B1(new_n487), .B2(G142), .ZN(new_n839));
  OAI221_X1 g414(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n477), .C2(G118), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n838), .B(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n766), .B(G164), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n754), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n782), .A2(KEYINPUT98), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n782), .B(KEYINPUT98), .Z(new_n847));
  OAI21_X1  g422(.A(new_n846), .B1(new_n844), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n842), .A2(new_n848), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n849), .A2(KEYINPUT100), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(KEYINPUT100), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n842), .A2(new_n848), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n836), .A2(new_n850), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(G37), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n852), .A2(new_n849), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n853), .B(new_n854), .C1(new_n836), .C2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT101), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT40), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(G395));
  NAND2_X1  g434(.A1(new_n816), .A2(new_n623), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n619), .B1(new_n591), .B2(new_n592), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n586), .A2(new_n590), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT81), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n586), .A2(KEYINPUT81), .A3(new_n590), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n864), .A2(new_n865), .A3(new_n620), .ZN(new_n866));
  AND3_X1   g441(.A1(new_n861), .A2(new_n866), .A3(KEYINPUT41), .ZN(new_n867));
  AOI21_X1  g442(.A(KEYINPUT41), .B1(new_n861), .B2(new_n866), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n825), .B(KEYINPUT102), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n632), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n861), .A2(new_n866), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n872), .B1(new_n873), .B2(new_n871), .ZN(new_n874));
  XNOR2_X1  g449(.A(G303), .B(G288), .ZN(new_n875));
  AOI21_X1  g450(.A(G290), .B1(new_n600), .B2(new_n604), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n600), .A2(new_n604), .A3(G290), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n875), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n875), .B1(new_n877), .B2(new_n878), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n882), .A2(KEYINPUT103), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT42), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n874), .B(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n860), .B1(new_n885), .B2(new_n623), .ZN(G295));
  OAI21_X1  g461(.A(new_n860), .B1(new_n885), .B2(new_n623), .ZN(G331));
  NAND3_X1  g462(.A1(G171), .A2(new_n542), .A3(new_n544), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(G171), .B1(new_n544), .B2(new_n542), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n825), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT105), .ZN(new_n892));
  NAND2_X1  g467(.A1(G168), .A2(G301), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n823), .A2(new_n824), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n893), .A2(new_n894), .A3(new_n888), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n891), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n893), .A2(new_n894), .A3(KEYINPUT105), .A4(new_n888), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT41), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n873), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n861), .A2(new_n866), .A3(KEYINPUT41), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n891), .A2(new_n895), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n873), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n881), .B1(new_n902), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n903), .B1(new_n867), .B2(new_n868), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n881), .B1(new_n898), .B2(new_n873), .ZN(new_n909));
  AOI21_X1  g484(.A(G37), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n911), .A2(KEYINPUT43), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n898), .A2(new_n873), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n908), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n881), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n913), .B1(new_n916), .B2(new_n910), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n912), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT109), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n916), .A2(new_n910), .A3(new_n913), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n916), .A2(new_n910), .A3(KEYINPUT106), .A4(new_n913), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n923), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n913), .B1(new_n911), .B2(KEYINPUT107), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n907), .A2(new_n910), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT108), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n904), .B1(new_n900), .B2(new_n901), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n914), .A2(new_n882), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n854), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n896), .A2(new_n897), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(new_n867), .B2(new_n868), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n882), .B1(new_n937), .B2(new_n905), .ZN(new_n938));
  OAI21_X1  g513(.A(KEYINPUT107), .B1(new_n935), .B2(new_n938), .ZN(new_n939));
  AND4_X1   g514(.A1(KEYINPUT108), .A2(new_n939), .A3(KEYINPUT43), .A4(new_n931), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n922), .B(new_n928), .C1(new_n932), .C2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n939), .A2(KEYINPUT43), .A3(new_n931), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT108), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n939), .A2(new_n931), .A3(KEYINPUT108), .A4(KEYINPUT43), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n922), .B1(new_n947), .B2(new_n928), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n921), .B1(new_n942), .B2(new_n948), .ZN(G397));
  INV_X1    g524(.A(new_n470), .ZN(new_n950));
  OAI21_X1  g525(.A(G125), .B1(new_n466), .B2(new_n467), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT70), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AOI22_X1  g528(.A1(new_n953), .A2(new_n474), .B1(G113), .B2(G2104), .ZN(new_n954));
  OAI211_X1 g529(.A(G40), .B(new_n950), .C1(new_n954), .C2(new_n477), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT111), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n476), .A2(new_n478), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT111), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n957), .A2(new_n958), .A3(G40), .A4(new_n950), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(KEYINPUT110), .B(G1384), .ZN(new_n961));
  NOR2_X1   g536(.A1(G164), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n962), .A2(KEYINPUT45), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G1996), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  XOR2_X1   g542(.A(new_n967), .B(KEYINPUT112), .Z(new_n968));
  OR2_X1    g543(.A1(new_n968), .A2(new_n754), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n766), .A2(G2067), .ZN(new_n970));
  INV_X1    g545(.A(G2067), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n764), .A2(new_n971), .A3(new_n765), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n973), .B1(new_n966), .B2(new_n755), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n964), .A2(new_n974), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n969), .A2(new_n705), .A3(new_n703), .A4(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n965), .B1(new_n976), .B2(new_n972), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n968), .B(KEYINPUT46), .ZN(new_n978));
  INV_X1    g553(.A(new_n973), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n964), .B1(new_n754), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  XOR2_X1   g556(.A(new_n981), .B(KEYINPUT47), .Z(new_n982));
  XNOR2_X1  g557(.A(new_n702), .B(new_n705), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n969), .B(new_n975), .C1(new_n965), .C2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n965), .A2(G1986), .A3(G290), .ZN(new_n986));
  XNOR2_X1  g561(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n986), .B(new_n987), .ZN(new_n988));
  AOI211_X1 g563(.A(new_n977), .B(new_n982), .C1(new_n985), .C2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n494), .A2(new_n496), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n990), .A2(new_n489), .A3(new_n491), .ZN(new_n991));
  INV_X1    g566(.A(G1384), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n994));
  AOI22_X1  g569(.A1(new_n956), .A2(new_n959), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n962), .A2(KEYINPUT45), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n718), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n993), .A2(KEYINPUT50), .ZN(new_n999));
  OR3_X1    g574(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n960), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n998), .B1(G2090), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(G303), .A2(G8), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1003), .B1(KEYINPUT113), .B2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g580(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1005), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1002), .A2(G8), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G8), .ZN(new_n1009));
  NOR2_X1   g584(.A1(G164), .A2(G1384), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1009), .B1(new_n960), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G1976), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1011), .B1(new_n1012), .B2(G288), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n721), .A2(G1976), .ZN(new_n1014));
  OR3_X1    g589(.A1(new_n1013), .A2(KEYINPUT52), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(KEYINPUT52), .ZN(new_n1016));
  NAND2_X1  g591(.A1(G305), .A2(G1981), .ZN(new_n1017));
  INV_X1    g592(.A(G1981), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n600), .A2(new_n1018), .A3(new_n604), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT49), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1017), .A2(KEYINPUT49), .A3(new_n1019), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(new_n1011), .A3(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1008), .A2(new_n1015), .A3(new_n1016), .A4(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT63), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1002), .A2(G8), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1007), .B1(new_n1028), .B2(KEYINPUT117), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1029), .B1(KEYINPUT117), .B2(new_n1028), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1001), .A2(G2084), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n1032));
  AOI22_X1  g607(.A1(new_n995), .A2(new_n1032), .B1(KEYINPUT45), .B2(new_n1010), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n958), .B1(G160), .B2(G40), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n955), .A2(KEYINPUT111), .ZN(new_n1035));
  OAI22_X1  g610(.A1(new_n1034), .A2(new_n1035), .B1(KEYINPUT45), .B2(new_n1010), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT116), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1033), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G1966), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1031), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1040), .A2(new_n1009), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(G168), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1027), .A2(new_n1030), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1000), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n956), .A2(new_n959), .B1(new_n993), .B2(KEYINPUT50), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1045), .B1(new_n1046), .B2(KEYINPUT115), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n960), .A2(new_n999), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT115), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(G2090), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1047), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n998), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1007), .B1(new_n1053), .B2(G8), .ZN(new_n1054));
  NOR3_X1   g629(.A1(new_n1042), .A2(new_n1025), .A3(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1044), .B1(new_n1055), .B2(KEYINPUT63), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1015), .A2(new_n1016), .A3(new_n1024), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1057), .A2(new_n1008), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1024), .A2(new_n1012), .A3(new_n721), .ZN(new_n1059));
  XOR2_X1   g634(.A(new_n1019), .B(KEYINPUT114), .Z(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1058), .B1(new_n1011), .B2(new_n1061), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n995), .A2(new_n996), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT53), .B1(new_n1063), .B2(new_n771), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1001), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1065), .A2(G1961), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1033), .A2(new_n1037), .A3(KEYINPUT53), .A4(new_n771), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1069), .A2(G301), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1041), .A2(G286), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n1073));
  NAND2_X1  g648(.A1(KEYINPUT121), .A2(G8), .ZN(new_n1074));
  AOI211_X1 g649(.A(new_n1073), .B(new_n1074), .C1(new_n1040), .C2(G168), .ZN(new_n1075));
  OAI22_X1  g650(.A1(new_n1036), .A2(KEYINPUT116), .B1(new_n994), .B2(new_n993), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n995), .A2(new_n1032), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1039), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1031), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1078), .A2(G168), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1074), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT51), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1072), .B1(new_n1075), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1071), .B1(new_n1083), .B2(KEYINPUT62), .ZN(new_n1084));
  AOI211_X1 g659(.A(G286), .B(new_n1031), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1073), .B1(new_n1085), .B2(new_n1074), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1080), .A2(KEYINPUT51), .A3(new_n1081), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT62), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1088), .A2(new_n1089), .A3(new_n1072), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT61), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT120), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT57), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1093), .B1(new_n586), .B2(new_n590), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n586), .A2(new_n1093), .A3(new_n590), .ZN(new_n1095));
  AOI21_X1  g670(.A(G1956), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT56), .B(G2072), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n995), .A2(new_n996), .A3(new_n1097), .ZN(new_n1098));
  OAI221_X1 g673(.A(new_n1092), .B1(new_n1094), .B2(new_n1095), .C1(new_n1096), .C2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G1956), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n960), .A2(KEYINPUT115), .A3(new_n999), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n1000), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1046), .A2(KEYINPUT115), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1100), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1095), .A2(new_n1094), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1098), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT120), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1105), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1091), .B(new_n1099), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n960), .A2(new_n1010), .ZN(new_n1112));
  XOR2_X1   g687(.A(KEYINPUT58), .B(G1341), .Z(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n995), .A2(new_n966), .A3(new_n996), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1111), .B1(new_n1116), .B2(new_n562), .ZN(new_n1117));
  AOI211_X1 g692(.A(KEYINPUT59), .B(new_n561), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT60), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1112), .A2(G2067), .ZN(new_n1121));
  AOI21_X1  g696(.A(G1348), .B1(new_n1046), .B2(new_n1000), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n620), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n960), .A2(new_n971), .A3(new_n1010), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n619), .B(new_n1124), .C1(new_n1065), .C2(G1348), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1120), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  NOR4_X1   g701(.A1(new_n1121), .A2(new_n1122), .A3(KEYINPUT60), .A4(new_n619), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1119), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT118), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1129), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1104), .A2(KEYINPUT118), .A3(new_n1106), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1094), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT119), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n586), .A2(new_n1093), .A3(new_n590), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT119), .B1(new_n1095), .B2(new_n1094), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1130), .A2(new_n1131), .A3(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1091), .B1(new_n1139), .B2(new_n1105), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1110), .A2(new_n1128), .A3(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1138), .A2(new_n1123), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(new_n1107), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  XOR2_X1   g720(.A(G301), .B(KEYINPUT54), .Z(new_n1146));
  NAND4_X1  g721(.A1(new_n950), .A2(KEYINPUT53), .A3(G40), .A4(new_n771), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1147), .B1(new_n962), .B2(KEYINPUT45), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n477), .B1(new_n476), .B2(KEYINPUT122), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1149), .B1(KEYINPUT122), .B2(new_n476), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1148), .B(new_n1150), .C1(KEYINPUT45), .C2(new_n962), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1146), .B1(new_n1151), .B2(KEYINPUT123), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1152), .B1(KEYINPUT123), .B2(new_n1151), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1067), .A2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1154), .B1(new_n1069), .B2(new_n1146), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1155), .B1(new_n1088), .B2(new_n1072), .ZN(new_n1156));
  AOI22_X1  g731(.A1(new_n1084), .A2(new_n1090), .B1(new_n1145), .B2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1025), .A2(new_n1054), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n1158), .B(KEYINPUT124), .ZN(new_n1159));
  OAI211_X1 g734(.A(new_n1056), .B(new_n1062), .C1(new_n1157), .C2(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g735(.A(G290), .B(G1986), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n984), .B1(new_n964), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(KEYINPUT125), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1145), .A2(new_n1156), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1083), .A2(KEYINPUT62), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1165), .A2(new_n1090), .A3(new_n1070), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1159), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1056), .A2(new_n1062), .ZN(new_n1168));
  OAI211_X1 g743(.A(KEYINPUT125), .B(new_n1162), .C1(new_n1167), .C2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n989), .B1(new_n1163), .B2(new_n1170), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g746(.A(G319), .ZN(new_n1173));
  OR3_X1    g747(.A1(G401), .A2(new_n1173), .A3(G227), .ZN(new_n1174));
  NOR4_X1   g748(.A1(new_n857), .A2(new_n918), .A3(G229), .A4(new_n1174), .ZN(G308));
  NOR3_X1   g749(.A1(new_n857), .A2(G229), .A3(new_n1174), .ZN(new_n1176));
  NAND2_X1  g750(.A1(new_n1176), .A2(new_n919), .ZN(G225));
endmodule


