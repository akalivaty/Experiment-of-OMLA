//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G143), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(new_n188), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT0), .B(G128), .ZN(new_n192));
  OAI21_X1  g006(.A(KEYINPUT66), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT11), .ZN(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(G137), .ZN(new_n196));
  INV_X1    g010(.A(G137), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT11), .A3(G134), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(G137), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n196), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G131), .ZN(new_n201));
  INV_X1    g015(.A(G131), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n196), .A2(new_n198), .A3(new_n202), .A4(new_n199), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n192), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT66), .ZN(new_n206));
  OR2_X1    g020(.A1(KEYINPUT65), .A2(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(KEYINPUT65), .A2(G143), .ZN(new_n208));
  AOI21_X1  g022(.A(G146), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n205), .B(new_n206), .C1(new_n209), .C2(new_n189), .ZN(new_n210));
  AND2_X1   g024(.A1(KEYINPUT0), .A2(G128), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n188), .A2(G143), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n211), .B(new_n212), .C1(new_n190), .C2(new_n188), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n193), .A2(new_n204), .A3(new_n210), .A4(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G128), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(KEYINPUT1), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n212), .B(new_n216), .C1(new_n190), .C2(new_n188), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n215), .B1(new_n212), .B2(KEYINPUT1), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n217), .B1(new_n191), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n197), .A2(KEYINPUT67), .A3(G134), .ZN(new_n220));
  INV_X1    g034(.A(new_n199), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n222), .B1(new_n195), .B2(G137), .ZN(new_n223));
  OAI211_X1 g037(.A(G131), .B(new_n220), .C1(new_n221), .C2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n219), .A2(new_n203), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n214), .A2(new_n225), .ZN(new_n226));
  XOR2_X1   g040(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT68), .ZN(new_n229));
  INV_X1    g043(.A(G119), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT69), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G119), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n231), .A2(new_n233), .A3(G116), .ZN(new_n234));
  INV_X1    g048(.A(G116), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G119), .ZN(new_n236));
  INV_X1    g050(.A(G113), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT2), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT2), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G113), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  AND3_X1   g055(.A1(new_n234), .A2(new_n236), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n241), .B1(new_n234), .B2(new_n236), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n214), .A2(new_n225), .A3(KEYINPUT30), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n226), .A2(new_n247), .A3(new_n227), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n229), .A2(new_n245), .A3(new_n246), .A4(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT31), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n214), .A2(new_n225), .A3(new_n244), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT70), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  XOR2_X1   g067(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n254));
  INV_X1    g068(.A(G237), .ZN(new_n255));
  INV_X1    g069(.A(G953), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n255), .A2(new_n256), .A3(G210), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n254), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT26), .B(G101), .ZN(new_n259));
  XOR2_X1   g073(.A(new_n258), .B(new_n259), .Z(new_n260));
  NAND4_X1  g074(.A1(new_n214), .A2(new_n225), .A3(new_n244), .A4(KEYINPUT70), .ZN(new_n261));
  AND3_X1   g075(.A1(new_n253), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n249), .A2(new_n250), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT28), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n251), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n226), .A2(new_n245), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n253), .A2(new_n261), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n266), .B1(new_n268), .B2(KEYINPUT28), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n263), .B1(new_n260), .B2(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n250), .B1(new_n249), .B2(new_n262), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n187), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT32), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n268), .A2(KEYINPUT28), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n260), .B1(new_n276), .B2(new_n265), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n249), .A2(new_n262), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT31), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n278), .A2(new_n280), .A3(new_n263), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(KEYINPUT72), .A3(new_n187), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n274), .A2(new_n275), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n187), .ZN(new_n284));
  AND3_X1   g098(.A1(new_n249), .A2(new_n250), .A3(new_n262), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n285), .A2(new_n277), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n284), .B1(new_n286), .B2(new_n280), .ZN(new_n287));
  INV_X1    g101(.A(G902), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n269), .A2(KEYINPUT29), .A3(new_n260), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n276), .A2(new_n260), .A3(new_n265), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT29), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AND2_X1   g106(.A1(new_n253), .A2(new_n261), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n260), .B1(new_n249), .B2(new_n293), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n288), .B(new_n289), .C1(new_n292), .C2(new_n294), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n287), .A2(KEYINPUT32), .B1(new_n295), .B2(G472), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n283), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n256), .A2(G221), .A3(G234), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n298), .B(KEYINPUT77), .ZN(new_n299));
  XNOR2_X1  g113(.A(KEYINPUT22), .B(G137), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n299), .B(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G110), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT24), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT24), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G110), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT74), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n303), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n306), .B1(new_n303), .B2(new_n305), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n230), .A2(G128), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT69), .B(G119), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n310), .B1(new_n311), .B2(G128), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT76), .B1(new_n309), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT23), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n314), .B1(new_n311), .B2(G128), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n302), .B(new_n315), .C1(new_n312), .C2(new_n314), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n231), .A2(new_n233), .A3(G128), .ZN(new_n317));
  INV_X1    g131(.A(new_n310), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT76), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n319), .B(new_n320), .C1(new_n307), .C2(new_n308), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n313), .A2(new_n316), .A3(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT16), .ZN(new_n323));
  INV_X1    g137(.A(G140), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(new_n324), .A3(G125), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(G125), .ZN(new_n326));
  INV_X1    g140(.A(G125), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G140), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  OAI211_X1 g143(.A(G146), .B(new_n325), .C1(new_n329), .C2(new_n323), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(G125), .B(G140), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n331), .B1(new_n188), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n322), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT78), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n314), .B1(new_n317), .B2(new_n318), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n231), .A2(new_n233), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT23), .B1(new_n337), .B2(new_n215), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT75), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT75), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n340), .B(new_n315), .C1(new_n312), .C2(new_n314), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n339), .A2(new_n341), .A3(G110), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n325), .B1(new_n329), .B2(new_n323), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n188), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n344), .A2(new_n330), .B1(new_n309), .B2(new_n312), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  AND3_X1   g160(.A1(new_n334), .A2(new_n335), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n335), .B1(new_n334), .B2(new_n346), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n301), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n301), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n334), .A2(new_n346), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n350), .B1(new_n351), .B2(KEYINPUT78), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT79), .ZN(new_n354));
  XOR2_X1   g168(.A(KEYINPUT73), .B(G217), .Z(new_n355));
  AOI21_X1  g169(.A(new_n355), .B1(G234), .B2(new_n288), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n356), .A2(G902), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT79), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n349), .A2(new_n358), .A3(new_n352), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n354), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n356), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n349), .A2(new_n288), .A3(new_n352), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT25), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n349), .A2(KEYINPUT25), .A3(new_n288), .A4(new_n352), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n361), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n360), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(KEYINPUT9), .B(G234), .ZN(new_n368));
  OAI21_X1  g182(.A(G221), .B1(new_n368), .B2(G902), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G104), .ZN(new_n371));
  OAI21_X1  g185(.A(KEYINPUT3), .B1(new_n371), .B2(G107), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT3), .ZN(new_n373));
  INV_X1    g187(.A(G107), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n374), .A3(G104), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n371), .A2(G107), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n372), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT4), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n378), .A3(G101), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n193), .A2(new_n210), .A3(new_n213), .A4(new_n379), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n377), .A2(G101), .ZN(new_n381));
  INV_X1    g195(.A(G101), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n372), .A2(new_n375), .A3(new_n382), .A4(new_n376), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT4), .ZN(new_n384));
  OAI21_X1  g198(.A(KEYINPUT80), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n377), .A2(G101), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT80), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n386), .A2(new_n387), .A3(KEYINPUT4), .A4(new_n383), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n380), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT10), .ZN(new_n390));
  INV_X1    g204(.A(G143), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(G146), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT1), .ZN(new_n393));
  OAI21_X1  g207(.A(G128), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n394), .B1(new_n209), .B2(new_n189), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n390), .B1(new_n395), .B2(new_n217), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n371), .A2(G107), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n374), .A2(G104), .ZN(new_n398));
  OAI21_X1  g212(.A(G101), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n383), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n212), .B1(new_n190), .B2(new_n188), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n393), .B1(new_n190), .B2(new_n188), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n403), .B1(new_n404), .B2(new_n215), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n400), .B1(new_n405), .B2(new_n217), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n402), .B1(new_n406), .B2(KEYINPUT10), .ZN(new_n407));
  OAI21_X1  g221(.A(KEYINPUT81), .B1(new_n389), .B2(new_n407), .ZN(new_n408));
  AND2_X1   g222(.A1(KEYINPUT65), .A2(G143), .ZN(new_n409));
  NOR2_X1   g223(.A1(KEYINPUT65), .A2(G143), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n188), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n189), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n192), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n213), .B1(new_n413), .B2(new_n206), .ZN(new_n414));
  INV_X1    g228(.A(new_n210), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n384), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n387), .B1(new_n417), .B2(new_n386), .ZN(new_n418));
  INV_X1    g232(.A(new_n388), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n416), .B(new_n379), .C1(new_n418), .C2(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n215), .B1(new_n411), .B2(KEYINPUT1), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n409), .A2(new_n410), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n392), .B1(new_n422), .B2(G146), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n217), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n401), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n425), .A2(new_n390), .B1(new_n401), .B2(new_n396), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT81), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n420), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n408), .A2(new_n428), .A3(new_n204), .ZN(new_n429));
  INV_X1    g243(.A(new_n204), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n420), .A2(new_n426), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(G110), .B(G140), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n256), .A2(G227), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n433), .B(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT82), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n395), .A2(new_n400), .A3(new_n217), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n425), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(KEYINPUT12), .B1(new_n439), .B2(new_n204), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT12), .ZN(new_n441));
  AOI211_X1 g255(.A(new_n441), .B(new_n430), .C1(new_n425), .C2(new_n438), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n437), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n438), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n204), .B1(new_n406), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n441), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n439), .A2(KEYINPUT12), .A3(new_n204), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(KEYINPUT82), .A3(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n435), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n443), .A2(new_n448), .A3(new_n431), .A4(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT83), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n431), .A2(new_n449), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n453), .A2(KEYINPUT83), .A3(new_n448), .A4(new_n443), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n436), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(G469), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(new_n456), .A3(new_n288), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n453), .A2(new_n429), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n446), .A2(new_n447), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n449), .B1(new_n459), .B2(new_n431), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(G469), .B1(new_n461), .B2(G902), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n370), .B1(new_n457), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(G210), .B1(G237), .B2(G902), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(G110), .B(G122), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(KEYINPUT8), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n242), .A2(new_n400), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n234), .A2(KEYINPUT5), .A3(new_n236), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(KEYINPUT84), .B1(new_n234), .B2(KEYINPUT5), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT84), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT5), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n311), .A2(new_n473), .A3(new_n474), .A4(G116), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n472), .A2(new_n475), .A3(G113), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT86), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n471), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n472), .A2(new_n475), .A3(KEYINPUT86), .A4(G113), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n469), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n472), .A2(new_n470), .A3(G113), .A4(new_n475), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n234), .A2(new_n236), .A3(new_n241), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n401), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n467), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n379), .B1(new_n242), .B2(new_n243), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n486), .B1(new_n418), .B2(new_n419), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n468), .A2(new_n481), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(new_n466), .A3(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(G125), .B1(new_n414), .B2(new_n415), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n395), .A2(new_n327), .A3(new_n217), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n256), .A2(G224), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n493), .B(KEYINPUT85), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT7), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n484), .A2(new_n489), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n491), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n193), .A2(new_n210), .A3(new_n213), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n500), .B1(new_n501), .B2(G125), .ZN(new_n502));
  AOI21_X1  g316(.A(KEYINPUT87), .B1(new_n502), .B2(new_n496), .ZN(new_n503));
  AND4_X1   g317(.A1(KEYINPUT87), .A2(new_n490), .A3(new_n491), .A4(new_n496), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n288), .B1(new_n499), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n466), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n485), .B1(new_n385), .B2(new_n388), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n468), .A2(new_n481), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n489), .A2(new_n510), .A3(KEYINPUT6), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT6), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n512), .B(new_n507), .C1(new_n508), .C2(new_n509), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n490), .A2(new_n491), .A3(new_n494), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n494), .B1(new_n490), .B2(new_n491), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n511), .A2(new_n513), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n465), .B1(new_n506), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT87), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n519), .B1(new_n492), .B2(new_n497), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n502), .A2(KEYINPUT87), .A3(new_n496), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n522), .A2(new_n489), .A3(new_n484), .A4(new_n498), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n511), .A2(new_n513), .A3(new_n516), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n523), .A2(new_n524), .A3(new_n288), .A4(new_n464), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n518), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(G952), .ZN(new_n527));
  OR2_X1    g341(.A1(new_n527), .A2(KEYINPUT93), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(KEYINPUT93), .ZN(new_n529));
  AOI21_X1  g343(.A(G953), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(G234), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n530), .B1(new_n531), .B2(new_n255), .ZN(new_n532));
  XOR2_X1   g346(.A(new_n532), .B(KEYINPUT94), .Z(new_n533));
  OAI211_X1 g347(.A(G902), .B(G953), .C1(new_n531), .C2(new_n255), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n534), .B(KEYINPUT95), .ZN(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT21), .B(G898), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(G214), .B1(G237), .B2(G902), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n526), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(G214), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n542), .A2(G237), .A3(G953), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(KEYINPUT89), .A3(G143), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT89), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n255), .A2(new_n256), .A3(G214), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n545), .B1(new_n546), .B2(new_n391), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NOR3_X1   g362(.A1(new_n190), .A2(new_n543), .A3(KEYINPUT88), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT88), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n550), .B1(new_n422), .B2(new_n546), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n548), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(G131), .ZN(new_n553));
  OAI21_X1  g367(.A(KEYINPUT88), .B1(new_n190), .B2(new_n543), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n422), .A2(new_n550), .A3(new_n546), .ZN(new_n555));
  AOI22_X1  g369(.A1(new_n554), .A2(new_n555), .B1(new_n547), .B2(new_n544), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n202), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT17), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n553), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n344), .A2(new_n330), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n554), .A2(new_n555), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n202), .B1(new_n561), .B2(new_n548), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n560), .B1(new_n562), .B2(KEYINPUT17), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(G113), .B(G122), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(new_n371), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(KEYINPUT91), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n332), .B(G146), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT18), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n569), .A2(new_n202), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n568), .B1(new_n556), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n552), .A2(KEYINPUT18), .A3(G131), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT90), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n574), .B1(new_n572), .B2(new_n573), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n564), .B(new_n567), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n568), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n578), .B1(new_n552), .B2(new_n570), .ZN(new_n579));
  NOR3_X1   g393(.A1(new_n556), .A2(new_n569), .A3(new_n202), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT90), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n581), .A2(new_n582), .B1(new_n559), .B2(new_n563), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n577), .B1(new_n583), .B2(new_n566), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n288), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(G475), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n553), .A2(new_n557), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n332), .B(KEYINPUT19), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n331), .B1(new_n188), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n581), .A2(new_n582), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n577), .B1(new_n590), .B2(new_n566), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT20), .ZN(new_n592));
  NOR2_X1   g406(.A1(G475), .A2(G902), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n592), .B1(new_n591), .B2(new_n593), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n586), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(G122), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(G116), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n235), .A2(G122), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(G107), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n207), .A2(G128), .A3(new_n208), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n215), .A2(G143), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n602), .A2(new_n195), .A3(new_n603), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n602), .A2(KEYINPUT13), .A3(new_n603), .ZN(new_n605));
  OAI21_X1  g419(.A(G134), .B1(new_n602), .B2(KEYINPUT13), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n601), .B(new_n604), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n374), .B1(new_n598), .B2(KEYINPUT14), .ZN(new_n608));
  OR2_X1    g422(.A1(new_n608), .A2(new_n600), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n600), .ZN(new_n610));
  INV_X1    g424(.A(new_n604), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n195), .B1(new_n602), .B2(new_n603), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n609), .B(new_n610), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n355), .A2(G953), .A3(new_n368), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n607), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n614), .B1(new_n607), .B2(new_n613), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n288), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(G478), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(KEYINPUT15), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  OAI221_X1 g434(.A(new_n288), .B1(KEYINPUT15), .B2(new_n618), .C1(new_n615), .C2(new_n616), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT92), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n541), .A2(new_n596), .A3(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n297), .A2(new_n367), .A3(new_n463), .A4(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G101), .ZN(G3));
  NAND2_X1  g441(.A1(new_n457), .A2(new_n462), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n628), .A2(new_n367), .A3(new_n369), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n288), .B1(new_n270), .B2(new_n271), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(G472), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n274), .A2(new_n631), .A3(new_n282), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT96), .ZN(new_n634));
  INV_X1    g448(.A(new_n540), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n635), .B1(new_n518), .B2(new_n525), .ZN(new_n636));
  OR2_X1    g450(.A1(new_n615), .A2(new_n616), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n637), .A2(new_n618), .A3(new_n288), .ZN(new_n638));
  NAND2_X1  g452(.A1(G478), .A2(G902), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n637), .B(KEYINPUT33), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n638), .B(new_n639), .C1(new_n640), .C2(new_n618), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n636), .A2(new_n596), .A3(new_n539), .A4(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n634), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT34), .B(G104), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G6));
  OAI211_X1 g461(.A(new_n624), .B(new_n586), .C1(new_n595), .C2(new_n594), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n541), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n634), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT35), .B(G107), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G9));
  AND3_X1   g466(.A1(new_n274), .A2(new_n631), .A3(new_n282), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n364), .A2(new_n365), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n356), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n350), .A2(KEYINPUT36), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n351), .A2(KEYINPUT97), .ZN(new_n658));
  AOI22_X1  g472(.A1(new_n322), .A2(new_n333), .B1(new_n342), .B2(new_n345), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT97), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n657), .B1(new_n658), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n351), .A2(KEYINPUT97), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n659), .A2(new_n660), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n663), .A2(new_n664), .A3(new_n656), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(KEYINPUT98), .B1(new_n666), .B2(new_n357), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT98), .ZN(new_n668));
  INV_X1    g482(.A(new_n357), .ZN(new_n669));
  AOI211_X1 g483(.A(new_n668), .B(new_n669), .C1(new_n662), .C2(new_n665), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n655), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n653), .A2(new_n625), .A3(new_n463), .A4(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT37), .B(G110), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G12));
  INV_X1    g489(.A(new_n297), .ZN(new_n676));
  INV_X1    g490(.A(G900), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n535), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n533), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n648), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n680), .A2(new_n463), .A3(new_n636), .A4(new_n672), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(new_n215), .ZN(G30));
  XOR2_X1   g497(.A(new_n679), .B(KEYINPUT39), .Z(new_n684));
  NAND2_X1  g498(.A1(new_n463), .A2(new_n684), .ZN(new_n685));
  OR2_X1    g499(.A1(new_n685), .A2(KEYINPUT40), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n281), .A2(KEYINPUT32), .A3(new_n187), .ZN(new_n687));
  INV_X1    g501(.A(new_n260), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n688), .B1(new_n249), .B2(new_n293), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n288), .B1(new_n268), .B2(new_n260), .ZN(new_n690));
  OAI21_X1  g504(.A(G472), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n692), .A2(new_n283), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n685), .A2(KEYINPUT40), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT38), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n526), .B(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n596), .A2(new_n624), .A3(new_n540), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n697), .A2(new_n672), .A3(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n686), .A2(new_n694), .A3(new_n695), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n190), .ZN(G45));
  NAND2_X1  g515(.A1(new_n591), .A2(new_n593), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(KEYINPUT20), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n704));
  AOI22_X1  g518(.A1(new_n703), .A2(new_n704), .B1(G475), .B2(new_n585), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n705), .A2(new_n641), .A3(new_n679), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n463), .A2(new_n706), .A3(new_n636), .A4(new_n672), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n676), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(new_n188), .ZN(G48));
  AND3_X1   g523(.A1(new_n455), .A2(new_n456), .A3(new_n288), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n456), .B1(new_n455), .B2(new_n288), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n710), .A2(new_n711), .A3(new_n370), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n297), .A2(new_n367), .A3(new_n644), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT41), .B(G113), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G15));
  NAND4_X1  g529(.A1(new_n297), .A2(new_n367), .A3(new_n649), .A4(new_n712), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT99), .B(G116), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G18));
  NOR3_X1   g532(.A1(new_n596), .A2(new_n624), .A3(new_n538), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n672), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n720), .B1(new_n283), .B2(new_n296), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT100), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n722), .B1(new_n712), .B2(new_n636), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n455), .A2(new_n288), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(G469), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n725), .A2(new_n369), .A3(new_n457), .A4(new_n636), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(KEYINPUT100), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n721), .B1(new_n723), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(KEYINPUT101), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n712), .A2(new_n722), .A3(new_n636), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n726), .A2(KEYINPUT100), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT101), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n732), .A2(new_n733), .A3(new_n721), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n729), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G119), .ZN(G21));
  NAND2_X1  g550(.A1(new_n631), .A2(new_n272), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n354), .A2(new_n359), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n655), .B1(new_n738), .B2(new_n669), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n636), .A2(new_n596), .A3(new_n624), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n740), .A2(new_n539), .A3(new_n712), .A4(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G122), .ZN(G24));
  NAND4_X1  g557(.A1(new_n706), .A2(new_n272), .A3(new_n672), .A4(new_n631), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n744), .B1(new_n730), .B2(new_n731), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n327), .ZN(G27));
  NAND3_X1  g560(.A1(new_n518), .A2(new_n540), .A3(new_n525), .ZN(new_n747));
  AOI211_X1 g561(.A(new_n370), .B(new_n747), .C1(new_n457), .C2(new_n462), .ZN(new_n748));
  INV_X1    g562(.A(new_n679), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n596), .A2(new_n642), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n750), .A2(KEYINPUT42), .ZN(new_n751));
  AND4_X1   g565(.A1(new_n297), .A2(new_n748), .A3(new_n367), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n272), .A2(new_n275), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n292), .A2(new_n294), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n289), .A2(new_n288), .ZN(new_n755));
  OAI21_X1  g569(.A(G472), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n753), .A2(new_n756), .A3(new_n687), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT102), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n757), .A2(new_n758), .A3(new_n367), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n758), .B1(new_n757), .B2(new_n367), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n706), .B(new_n748), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n752), .B1(new_n761), .B2(KEYINPUT42), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G131), .ZN(G33));
  NAND4_X1  g577(.A1(new_n297), .A2(new_n748), .A3(new_n367), .A4(new_n680), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G134), .ZN(G36));
  NOR3_X1   g579(.A1(new_n366), .A2(new_n667), .A3(new_n670), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n653), .A2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT43), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n705), .A2(new_n768), .A3(new_n642), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT104), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n641), .B1(new_n596), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n705), .A2(KEYINPUT104), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n770), .B1(new_n774), .B2(KEYINPUT43), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n767), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT44), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT107), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n776), .A2(KEYINPUT107), .A3(new_n777), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n767), .A2(new_n775), .A3(KEYINPUT44), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT106), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n747), .B(KEYINPUT105), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n784), .B1(new_n783), .B2(new_n785), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n782), .A2(new_n786), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT108), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n461), .A2(KEYINPUT45), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT45), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n793), .B1(new_n458), .B2(new_n460), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n792), .A2(G469), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(G469), .A2(G902), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT46), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT103), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n795), .A2(KEYINPUT46), .A3(new_n796), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n800), .A2(new_n457), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n797), .A2(new_n798), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n799), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n369), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n684), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n782), .A2(KEYINPUT108), .A3(new_n786), .A4(new_n788), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n791), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G137), .ZN(G39));
  NOR4_X1   g624(.A1(new_n297), .A2(new_n750), .A3(new_n367), .A4(new_n747), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(KEYINPUT109), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT47), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n804), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n803), .A2(KEYINPUT47), .A3(new_n369), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n813), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G140), .ZN(G42));
  INV_X1    g633(.A(new_n697), .ZN(new_n820));
  OR4_X1    g634(.A1(new_n739), .A2(new_n774), .A3(new_n370), .A4(new_n635), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(KEYINPUT110), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n710), .A2(new_n711), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  AOI211_X1 g638(.A(new_n820), .B(new_n822), .C1(KEYINPUT49), .C2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(KEYINPUT49), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT111), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(KEYINPUT111), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n828), .B1(KEYINPUT110), .B2(new_n821), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n825), .A2(new_n693), .A3(new_n827), .A4(new_n829), .ZN(new_n830));
  AOI211_X1 g644(.A(new_n533), .B(new_n770), .C1(KEYINPUT43), .C2(new_n774), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(new_n740), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n824), .A2(new_n369), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n785), .B(new_n833), .C1(new_n817), .C2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n712), .A2(new_n635), .A3(new_n697), .ZN(new_n836));
  OR4_X1    g650(.A1(KEYINPUT116), .A2(new_n832), .A3(KEYINPUT50), .A4(new_n836), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n824), .A2(new_n370), .A3(new_n747), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n739), .A2(new_n533), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n838), .A2(new_n693), .A3(new_n839), .ZN(new_n840));
  OR3_X1    g654(.A1(new_n840), .A2(new_n596), .A3(new_n642), .ZN(new_n841));
  XOR2_X1   g655(.A(KEYINPUT116), .B(KEYINPUT50), .Z(new_n842));
  OAI21_X1  g656(.A(new_n842), .B1(new_n832), .B2(new_n836), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n831), .A2(new_n838), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n737), .A2(new_n766), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n841), .A2(new_n843), .A3(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n835), .A2(new_n837), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT51), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n848), .A2(KEYINPUT115), .A3(new_n849), .ZN(new_n850));
  OR2_X1    g664(.A1(new_n759), .A2(new_n760), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n844), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(KEYINPUT48), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n596), .A2(new_n642), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n530), .B1(new_n840), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n855), .B1(new_n732), .B2(new_n833), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n850), .A2(new_n853), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT54), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n681), .A2(new_n707), .B1(new_n283), .B2(new_n296), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n741), .A2(new_n463), .A3(new_n766), .A4(new_n749), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n693), .A2(new_n861), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n745), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n863), .A2(KEYINPUT114), .A3(KEYINPUT52), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT52), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n706), .B(new_n845), .C1(new_n723), .C2(new_n727), .ZN(new_n866));
  INV_X1    g680(.A(new_n862), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n463), .A2(new_n636), .A3(new_n672), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n868), .B(new_n297), .C1(new_n680), .C2(new_n706), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n866), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT114), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n865), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n864), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT112), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n586), .B(new_n622), .C1(new_n594), .C2(new_n595), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n874), .B1(new_n541), .B2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n875), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n877), .A2(KEYINPUT112), .A3(new_n539), .A4(new_n636), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n876), .A2(new_n878), .A3(new_n643), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n633), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n880), .A2(new_n713), .A3(new_n716), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n626), .A2(new_n742), .A3(new_n673), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n622), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n705), .A2(new_n884), .A3(new_n749), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n766), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n297), .A2(new_n748), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n764), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n845), .A2(new_n748), .A3(new_n706), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT113), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n845), .A2(new_n748), .A3(KEYINPUT113), .A4(new_n706), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n888), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n735), .A2(new_n883), .A3(new_n893), .A4(new_n762), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n859), .B1(new_n873), .B2(new_n894), .ZN(new_n895));
  AND4_X1   g709(.A1(new_n735), .A2(new_n883), .A3(new_n893), .A4(new_n762), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n745), .A2(new_n860), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT52), .B1(new_n897), .B2(new_n867), .ZN(new_n898));
  NOR4_X1   g712(.A1(new_n745), .A2(new_n860), .A3(new_n862), .A4(new_n865), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n896), .B(KEYINPUT53), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n858), .B1(new_n895), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(KEYINPUT52), .B1(new_n863), .B2(KEYINPUT114), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n870), .A2(new_n871), .A3(new_n865), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n904), .A2(new_n896), .A3(KEYINPUT53), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n898), .A2(new_n899), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n859), .B1(new_n906), .B2(new_n894), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n905), .A2(new_n858), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n849), .B1(new_n848), .B2(KEYINPUT115), .ZN(new_n909));
  NOR4_X1   g723(.A1(new_n857), .A2(new_n901), .A3(new_n908), .A4(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(G952), .A2(G953), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n830), .B1(new_n910), .B2(new_n911), .ZN(G75));
  NOR2_X1   g726(.A1(new_n256), .A2(G952), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n288), .B1(new_n905), .B2(new_n907), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT56), .B1(new_n915), .B2(G210), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n511), .A2(new_n513), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(new_n516), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT55), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n914), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n920), .B1(new_n916), .B2(new_n919), .ZN(G51));
  INV_X1    g735(.A(new_n795), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n915), .A2(new_n922), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT118), .Z(new_n924));
  XNOR2_X1  g738(.A(new_n455), .B(KEYINPUT117), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n905), .A2(new_n907), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(KEYINPUT54), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n905), .A2(new_n907), .A3(new_n858), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n796), .B(KEYINPUT57), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n925), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n913), .B1(new_n924), .B2(new_n932), .ZN(G54));
  AND2_X1   g747(.A1(KEYINPUT58), .A2(G475), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n915), .A2(new_n591), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n591), .B1(new_n915), .B2(new_n934), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n935), .A2(new_n936), .A3(new_n913), .ZN(G60));
  INV_X1    g751(.A(KEYINPUT120), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n639), .B(KEYINPUT59), .Z(new_n939));
  AOI21_X1  g753(.A(KEYINPUT53), .B1(new_n904), .B2(new_n896), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n906), .A2(new_n894), .A3(new_n859), .ZN(new_n941));
  OAI21_X1  g755(.A(KEYINPUT54), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n939), .B1(new_n942), .B2(new_n928), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n938), .B1(new_n943), .B2(new_n640), .ZN(new_n944));
  INV_X1    g758(.A(new_n640), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n945), .A2(new_n939), .ZN(new_n946));
  AOI21_X1  g760(.A(KEYINPUT119), .B1(new_n929), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n858), .B1(new_n905), .B2(new_n907), .ZN(new_n948));
  OAI211_X1 g762(.A(KEYINPUT119), .B(new_n946), .C1(new_n908), .C2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n944), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n939), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n952), .B1(new_n901), .B2(new_n908), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n953), .A2(KEYINPUT120), .A3(new_n945), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n914), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n951), .A2(new_n955), .ZN(G63));
  XNOR2_X1  g770(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n957));
  NAND2_X1  g771(.A1(G217), .A2(G902), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n957), .B(new_n958), .Z(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n905), .B2(new_n907), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n913), .B1(new_n962), .B2(new_n738), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n666), .B(KEYINPUT122), .Z(new_n964));
  AND3_X1   g778(.A1(new_n961), .A2(KEYINPUT123), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(KEYINPUT123), .B1(new_n961), .B2(new_n964), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n963), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT61), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n963), .B(KEYINPUT61), .C1(new_n965), .C2(new_n966), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(G66));
  INV_X1    g785(.A(G224), .ZN(new_n972));
  OAI21_X1  g786(.A(G953), .B1(new_n536), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n735), .A2(new_n883), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n973), .B1(new_n975), .B2(G953), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n917), .B1(G898), .B2(new_n256), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n976), .B(new_n977), .ZN(G69));
  INV_X1    g792(.A(KEYINPUT126), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n805), .A2(new_n684), .A3(new_n851), .A4(new_n741), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n815), .A2(new_n816), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n764), .B(new_n980), .C1(new_n981), .C2(new_n812), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT124), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n897), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(KEYINPUT124), .B1(new_n745), .B2(new_n860), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(new_n762), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n982), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n988), .A2(new_n809), .A3(new_n256), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n229), .A2(new_n246), .A3(new_n248), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(new_n588), .Z(new_n991));
  NAND2_X1  g805(.A1(G900), .A2(G953), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n979), .B1(new_n989), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n297), .A2(new_n367), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n854), .A2(new_n875), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  NOR4_X1   g811(.A1(new_n995), .A2(new_n997), .A3(new_n685), .A4(new_n747), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n998), .B1(new_n813), .B2(new_n817), .ZN(new_n999));
  INV_X1    g813(.A(new_n700), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n1000), .B1(new_n984), .B2(new_n985), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n1001), .A2(KEYINPUT62), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT62), .ZN(new_n1003));
  AOI211_X1 g817(.A(new_n1003), .B(new_n1000), .C1(new_n984), .C2(new_n985), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n999), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n808), .A2(new_n807), .ZN(new_n1006));
  INV_X1    g820(.A(new_n786), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n1007), .A2(new_n787), .ZN(new_n1008));
  AOI21_X1  g822(.A(KEYINPUT108), .B1(new_n1008), .B2(new_n782), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(KEYINPUT125), .B1(new_n1005), .B2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1001), .B(KEYINPUT62), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT125), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n1012), .A2(new_n809), .A3(new_n1013), .A4(new_n999), .ZN(new_n1014));
  AOI21_X1  g828(.A(G953), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n994), .B1(new_n1015), .B2(new_n991), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n256), .B1(G227), .B2(G900), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g832(.A(new_n1017), .ZN(new_n1019));
  OAI211_X1 g833(.A(new_n1019), .B(new_n994), .C1(new_n1015), .C2(new_n991), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1018), .A2(new_n1020), .ZN(G72));
  NAND3_X1  g835(.A1(new_n988), .A2(new_n809), .A3(new_n975), .ZN(new_n1022));
  NAND2_X1  g836(.A1(G472), .A2(G902), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n1023), .B(KEYINPUT63), .Z(new_n1024));
  NAND3_X1  g838(.A1(new_n1022), .A2(KEYINPUT127), .A3(new_n1024), .ZN(new_n1025));
  AND3_X1   g839(.A1(new_n249), .A2(new_n688), .A3(new_n293), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g841(.A(KEYINPUT127), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g843(.A(new_n689), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n1011), .A2(new_n975), .A3(new_n1014), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1030), .B1(new_n1031), .B2(new_n1024), .ZN(new_n1032));
  INV_X1    g846(.A(new_n1024), .ZN(new_n1033));
  NOR3_X1   g847(.A1(new_n1026), .A2(new_n689), .A3(new_n1033), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1034), .B1(new_n940), .B2(new_n941), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1035), .A2(new_n914), .ZN(new_n1036));
  NOR3_X1   g850(.A1(new_n1029), .A2(new_n1032), .A3(new_n1036), .ZN(G57));
endmodule


