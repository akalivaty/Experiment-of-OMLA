//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 0 1 0 0 0 1 0 0 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 0 0 0 0 1 1 1 1 1 1 1 0 1 0 1 0 1 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1261,
    new_n1262, new_n1263, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  INV_X1    g0012(.A(G58), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n207), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n221));
  INV_X1    g0021(.A(G226), .ZN(new_n222));
  INV_X1    g0022(.A(G116), .ZN(new_n223));
  INV_X1    g0023(.A(G270), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n221), .B1(new_n202), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n209), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n212), .B(new_n220), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n202), .A2(G68), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n214), .A2(G50), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n243), .B(new_n248), .Z(G351));
  NAND2_X1  g0049(.A1(G33), .A2(G41), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(KEYINPUT64), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT64), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n252), .A2(G33), .A3(G41), .ZN(new_n253));
  INV_X1    g0053(.A(new_n218), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n251), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G41), .ZN(new_n256));
  INV_X1    g0056(.A(G45), .ZN(new_n257));
  AOI21_X1  g0057(.A(G1), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n255), .A2(G274), .A3(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n258), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n255), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n259), .B1(new_n261), .B2(new_n222), .ZN(new_n262));
  OR2_X1    g0062(.A1(new_n262), .A2(KEYINPUT65), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT3), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(G1698), .B1(new_n266), .B2(new_n267), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n269), .A2(G77), .B1(new_n270), .B2(G222), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n268), .A2(G1698), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT66), .B(G223), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n254), .A2(new_n250), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n262), .A2(KEYINPUT65), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n263), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G179), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  XOR2_X1   g0082(.A(KEYINPUT8), .B(G58), .Z(new_n283));
  NOR2_X1   g0083(.A1(new_n265), .A2(G20), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G20), .A2(G33), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n283), .A2(new_n284), .B1(G150), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT67), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n286), .A2(new_n287), .B1(G20), .B2(new_n203), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n288), .B1(new_n287), .B2(new_n286), .ZN(new_n289));
  NAND3_X1  g0089(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n218), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G13), .ZN(new_n293));
  NOR3_X1   g0093(.A1(new_n293), .A2(new_n207), .A3(G1), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(new_n291), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n202), .B1(new_n206), .B2(G20), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n295), .A2(new_n296), .B1(new_n202), .B2(new_n294), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G169), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n279), .A2(new_n299), .ZN(new_n300));
  AND3_X1   g0100(.A1(new_n282), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT70), .ZN(new_n302));
  INV_X1    g0102(.A(new_n298), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n302), .B1(new_n303), .B2(KEYINPUT9), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT9), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n298), .A2(KEYINPUT70), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n280), .A2(G190), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n303), .A2(KEYINPUT9), .B1(G200), .B2(new_n279), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT10), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT10), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n307), .A2(new_n312), .A3(new_n308), .A4(new_n309), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n301), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n206), .A2(G20), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n283), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT8), .B(G58), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n317), .A2(new_n295), .B1(new_n294), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n291), .ZN(new_n321));
  NAND2_X1  g0121(.A1(G58), .A2(G68), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(G20), .B1(new_n323), .B2(new_n201), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT75), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n285), .A2(G159), .ZN(new_n327));
  OAI211_X1 g0127(.A(KEYINPUT75), .B(G20), .C1(new_n323), .C2(new_n201), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  AND2_X1   g0129(.A1(KEYINPUT3), .A2(G33), .ZN(new_n330));
  NOR2_X1   g0130(.A1(KEYINPUT3), .A2(G33), .ZN(new_n331));
  NOR3_X1   g0131(.A1(new_n330), .A2(new_n331), .A3(G20), .ZN(new_n332));
  OAI21_X1  g0132(.A(KEYINPUT74), .B1(new_n332), .B2(KEYINPUT7), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT7), .ZN(new_n334));
  NOR4_X1   g0134(.A1(new_n330), .A2(new_n331), .A3(new_n334), .A4(G20), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n266), .A2(new_n207), .A3(new_n267), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT74), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n337), .A2(new_n338), .A3(new_n334), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n333), .A2(new_n336), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n329), .B1(new_n340), .B2(G68), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n321), .B1(new_n341), .B2(KEYINPUT16), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT16), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n337), .A2(new_n334), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n335), .B1(KEYINPUT76), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT76), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n337), .A2(new_n346), .A3(new_n334), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n214), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n343), .B1(new_n348), .B2(new_n329), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n320), .B1(new_n342), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n259), .B1(new_n261), .B2(new_n233), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT77), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT77), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n259), .B(new_n353), .C1(new_n261), .C2(new_n233), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n222), .A2(G1698), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n268), .B(new_n356), .C1(G223), .C2(G1698), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G33), .A2(G87), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n275), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n359), .A2(G179), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  OR2_X1    g0161(.A1(new_n359), .A2(new_n351), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n299), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(KEYINPUT18), .B1(new_n350), .B2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n329), .ZN(new_n366));
  AND3_X1   g0166(.A1(new_n337), .A2(new_n338), .A3(new_n334), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n338), .B1(new_n337), .B2(new_n334), .ZN(new_n368));
  NOR3_X1   g0168(.A1(new_n367), .A2(new_n368), .A3(new_n335), .ZN(new_n369));
  OAI211_X1 g0169(.A(KEYINPUT16), .B(new_n366), .C1(new_n369), .C2(new_n214), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n291), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n344), .A2(KEYINPUT76), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n372), .A2(new_n347), .A3(new_n336), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(G68), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT16), .B1(new_n374), .B2(new_n366), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n319), .B1(new_n371), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT18), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n355), .A2(new_n360), .B1(new_n299), .B2(new_n362), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n365), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n359), .A2(G190), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n381), .A2(new_n352), .A3(new_n354), .ZN(new_n382));
  INV_X1    g0182(.A(G200), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(new_n359), .B2(new_n351), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n385), .B(new_n319), .C1(new_n371), .C2(new_n375), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT17), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n350), .A2(KEYINPUT17), .A3(new_n385), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n380), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n270), .A2(G232), .ZN(new_n392));
  INV_X1    g0192(.A(G107), .ZN(new_n393));
  INV_X1    g0193(.A(G238), .ZN(new_n394));
  OAI221_X1 g0194(.A(new_n392), .B1(new_n393), .B2(new_n268), .C1(new_n394), .C2(new_n272), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n276), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n255), .A2(G244), .A3(new_n260), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n396), .A2(new_n281), .A3(new_n259), .A4(new_n397), .ZN(new_n398));
  XOR2_X1   g0198(.A(new_n398), .B(KEYINPUT69), .Z(new_n399));
  NAND3_X1  g0199(.A1(new_n396), .A2(new_n259), .A3(new_n397), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n299), .ZN(new_n401));
  INV_X1    g0201(.A(new_n285), .ZN(new_n402));
  INV_X1    g0202(.A(G77), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n318), .A2(new_n402), .B1(new_n207), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g0204(.A(KEYINPUT15), .B(G87), .ZN(new_n405));
  INV_X1    g0205(.A(new_n284), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n291), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  XNOR2_X1  g0208(.A(new_n408), .B(KEYINPUT68), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n403), .B1(new_n206), .B2(G20), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n295), .A2(new_n410), .B1(new_n403), .B2(new_n294), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n401), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n399), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n412), .B1(G200), .B2(new_n400), .ZN(new_n416));
  INV_X1    g0216(.A(G190), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n416), .B1(new_n417), .B2(new_n400), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n314), .A2(new_n391), .A3(new_n415), .A4(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(G33), .A2(G97), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n233), .A2(G1698), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(G226), .B2(G1698), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n420), .B1(new_n422), .B2(new_n269), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n276), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n255), .A2(G238), .A3(new_n260), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT71), .ZN(new_n426));
  AND3_X1   g0226(.A1(new_n259), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n426), .B1(new_n259), .B2(new_n425), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n424), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT13), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT13), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n424), .B(new_n431), .C1(new_n427), .C2(new_n428), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n430), .A2(KEYINPUT72), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT72), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n429), .A2(new_n434), .A3(KEYINPUT13), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n433), .A2(G169), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT73), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT14), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n430), .A2(G179), .A3(new_n432), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n433), .A2(G169), .A3(new_n435), .A4(new_n438), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n294), .A2(new_n214), .ZN(new_n444));
  XNOR2_X1  g0244(.A(new_n444), .B(KEYINPUT12), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n285), .A2(G50), .B1(G20), .B2(new_n214), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(new_n406), .B2(new_n403), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n447), .A2(KEYINPUT11), .A3(new_n291), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n295), .A2(G68), .A3(new_n315), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n445), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(KEYINPUT11), .B1(new_n447), .B2(new_n291), .ZN(new_n451));
  OR2_X1    g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n443), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n433), .A2(G200), .A3(new_n435), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n432), .A2(G190), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n452), .B1(new_n455), .B2(new_n430), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n419), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(G250), .B(G1698), .C1(new_n330), .C2(new_n331), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G283), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(G1698), .ZN(new_n464));
  OAI211_X1 g0264(.A(G244), .B(new_n464), .C1(new_n330), .C2(new_n331), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT4), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n465), .A2(KEYINPUT80), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n466), .B1(new_n465), .B2(KEYINPUT80), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n276), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n257), .A2(G1), .ZN(new_n471));
  XNOR2_X1  g0271(.A(KEYINPUT5), .B(G41), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n255), .A2(G274), .A3(new_n471), .A4(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(KEYINPUT5), .A2(G41), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(KEYINPUT5), .A2(G41), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n471), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n255), .A2(new_n477), .A3(G257), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT81), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n473), .A2(new_n478), .A3(KEYINPUT81), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n470), .A2(new_n281), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT83), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n482), .ZN(new_n486));
  AOI21_X1  g0286(.A(KEYINPUT81), .B1(new_n473), .B2(new_n478), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n488), .A2(KEYINPUT83), .A3(new_n281), .A4(new_n470), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n393), .B1(new_n345), .B2(new_n347), .ZN(new_n491));
  XNOR2_X1  g0291(.A(KEYINPUT78), .B(G107), .ZN(new_n492));
  INV_X1    g0292(.A(G97), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n493), .A2(new_n393), .A3(KEYINPUT6), .ZN(new_n494));
  OR2_X1    g0294(.A1(new_n493), .A2(KEYINPUT6), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n492), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n393), .A2(KEYINPUT78), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT78), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G107), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n495), .A2(new_n494), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(G20), .B1(new_n496), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n285), .A2(G77), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n291), .B1(new_n491), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n293), .A2(G1), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G20), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n206), .A2(G33), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n321), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT79), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n295), .A2(KEYINPUT79), .A3(new_n507), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n510), .A2(new_n511), .A3(G97), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n294), .A2(new_n493), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n479), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n470), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n504), .A2(new_n515), .B1(new_n517), .B2(new_n299), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n490), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n481), .A2(new_n482), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n461), .A2(new_n462), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT80), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n522), .B1(new_n270), .B2(G244), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n521), .B1(new_n523), .B2(new_n466), .ZN(new_n524));
  INV_X1    g0324(.A(new_n469), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n275), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(KEYINPUT82), .B1(new_n520), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT82), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n470), .A2(new_n528), .A3(new_n481), .A4(new_n482), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n527), .A2(G200), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n470), .A2(G190), .A3(new_n516), .ZN(new_n531));
  AND3_X1   g0331(.A1(new_n504), .A2(new_n531), .A3(new_n515), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n510), .A2(new_n511), .A3(G87), .ZN(new_n534));
  AOI21_X1  g0334(.A(G20), .B1(new_n266), .B2(new_n267), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G68), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT19), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(new_n406), .B2(new_n493), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n207), .B1(new_n420), .B2(new_n537), .ZN(new_n539));
  INV_X1    g0339(.A(G87), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n540), .A2(new_n493), .A3(new_n393), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n536), .A2(new_n538), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n291), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n405), .A2(new_n294), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n534), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT85), .ZN(new_n547));
  OAI211_X1 g0347(.A(G238), .B(new_n464), .C1(new_n330), .C2(new_n331), .ZN(new_n548));
  OAI211_X1 g0348(.A(G244), .B(G1698), .C1(new_n330), .C2(new_n331), .ZN(new_n549));
  NAND2_X1  g0349(.A1(KEYINPUT84), .A2(G116), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(KEYINPUT84), .A2(G116), .ZN(new_n552));
  OAI21_X1  g0352(.A(G33), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n548), .A2(new_n549), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n276), .ZN(new_n555));
  INV_X1    g0355(.A(G274), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n206), .A2(new_n556), .A3(G45), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(new_n471), .B2(G250), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n255), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n547), .B1(new_n561), .B2(new_n417), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n554), .A2(new_n276), .B1(new_n255), .B2(new_n559), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n563), .A2(KEYINPUT85), .A3(G190), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n546), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n561), .A2(G200), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n555), .A2(new_n281), .A3(new_n560), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n567), .B1(new_n299), .B2(new_n561), .ZN(new_n568));
  INV_X1    g0368(.A(new_n405), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n510), .A2(new_n511), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n570), .A2(new_n544), .A3(new_n545), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n565), .A2(new_n566), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n519), .A2(new_n533), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n473), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n255), .A2(new_n477), .A3(G270), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT86), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n255), .A2(new_n477), .A3(KEYINPUT86), .A4(G270), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n574), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(G264), .B(G1698), .C1(new_n330), .C2(new_n331), .ZN(new_n580));
  OAI211_X1 g0380(.A(G257), .B(new_n464), .C1(new_n330), .C2(new_n331), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n266), .A2(G303), .A3(new_n267), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT87), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n580), .A2(new_n581), .A3(KEYINPUT87), .A4(new_n582), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n585), .A2(new_n276), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n579), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(G190), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n321), .A2(new_n506), .A3(G116), .A4(new_n507), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT84), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n223), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n593), .A2(G20), .A3(new_n550), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n462), .B(new_n207), .C1(G33), .C2(new_n493), .ZN(new_n595));
  NOR2_X1   g0395(.A1(KEYINPUT88), .A2(KEYINPUT20), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n594), .A2(new_n291), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n591), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n594), .A2(new_n291), .A3(new_n595), .ZN(new_n599));
  XOR2_X1   g0399(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n600));
  NOR2_X1   g0400(.A1(new_n551), .A2(new_n552), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n599), .A2(new_n600), .B1(new_n601), .B2(new_n294), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n603), .B1(new_n588), .B2(G200), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n590), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n589), .A2(G179), .A3(new_n603), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n299), .B1(new_n598), .B2(new_n602), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n588), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(KEYINPUT21), .B1(new_n608), .B2(KEYINPUT89), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT89), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT21), .ZN(new_n611));
  AOI211_X1 g0411(.A(new_n610), .B(new_n611), .C1(new_n588), .C2(new_n607), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n605), .B(new_n606), .C1(new_n609), .C2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT23), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n616), .A2(new_n393), .A3(G20), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n265), .B1(new_n593), .B2(new_n550), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n618), .B1(new_n207), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT22), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n621), .B1(new_n535), .B2(G87), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n207), .B(G87), .C1(new_n330), .C2(new_n331), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n623), .A2(KEYINPUT22), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n620), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(KEYINPUT90), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n623), .A2(KEYINPUT22), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n268), .A2(new_n621), .A3(new_n207), .A4(G87), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT90), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n629), .A2(new_n630), .A3(new_n620), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n626), .A2(KEYINPUT24), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n630), .B1(new_n629), .B2(new_n620), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT24), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n321), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n506), .A2(G107), .ZN(new_n637));
  XNOR2_X1  g0437(.A(new_n637), .B(KEYINPUT25), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n510), .A2(new_n511), .A3(G107), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  OAI211_X1 g0441(.A(G257), .B(G1698), .C1(new_n330), .C2(new_n331), .ZN(new_n642));
  OAI211_X1 g0442(.A(G250), .B(new_n464), .C1(new_n330), .C2(new_n331), .ZN(new_n643));
  NAND2_X1  g0443(.A1(G33), .A2(G294), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n276), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n255), .A2(new_n477), .A3(G264), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n646), .A2(new_n473), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n383), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(G190), .B2(new_n648), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n636), .A2(new_n641), .A3(new_n650), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n646), .A2(G179), .A3(new_n647), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n652), .A2(new_n473), .B1(new_n648), .B2(G169), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n653), .B1(new_n636), .B2(new_n641), .ZN(new_n654));
  OAI21_X1  g0454(.A(KEYINPUT91), .B1(new_n651), .B2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n640), .B1(new_n632), .B2(new_n635), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n650), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT91), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n657), .B(new_n658), .C1(new_n656), .C2(new_n653), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n573), .A2(new_n614), .A3(new_n655), .A4(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n460), .A2(new_n660), .ZN(G372));
  INV_X1    g0461(.A(KEYINPUT93), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT92), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n559), .A2(new_n663), .A3(new_n255), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n251), .A2(new_n253), .A3(new_n254), .ZN(new_n665));
  OAI21_X1  g0465(.A(KEYINPUT92), .B1(new_n665), .B2(new_n558), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(G169), .B1(new_n667), .B2(new_n555), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n662), .B1(new_n668), .B2(new_n567), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n563), .A2(new_n281), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n664), .A2(new_n666), .B1(new_n276), .B2(new_n554), .ZN(new_n671));
  OAI211_X1 g0471(.A(new_n670), .B(KEYINPUT93), .C1(new_n671), .C2(G169), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n571), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n606), .B1(new_n609), .B2(new_n612), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(new_n654), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n671), .A2(new_n383), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n565), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n519), .A2(new_n533), .A3(new_n657), .A4(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n674), .B1(new_n676), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n373), .A2(G107), .ZN(new_n681));
  INV_X1    g0481(.A(new_n492), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n495), .A2(new_n494), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n492), .A2(new_n494), .A3(new_n495), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n686), .A2(G20), .B1(G77), .B2(new_n285), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n321), .B1(new_n681), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n524), .A2(new_n525), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n479), .B1(new_n689), .B2(new_n276), .ZN(new_n690));
  OAI22_X1  g0490(.A1(new_n688), .A2(new_n514), .B1(new_n690), .B2(G169), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(new_n485), .B2(new_n489), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n673), .A2(new_n571), .B1(new_n565), .B2(new_n677), .ZN(new_n693));
  AOI21_X1  g0493(.A(KEYINPUT26), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n562), .A2(new_n564), .ZN(new_n695));
  INV_X1    g0495(.A(new_n546), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(new_n566), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n568), .A2(new_n571), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n490), .A2(new_n518), .A3(new_n697), .A4(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT26), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n694), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n680), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n460), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT94), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n398), .B(KEYINPUT69), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(new_n413), .ZN(new_n707));
  AOI22_X1  g0507(.A1(new_n443), .A2(new_n452), .B1(new_n457), .B2(new_n707), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n365), .B(new_n379), .C1(new_n708), .C2(new_n390), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n311), .A2(new_n313), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n301), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n705), .A2(new_n711), .ZN(G369));
  INV_X1    g0512(.A(new_n675), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n505), .A2(new_n207), .ZN(new_n714));
  OR2_X1    g0514(.A1(new_n714), .A2(KEYINPUT27), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(KEYINPUT27), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n715), .A2(new_n716), .A3(G213), .ZN(new_n717));
  INV_X1    g0517(.A(G343), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n603), .A2(new_n719), .ZN(new_n720));
  MUX2_X1   g0520(.A(new_n713), .B(new_n613), .S(new_n720), .Z(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT95), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n722), .A2(G330), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n655), .A2(new_n659), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n719), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n725), .B1(new_n656), .B2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n654), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n727), .B1(new_n728), .B2(new_n726), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n723), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n713), .A2(new_n719), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n725), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(new_n728), .B2(new_n719), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n731), .A2(new_n734), .ZN(G399));
  INV_X1    g0535(.A(new_n210), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G41), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n541), .A2(G116), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n738), .A2(G1), .A3(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(new_n216), .B2(new_n738), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT28), .ZN(new_n742));
  INV_X1    g0542(.A(new_n674), .ZN(new_n743));
  INV_X1    g0543(.A(new_n679), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n728), .B(new_n606), .C1(new_n609), .C2(new_n612), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n699), .A2(new_n700), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(KEYINPUT97), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n692), .A2(new_n693), .A3(KEYINPUT26), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT97), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n699), .A2(new_n750), .A3(new_n700), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n748), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n719), .B1(new_n746), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(KEYINPUT29), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT29), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(new_n703), .B2(new_n719), .ZN(new_n756));
  AND2_X1   g0556(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(G330), .ZN(new_n758));
  OAI21_X1  g0558(.A(KEYINPUT96), .B1(new_n660), .B2(new_n719), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n490), .A2(new_n518), .B1(new_n530), .B2(new_n532), .ZN(new_n760));
  AND4_X1   g0560(.A1(new_n655), .A2(new_n760), .A3(new_n659), .A4(new_n572), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT96), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n761), .A2(new_n762), .A3(new_n614), .A4(new_n726), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  AND2_X1   g0564(.A1(new_n652), .A2(new_n563), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n765), .A2(new_n589), .A3(new_n690), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT30), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n765), .A2(new_n589), .A3(KEYINPUT30), .A4(new_n690), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n488), .A2(new_n470), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n671), .A2(G179), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n770), .A2(new_n588), .A3(new_n648), .A4(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n768), .A2(new_n769), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(new_n719), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT31), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n774), .B(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n758), .B1(new_n764), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n757), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n742), .B1(new_n779), .B2(G1), .ZN(G364));
  NOR2_X1   g0580(.A1(new_n293), .A2(G20), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n206), .B1(new_n781), .B2(G45), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n737), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n723), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(G330), .B2(new_n722), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n218), .B1(G20), .B2(new_n299), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n207), .A2(G179), .ZN(new_n788));
  NOR2_X1   g0588(.A1(G190), .A2(G200), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G159), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n788), .A2(new_n417), .A3(G200), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n792), .A2(KEYINPUT32), .B1(G107), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n207), .A2(new_n281), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G200), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n417), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR3_X1   g0599(.A1(new_n417), .A2(G179), .A3(G200), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n207), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n795), .B1(new_n202), .B2(new_n799), .C1(new_n493), .C2(new_n801), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n788), .A2(G190), .A3(G200), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(G87), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n797), .A2(G190), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n805), .B1(new_n792), .B2(KEYINPUT32), .C1(new_n807), .C2(new_n214), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n796), .A2(new_n789), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n796), .A2(G190), .A3(new_n383), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n268), .B1(new_n809), .B2(new_n403), .C1(new_n213), .C2(new_n810), .ZN(new_n811));
  NOR3_X1   g0611(.A1(new_n802), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n810), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n813), .A2(G322), .B1(new_n791), .B2(G329), .ZN(new_n814));
  INV_X1    g0614(.A(G311), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n814), .B(new_n269), .C1(new_n815), .C2(new_n809), .ZN(new_n816));
  INV_X1    g0616(.A(G317), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(KEYINPUT33), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n817), .A2(KEYINPUT33), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n806), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n798), .A2(G326), .ZN(new_n821));
  INV_X1    g0621(.A(G303), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n820), .B(new_n821), .C1(new_n822), .C2(new_n803), .ZN(new_n823));
  INV_X1    g0623(.A(G294), .ZN(new_n824));
  INV_X1    g0624(.A(G283), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n801), .A2(new_n824), .B1(new_n793), .B2(new_n825), .ZN(new_n826));
  NOR3_X1   g0626(.A1(new_n816), .A2(new_n823), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n787), .B1(new_n812), .B2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n784), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n210), .A2(G355), .A3(new_n268), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n736), .A2(new_n268), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(G45), .B2(new_n216), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n248), .A2(new_n257), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n830), .B1(G116), .B2(new_n210), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(G13), .A2(G33), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n836), .A2(G20), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n837), .A2(new_n787), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n829), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n837), .B(KEYINPUT98), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n828), .B(new_n839), .C1(new_n722), .C2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n786), .A2(new_n841), .ZN(G396));
  NOR2_X1   g0642(.A1(new_n787), .A2(new_n835), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT99), .Z(new_n844));
  OAI21_X1  g0644(.A(new_n784), .B1(new_n844), .B2(G77), .ZN(new_n845));
  INV_X1    g0645(.A(new_n809), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n813), .A2(G143), .B1(new_n846), .B2(G159), .ZN(new_n847));
  INV_X1    g0647(.A(G150), .ZN(new_n848));
  INV_X1    g0648(.A(G137), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n847), .B1(new_n807), .B2(new_n848), .C1(new_n849), .C2(new_n799), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT34), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n794), .A2(G68), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n269), .B1(new_n791), .B2(G132), .ZN(new_n854));
  INV_X1    g0654(.A(new_n801), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n855), .A2(G58), .B1(new_n804), .B2(G50), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n852), .A2(new_n853), .A3(new_n854), .A4(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n850), .A2(new_n851), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n793), .A2(new_n540), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(G303), .B2(new_n798), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n393), .B2(new_n803), .ZN(new_n861));
  AOI22_X1  g0661(.A1(G97), .A2(new_n855), .B1(new_n806), .B2(G283), .ZN(new_n862));
  INV_X1    g0662(.A(new_n601), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n268), .B1(new_n846), .B2(new_n863), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n813), .A2(G294), .B1(new_n791), .B2(G311), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n862), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n857), .A2(new_n858), .B1(new_n861), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT100), .ZN(new_n868));
  OR2_X1    g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n787), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n867), .B2(new_n868), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n845), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n412), .A2(new_n719), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n415), .A2(new_n418), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n707), .A2(new_n412), .A3(new_n719), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n872), .B1(new_n876), .B2(new_n836), .ZN(new_n877));
  INV_X1    g0677(.A(new_n876), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(new_n703), .B2(new_n719), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n876), .B(new_n726), .C1(new_n680), .C2(new_n702), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n881), .A2(new_n778), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n829), .B1(new_n881), .B2(new_n778), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n877), .B1(new_n882), .B2(new_n883), .ZN(G384));
  NOR2_X1   g0684(.A1(new_n781), .A2(new_n206), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n519), .A2(new_n533), .A3(new_n572), .ZN(new_n886));
  NOR3_X1   g0686(.A1(new_n724), .A2(new_n613), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n762), .B1(new_n887), .B2(new_n726), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n655), .A2(new_n760), .A3(new_n659), .A4(new_n572), .ZN(new_n889));
  NOR4_X1   g0689(.A1(new_n889), .A2(KEYINPUT96), .A3(new_n613), .A4(new_n719), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n777), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n343), .B1(new_n341), .B2(KEYINPUT101), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT101), .ZN(new_n893));
  AOI211_X1 g0693(.A(new_n893), .B(new_n329), .C1(new_n340), .C2(G68), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n342), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n717), .B1(new_n895), .B2(new_n319), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n380), .B2(new_n390), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT37), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n895), .A2(new_n319), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n899), .A2(new_n378), .B1(new_n350), .B2(new_n385), .ZN(new_n900));
  INV_X1    g0700(.A(new_n896), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n376), .A2(new_n378), .ZN(new_n903));
  XOR2_X1   g0703(.A(new_n717), .B(KEYINPUT102), .Z(new_n904));
  NAND2_X1  g0704(.A1(new_n376), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n903), .A2(new_n905), .A3(new_n898), .A4(new_n386), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n897), .B1(new_n902), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT38), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n897), .B(KEYINPUT38), .C1(new_n902), .C2(new_n907), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n452), .A2(new_n719), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n453), .A2(new_n457), .A3(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n457), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n452), .B(new_n719), .C1(new_n443), .C2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n891), .A2(new_n912), .A3(new_n876), .A4(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT40), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n386), .B1(new_n350), .B2(new_n364), .ZN(new_n921));
  INV_X1    g0721(.A(new_n904), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n350), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(KEYINPUT37), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n906), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n923), .B1(new_n380), .B2(new_n390), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n909), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n919), .B1(new_n928), .B2(new_n911), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n891), .A2(new_n929), .A3(new_n876), .A4(new_n917), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n920), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n776), .B1(new_n759), .B2(new_n763), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n460), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n758), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n931), .B2(new_n933), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n757), .A2(new_n459), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n711), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n707), .A2(new_n726), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n880), .A2(new_n938), .B1(new_n914), .B2(new_n916), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n939), .A2(new_n912), .B1(new_n380), .B2(new_n922), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT39), .ZN(new_n941));
  INV_X1    g0741(.A(new_n911), .ZN(new_n942));
  AOI21_X1  g0742(.A(KEYINPUT38), .B1(new_n925), .B2(new_n926), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n453), .A2(new_n719), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n910), .A2(KEYINPUT39), .A3(new_n911), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n940), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n937), .B(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n885), .B1(new_n935), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n949), .B2(new_n935), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n219), .A2(G116), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(new_n686), .B2(KEYINPUT35), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(KEYINPUT35), .B2(new_n686), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT36), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n322), .A2(G77), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n244), .B1(new_n216), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n957), .A2(G1), .A3(new_n293), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n951), .A2(new_n955), .A3(new_n958), .ZN(G367));
  NAND2_X1  g0759(.A1(new_n546), .A2(new_n719), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n674), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(new_n693), .B2(new_n960), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT43), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n719), .B1(new_n688), .B2(new_n514), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n760), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n519), .B2(new_n726), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT103), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n967), .A2(new_n968), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n972), .A2(new_n733), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT42), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n971), .A2(new_n654), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n719), .B1(new_n975), .B2(new_n519), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n964), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n962), .A2(new_n963), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n978), .B(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n730), .A2(new_n972), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n980), .B(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n737), .B(new_n983), .Z(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n972), .A2(new_n734), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT44), .Z(new_n987));
  NOR2_X1   g0787(.A1(new_n972), .A2(new_n734), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT45), .ZN(new_n989));
  AND3_X1   g0789(.A1(new_n987), .A2(new_n730), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n730), .B1(new_n987), .B2(new_n989), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n733), .B1(new_n729), .B2(new_n732), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n723), .B(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n992), .A2(new_n779), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n985), .B1(new_n995), .B2(new_n779), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n982), .B1(new_n996), .B2(new_n783), .ZN(new_n997));
  INV_X1    g0797(.A(new_n831), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n838), .B1(new_n210), .B2(new_n405), .C1(new_n998), .C2(new_n239), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n810), .A2(new_n822), .B1(new_n809), .B2(new_n825), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n268), .B(new_n1000), .C1(G317), .C2(new_n791), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n806), .A2(G294), .B1(new_n794), .B2(G97), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n803), .A2(new_n601), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1001), .B(new_n1002), .C1(KEYINPUT46), .C2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n804), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n393), .B2(new_n801), .C1(new_n799), .C2(new_n815), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n801), .A2(new_n214), .B1(new_n810), .B2(new_n848), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT105), .Z(new_n1008));
  OAI22_X1  g0808(.A1(new_n809), .A2(new_n202), .B1(new_n790), .B2(new_n849), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(G143), .B2(new_n798), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n268), .B1(new_n793), .B2(new_n403), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT106), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n806), .A2(G159), .B1(new_n804), .B2(G58), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1010), .A2(new_n1013), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n1004), .A2(new_n1006), .B1(new_n1008), .B2(new_n1016), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT47), .Z(new_n1018));
  OAI211_X1 g0818(.A(new_n784), .B(new_n999), .C1(new_n1018), .C2(new_n870), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n840), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1019), .B1(new_n1020), .B2(new_n962), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n997), .A2(new_n1022), .ZN(G387));
  OR2_X1    g0823(.A1(new_n729), .A2(new_n840), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n739), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1025), .A2(new_n210), .A3(new_n268), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(G107), .B2(new_n210), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n236), .A2(new_n257), .ZN(new_n1028));
  AOI211_X1 g0828(.A(G45), .B(new_n1025), .C1(G68), .C2(G77), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n318), .A2(G50), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT50), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n998), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1027), .B1(new_n1028), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n838), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n784), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n809), .A2(new_n214), .B1(new_n790), .B2(new_n848), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n269), .B(new_n1036), .C1(G50), .C2(new_n813), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n804), .A2(G77), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n569), .A2(new_n855), .B1(new_n806), .B2(new_n283), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n798), .A2(G159), .B1(new_n794), .B2(G97), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n268), .B1(new_n791), .B2(G326), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n801), .A2(new_n825), .B1(new_n803), .B2(new_n824), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n813), .A2(G317), .B1(new_n846), .B2(G303), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n798), .A2(G322), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1044), .B(new_n1045), .C1(new_n815), .C2(new_n807), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT48), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1043), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n1047), .B2(new_n1046), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT49), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1042), .B1(new_n601), .B2(new_n793), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  AND2_X1   g0851(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1041), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1035), .B1(new_n1053), .B2(new_n787), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n994), .A2(new_n783), .B1(new_n1024), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n994), .A2(new_n779), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n737), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n994), .A2(new_n779), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1055), .B1(new_n1057), .B2(new_n1058), .ZN(G393));
  OAI21_X1  g0859(.A(new_n1056), .B1(new_n990), .B2(new_n991), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n995), .A2(new_n737), .A3(new_n1060), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n807), .A2(new_n202), .B1(new_n809), .B2(new_n318), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1062), .A2(KEYINPUT107), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(KEYINPUT107), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n269), .B(new_n859), .C1(G143), .C2(new_n791), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n801), .A2(new_n403), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(G68), .B2(new_n804), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .A4(new_n1067), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(G150), .A2(new_n798), .B1(new_n813), .B2(G159), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT51), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n855), .A2(new_n863), .B1(new_n804), .B2(G283), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n806), .A2(G303), .B1(new_n794), .B2(G107), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n846), .A2(G294), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n268), .B1(new_n791), .B2(G322), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(G317), .A2(new_n798), .B1(new_n813), .B2(G311), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT52), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n1068), .A2(new_n1070), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n787), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n831), .A2(new_n243), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1080), .B(new_n838), .C1(new_n493), .C2(new_n210), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1079), .A2(new_n784), .A3(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n972), .B2(new_n837), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n992), .B2(new_n783), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1061), .A2(new_n1084), .ZN(G390));
  NAND4_X1  g0885(.A1(new_n778), .A2(KEYINPUT108), .A3(new_n876), .A4(new_n917), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n880), .A2(new_n938), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n917), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n945), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n1088), .A2(new_n1089), .B1(new_n944), .B2(new_n946), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1089), .B1(new_n942), .B2(new_n943), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n749), .A2(new_n751), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n750), .B1(new_n699), .B2(new_n700), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n726), .B(new_n876), .C1(new_n1094), .C2(new_n680), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n938), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1091), .B1(new_n917), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1086), .B1(new_n1090), .B2(new_n1097), .ZN(new_n1098));
  AND3_X1   g0898(.A1(new_n910), .A2(KEYINPUT39), .A3(new_n911), .ZN(new_n1099));
  AOI21_X1  g0899(.A(KEYINPUT39), .B1(new_n928), .B2(new_n911), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n1099), .A2(new_n1100), .B1(new_n939), .B2(new_n945), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n914), .A2(new_n916), .ZN(new_n1102));
  NOR4_X1   g0902(.A1(new_n932), .A2(new_n1102), .A3(new_n758), .A4(new_n878), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n945), .B1(new_n928), .B2(new_n911), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n938), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n753), .B2(new_n876), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1104), .B1(new_n1106), .B2(new_n1102), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1101), .A2(new_n1103), .A3(KEYINPUT108), .A4(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1098), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n778), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n936), .B(new_n711), .C1(new_n460), .C2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n917), .B1(new_n778), .B2(new_n876), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1087), .B1(new_n1112), .B2(new_n1103), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n891), .A2(G330), .A3(new_n876), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n1102), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n778), .A2(new_n876), .A3(new_n917), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1115), .A2(new_n1116), .A3(new_n1106), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1111), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT109), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1109), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n460), .A2(new_n1110), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n937), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1124), .A2(KEYINPUT109), .A3(new_n1098), .A4(new_n1108), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1120), .A2(new_n1125), .A3(new_n737), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n784), .B1(new_n844), .B2(new_n283), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n836), .B1(new_n944), .B2(new_n946), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n791), .A2(G125), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n269), .B(new_n1129), .C1(G132), .C2(new_n813), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(G159), .A2(new_n855), .B1(new_n798), .B2(G128), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n806), .A2(G137), .B1(new_n794), .B2(G50), .ZN(new_n1132));
  XOR2_X1   g0932(.A(KEYINPUT54), .B(G143), .Z(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT111), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n846), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .A4(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n804), .A2(G150), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT53), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n810), .A2(new_n223), .B1(new_n790), .B2(new_n824), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n268), .B(new_n1139), .C1(G97), .C2(new_n846), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1140), .A2(new_n805), .A3(new_n853), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1066), .B1(G283), .B2(new_n798), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n393), .B2(new_n807), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n1136), .A2(new_n1138), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1127), .B(new_n1128), .C1(new_n787), .C2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1109), .A2(new_n783), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(KEYINPUT110), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT110), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1109), .A2(new_n1148), .A3(new_n783), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1145), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1126), .A2(new_n1150), .ZN(G378));
  INV_X1    g0951(.A(new_n301), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n710), .A2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n303), .A2(new_n717), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1154), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n314), .A2(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1155), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1158), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n314), .A2(new_n1156), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n301), .B(new_n1154), .C1(new_n311), .C2(new_n313), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1160), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  AND2_X1   g0963(.A1(new_n1159), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n835), .ZN(new_n1165));
  AOI211_X1 g0965(.A(G41), .B(new_n268), .C1(new_n791), .C2(G283), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1166), .B(new_n1038), .C1(new_n213), .C2(new_n793), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT112), .Z(new_n1168));
  OAI22_X1  g0968(.A1(new_n810), .A2(new_n393), .B1(new_n809), .B2(new_n405), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(G68), .B2(new_n855), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G97), .A2(new_n806), .B1(new_n798), .B2(G116), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1168), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT58), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(G33), .A2(G41), .ZN(new_n1174));
  AOI211_X1 g0974(.A(G50), .B(new_n1174), .C1(new_n269), .C2(new_n256), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1134), .A2(new_n804), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n806), .A2(G132), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n813), .A2(G128), .B1(new_n846), .B2(G137), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(G150), .A2(new_n855), .B1(new_n798), .B2(G125), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1180), .A2(KEYINPUT59), .ZN(new_n1181));
  INV_X1    g0981(.A(G124), .ZN(new_n1182));
  INV_X1    g0982(.A(G159), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1174), .B1(new_n790), .B2(new_n1182), .C1(new_n1183), .C2(new_n793), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n1180), .B2(KEYINPUT59), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1175), .B1(new_n1181), .B2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1173), .A2(KEYINPUT113), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(KEYINPUT113), .B1(new_n1173), .B2(new_n1186), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1188), .A2(new_n870), .A3(new_n1189), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n829), .B(new_n1190), .C1(new_n202), .C2(new_n843), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1165), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1159), .A2(new_n1163), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n932), .A2(new_n1102), .A3(new_n878), .ZN(new_n1194));
  AOI21_X1  g0994(.A(KEYINPUT40), .B1(new_n1194), .B2(new_n912), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n930), .A2(G330), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1193), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n758), .B1(new_n1194), .B2(new_n929), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1198), .A2(new_n1164), .A3(new_n920), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n948), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT115), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n948), .ZN(new_n1203));
  OR2_X1    g1003(.A1(new_n1203), .A2(KEYINPUT114), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n1200), .A2(KEYINPUT115), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1192), .B1(new_n1207), .B2(new_n782), .ZN(new_n1208));
  NOR3_X1   g1008(.A1(new_n1195), .A2(new_n1196), .A3(new_n1193), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1164), .B1(new_n1198), .B2(new_n920), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1203), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT116), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1197), .A2(new_n948), .A3(new_n1199), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT57), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1109), .A2(new_n1121), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1215), .B1(new_n1216), .B2(new_n1123), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1197), .A2(new_n1199), .A3(KEYINPUT116), .A4(new_n948), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1214), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n737), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1216), .A2(new_n1123), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1220), .A2(KEYINPUT117), .B1(new_n1222), .B2(new_n1215), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT117), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1219), .A2(new_n1224), .A3(new_n737), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1208), .B1(new_n1223), .B2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(G375));
  NAND3_X1  g1027(.A1(new_n1111), .A2(new_n1113), .A3(new_n1117), .ZN(new_n1228));
  XOR2_X1   g1028(.A(new_n984), .B(KEYINPUT118), .Z(new_n1229));
  NAND3_X1  g1029(.A1(new_n1124), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1102), .A2(new_n835), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n784), .B1(new_n844), .B2(G68), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n801), .A2(new_n405), .B1(new_n810), .B2(new_n825), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT120), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n809), .A2(new_n393), .B1(new_n790), .B2(new_n822), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G294), .B2(new_n798), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n806), .A2(new_n863), .B1(new_n804), .B2(G97), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1234), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n268), .B1(new_n794), .B2(G77), .ZN(new_n1239));
  XOR2_X1   g1039(.A(new_n1239), .B(KEYINPUT119), .Z(new_n1240));
  NAND2_X1  g1040(.A1(new_n798), .A2(G132), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1241), .B(KEYINPUT121), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n801), .A2(new_n202), .B1(new_n793), .B2(new_n213), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(G159), .B2(new_n804), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1134), .A2(new_n806), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n269), .B1(new_n791), .B2(G128), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n813), .A2(G137), .B1(new_n846), .B2(G150), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .A4(new_n1247), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n1238), .A2(new_n1240), .B1(new_n1242), .B2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1232), .B1(new_n1249), .B2(new_n787), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n1121), .A2(new_n783), .B1(new_n1231), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1230), .A2(new_n1251), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n1252), .B(KEYINPUT122), .ZN(G381));
  OR4_X1    g1053(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1254));
  NOR3_X1   g1054(.A1(new_n1254), .A2(G387), .A3(G381), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1126), .A2(KEYINPUT123), .A3(new_n1150), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(KEYINPUT123), .B1(new_n1126), .B2(new_n1150), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1255), .A2(new_n1226), .A3(new_n1259), .ZN(G407));
  NAND2_X1  g1060(.A1(new_n718), .A2(G213), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1226), .A2(new_n1259), .A3(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(G407), .A2(G213), .A3(new_n1263), .ZN(G409));
  INV_X1    g1064(.A(G390), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(G387), .A2(new_n1265), .ZN(new_n1266));
  XOR2_X1   g1066(.A(G393), .B(G396), .Z(new_n1267));
  NAND3_X1  g1067(.A1(new_n997), .A2(new_n1022), .A3(G390), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1266), .A2(new_n1267), .A3(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1267), .B1(new_n1266), .B2(new_n1268), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1124), .A2(KEYINPUT60), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1228), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1111), .A2(KEYINPUT60), .A3(new_n1113), .A4(new_n1117), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1274), .A2(new_n737), .A3(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT125), .ZN(new_n1277));
  OR2_X1    g1077(.A1(G384), .A2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1251), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1276), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(G384), .A2(new_n1277), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(new_n1281), .B(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(G378), .ZN(new_n1285));
  AOI211_X1 g1085(.A(new_n1285), .B(new_n1208), .C1(new_n1223), .C2(new_n1225), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT123), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(G378), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n1256), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1214), .A2(new_n783), .A3(new_n1218), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT124), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1290), .A2(new_n1291), .A3(new_n1192), .ZN(new_n1292));
  OAI211_X1 g1092(.A(new_n1221), .B(new_n1229), .C1(new_n1205), .C2(new_n1206), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1291), .B1(new_n1290), .B2(new_n1192), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1289), .B1(new_n1292), .B2(new_n1296), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1261), .B(new_n1284), .C1(new_n1286), .C2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(KEYINPUT126), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1220), .A2(KEYINPUT117), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1222), .A2(new_n1215), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1300), .A2(new_n1225), .A3(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1208), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1302), .A2(G378), .A3(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1290), .A2(new_n1192), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(KEYINPUT124), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1306), .A2(new_n1292), .A3(new_n1293), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(new_n1259), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1262), .B1(new_n1304), .B2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT126), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1309), .A2(new_n1310), .A3(new_n1284), .ZN(new_n1311));
  AOI21_X1  g1111(.A(KEYINPUT62), .B1(new_n1299), .B2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1281), .A2(new_n1277), .A3(G384), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1276), .A2(new_n1280), .A3(new_n1282), .ZN(new_n1314));
  AND2_X1   g1114(.A1(new_n1262), .A2(G2897), .ZN(new_n1315));
  AND3_X1   g1115(.A1(new_n1313), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1315), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  AOI22_X1  g1118(.A1(new_n1226), .A2(G378), .B1(new_n1259), .B2(new_n1307), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1318), .B1(new_n1319), .B2(new_n1262), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT61), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT62), .ZN(new_n1322));
  AOI211_X1 g1122(.A(new_n1262), .B(new_n1283), .C1(new_n1304), .C2(new_n1308), .ZN(new_n1323));
  OAI211_X1 g1123(.A(new_n1320), .B(new_n1321), .C1(new_n1322), .C2(new_n1323), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1272), .B1(new_n1312), .B2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT63), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1299), .A2(new_n1326), .A3(new_n1311), .ZN(new_n1327));
  AND2_X1   g1127(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1323), .A2(KEYINPUT63), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1327), .A2(new_n1328), .A3(new_n1271), .A4(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1325), .A2(new_n1330), .ZN(G405));
  INV_X1    g1131(.A(KEYINPUT127), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1226), .A2(new_n1289), .ZN(new_n1333));
  OR4_X1    g1133(.A1(new_n1332), .A2(new_n1333), .A3(new_n1286), .A4(new_n1283), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1332), .B1(new_n1333), .B2(new_n1286), .ZN(new_n1335));
  OAI211_X1 g1135(.A(new_n1304), .B(KEYINPUT127), .C1(new_n1226), .C2(new_n1289), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1335), .A2(new_n1283), .A3(new_n1336), .ZN(new_n1337));
  AND3_X1   g1137(.A1(new_n1334), .A2(new_n1271), .A3(new_n1337), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1271), .B1(new_n1334), .B2(new_n1337), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1338), .A2(new_n1339), .ZN(G402));
endmodule


