

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765;

  AND2_X1 U377 ( .A1(n440), .A2(n439), .ZN(n637) );
  OR2_X1 U378 ( .A1(n762), .A2(KEYINPUT44), .ZN(n421) );
  NAND2_X1 U379 ( .A1(n609), .A2(n434), .ZN(n610) );
  NAND2_X1 U380 ( .A1(n355), .A2(n386), .ZN(n608) );
  AND2_X1 U381 ( .A1(n601), .A2(n425), .ZN(n609) );
  INV_X1 U382 ( .A(n596), .ZN(n648) );
  XNOR2_X1 U383 ( .A(n541), .B(n540), .ZN(n596) );
  NOR2_X1 U384 ( .A1(n682), .A2(G902), .ZN(n541) );
  XNOR2_X1 U385 ( .A(n537), .B(n539), .ZN(n357) );
  NAND2_X1 U386 ( .A1(n384), .A2(n385), .ZN(n355) );
  XNOR2_X2 U387 ( .A(n518), .B(n474), .ZN(n484) );
  XNOR2_X2 U388 ( .A(n356), .B(G143), .ZN(n518) );
  INV_X4 U389 ( .A(G128), .ZN(n356) );
  NAND2_X1 U390 ( .A1(n703), .A2(n613), .ZN(n614) );
  NAND2_X1 U391 ( .A1(n422), .A2(n612), .ZN(n703) );
  XNOR2_X1 U392 ( .A(n357), .B(n538), .ZN(n682) );
  INV_X1 U393 ( .A(n434), .ZN(n629) );
  INV_X1 U394 ( .A(G953), .ZN(n377) );
  NOR2_X1 U395 ( .A1(n665), .A2(n662), .ZN(n593) );
  XNOR2_X1 U396 ( .A(KEYINPUT38), .B(n629), .ZN(n660) );
  NOR2_X1 U397 ( .A1(n714), .A2(n359), .ZN(n461) );
  AND2_X1 U398 ( .A1(n579), .A2(n364), .ZN(n425) );
  XNOR2_X1 U399 ( .A(n402), .B(KEYINPUT67), .ZN(n620) );
  XNOR2_X1 U400 ( .A(n382), .B(n557), .ZN(n645) );
  XNOR2_X1 U401 ( .A(n467), .B(n465), .ZN(n571) );
  XNOR2_X1 U402 ( .A(n539), .B(n493), .ZN(n744) );
  XOR2_X1 U403 ( .A(G116), .B(G107), .Z(n521) );
  XNOR2_X1 U404 ( .A(G146), .B(G125), .ZN(n506) );
  NOR2_X2 U405 ( .A1(n705), .A2(n447), .ZN(n446) );
  INV_X1 U406 ( .A(n761), .ZN(n439) );
  NOR2_X1 U407 ( .A1(n645), .A2(n450), .ZN(n402) );
  XNOR2_X1 U408 ( .A(n517), .B(n466), .ZN(n465) );
  OR2_X1 U409 ( .A1(n726), .A2(G902), .ZN(n467) );
  INV_X1 U410 ( .A(G475), .ZN(n466) );
  XNOR2_X1 U411 ( .A(n566), .B(n565), .ZN(n643) );
  AND2_X1 U412 ( .A1(n369), .A2(n619), .ZN(n566) );
  XNOR2_X1 U413 ( .A(KEYINPUT69), .B(KEYINPUT34), .ZN(n567) );
  XNOR2_X1 U414 ( .A(n526), .B(n525), .ZN(n572) );
  OR2_X1 U415 ( .A1(n687), .A2(G472), .ZN(n430) );
  XOR2_X1 U416 ( .A(G140), .B(G113), .Z(n513) );
  XNOR2_X1 U417 ( .A(n488), .B(n487), .ZN(n489) );
  INV_X1 U418 ( .A(KEYINPUT17), .ZN(n487) );
  XOR2_X1 U419 ( .A(KEYINPUT25), .B(KEYINPUT72), .Z(n555) );
  XNOR2_X1 U420 ( .A(KEYINPUT81), .B(KEYINPUT45), .ZN(n586) );
  XNOR2_X1 U421 ( .A(n489), .B(n486), .ZN(n394) );
  XNOR2_X1 U422 ( .A(n484), .B(n505), .ZN(n485) );
  INV_X1 U423 ( .A(n506), .ZN(n505) );
  XNOR2_X1 U424 ( .A(n489), .B(n397), .ZN(n396) );
  INV_X1 U425 ( .A(n486), .ZN(n397) );
  XNOR2_X1 U426 ( .A(n406), .B(n499), .ZN(n501) );
  NAND2_X1 U427 ( .A1(G234), .A2(G237), .ZN(n499) );
  XNOR2_X1 U428 ( .A(KEYINPUT14), .B(KEYINPUT88), .ZN(n406) );
  NAND2_X1 U429 ( .A1(n374), .A2(n373), .ZN(n372) );
  INV_X1 U430 ( .A(KEYINPUT28), .ZN(n389) );
  XOR2_X1 U431 ( .A(G101), .B(KEYINPUT3), .Z(n490) );
  XNOR2_X1 U432 ( .A(n405), .B(n361), .ZN(n726) );
  XNOR2_X1 U433 ( .A(n368), .B(n477), .ZN(n367) );
  XNOR2_X1 U434 ( .A(n459), .B(G101), .ZN(n368) );
  NAND2_X1 U435 ( .A1(n360), .A2(n707), .ZN(n627) );
  INV_X1 U436 ( .A(n659), .ZN(n464) );
  NOR2_X1 U437 ( .A1(n456), .A2(n455), .ZN(n400) );
  XNOR2_X1 U438 ( .A(n436), .B(n470), .ZN(n561) );
  INV_X1 U439 ( .A(KEYINPUT22), .ZN(n470) );
  BUF_X1 U440 ( .A(n435), .Z(n434) );
  BUF_X1 U441 ( .A(n648), .Z(n416) );
  NAND2_X1 U442 ( .A1(n428), .A2(n427), .ZN(n426) );
  INV_X1 U443 ( .A(n687), .ZN(n427) );
  XNOR2_X1 U444 ( .A(n552), .B(n749), .ZN(n735) );
  XNOR2_X1 U445 ( .A(n522), .B(n420), .ZN(n524) );
  XNOR2_X1 U446 ( .A(n521), .B(n365), .ZN(n420) );
  XNOR2_X1 U447 ( .A(n726), .B(KEYINPUT59), .ZN(n729) );
  BUF_X2 U448 ( .A(n727), .Z(n733) );
  XOR2_X1 U449 ( .A(KEYINPUT86), .B(n688), .Z(n730) );
  XNOR2_X1 U450 ( .A(n380), .B(n379), .ZN(n378) );
  INV_X1 U451 ( .A(KEYINPUT79), .ZN(n379) );
  NAND2_X1 U452 ( .A1(n642), .A2(n641), .ZN(n380) );
  INV_X1 U453 ( .A(KEYINPUT74), .ZN(n424) );
  INV_X1 U454 ( .A(KEYINPUT47), .ZN(n447) );
  XNOR2_X1 U455 ( .A(n604), .B(KEYINPUT46), .ZN(n442) );
  INV_X1 U456 ( .A(KEYINPUT77), .ZN(n373) );
  INV_X1 U457 ( .A(KEYINPUT105), .ZN(n419) );
  OR2_X1 U458 ( .A1(G237), .A2(G902), .ZN(n497) );
  XNOR2_X1 U459 ( .A(G137), .B(G119), .ZN(n535) );
  XNOR2_X1 U460 ( .A(n484), .B(n476), .ZN(n748) );
  XNOR2_X1 U461 ( .A(n449), .B(n448), .ZN(n542) );
  INV_X1 U462 ( .A(KEYINPUT8), .ZN(n448) );
  NAND2_X1 U463 ( .A1(n377), .A2(G234), .ZN(n449) );
  XNOR2_X1 U464 ( .A(G143), .B(G131), .ZN(n512) );
  XOR2_X1 U465 ( .A(G107), .B(KEYINPUT68), .Z(n481) );
  INV_X1 U466 ( .A(G104), .ZN(n478) );
  XNOR2_X1 U467 ( .A(n381), .B(G140), .ZN(n551) );
  INV_X1 U468 ( .A(G137), .ZN(n381) );
  XNOR2_X1 U469 ( .A(n748), .B(G146), .ZN(n538) );
  XNOR2_X1 U470 ( .A(G902), .B(KEYINPUT15), .ZN(n683) );
  INV_X1 U471 ( .A(n612), .ZN(n455) );
  INV_X1 U472 ( .A(n644), .ZN(n438) );
  AND2_X1 U473 ( .A1(G953), .A2(G902), .ZN(n500) );
  XNOR2_X1 U474 ( .A(n564), .B(n452), .ZN(n369) );
  NAND2_X1 U475 ( .A1(G214), .A2(n497), .ZN(n659) );
  NOR2_X1 U476 ( .A1(n735), .A2(G902), .ZN(n382) );
  XOR2_X1 U477 ( .A(G104), .B(G122), .Z(n507) );
  INV_X1 U478 ( .A(KEYINPUT23), .ZN(n546) );
  XNOR2_X1 U479 ( .A(n409), .B(n744), .ZN(n719) );
  NAND2_X1 U480 ( .A1(n398), .A2(n396), .ZN(n395) );
  NAND2_X1 U481 ( .A1(n485), .A2(n394), .ZN(n393) );
  NOR2_X1 U482 ( .A1(n634), .A2(n633), .ZN(n642) );
  INV_X1 U483 ( .A(KEYINPUT6), .ZN(n418) );
  XNOR2_X1 U484 ( .A(n482), .B(G469), .ZN(n606) );
  NOR2_X1 U485 ( .A1(n721), .A2(G902), .ZN(n482) );
  AND2_X1 U486 ( .A1(n388), .A2(n387), .ZN(n386) );
  XOR2_X1 U487 ( .A(n571), .B(KEYINPUT100), .Z(n573) );
  XNOR2_X1 U488 ( .A(n391), .B(n414), .ZN(n578) );
  INV_X1 U489 ( .A(KEYINPUT89), .ZN(n414) );
  INV_X1 U490 ( .A(n416), .ZN(n451) );
  AND2_X1 U491 ( .A1(n462), .A2(n626), .ZN(n714) );
  XNOR2_X1 U492 ( .A(n458), .B(n568), .ZN(n762) );
  XNOR2_X1 U493 ( .A(n560), .B(KEYINPUT32), .ZN(n763) );
  NAND2_X1 U494 ( .A1(n561), .A2(n469), .ZN(n560) );
  AND2_X1 U495 ( .A1(n559), .A2(n626), .ZN(n469) );
  AND2_X1 U496 ( .A1(n582), .A2(n558), .ZN(n559) );
  NAND2_X1 U497 ( .A1(n363), .A2(n358), .ZN(n699) );
  AND2_X1 U498 ( .A1(n431), .A2(n366), .ZN(n429) );
  XNOR2_X1 U499 ( .A(n734), .B(n735), .ZN(n403) );
  XNOR2_X1 U500 ( .A(n731), .B(n732), .ZN(n412) );
  INV_X1 U501 ( .A(KEYINPUT60), .ZN(n407) );
  XNOR2_X1 U502 ( .A(n724), .B(n725), .ZN(n404) );
  AND2_X1 U503 ( .A1(n679), .A2(n377), .ZN(n376) );
  AND2_X1 U504 ( .A1(n416), .A2(n558), .ZN(n358) );
  XOR2_X1 U505 ( .A(n618), .B(KEYINPUT70), .Z(n359) );
  AND2_X1 U506 ( .A1(n619), .A2(n463), .ZN(n360) );
  XNOR2_X1 U507 ( .A(n606), .B(n483), .ZN(n649) );
  INV_X1 U508 ( .A(n649), .ZN(n626) );
  XOR2_X1 U509 ( .A(n511), .B(n510), .Z(n361) );
  XNOR2_X1 U510 ( .A(n494), .B(n496), .ZN(n362) );
  AND2_X1 U511 ( .A1(n561), .A2(n649), .ZN(n363) );
  XNOR2_X1 U512 ( .A(n648), .B(n418), .ZN(n582) );
  OR2_X1 U513 ( .A1(n592), .A2(n591), .ZN(n364) );
  XOR2_X1 U514 ( .A(G134), .B(G122), .Z(n365) );
  BUF_X1 U515 ( .A(n645), .Z(n411) );
  XOR2_X1 U516 ( .A(KEYINPUT18), .B(KEYINPUT68), .Z(n486) );
  AND2_X1 U517 ( .A1(n430), .A2(n730), .ZN(n366) );
  XNOR2_X1 U518 ( .A(n538), .B(n367), .ZN(n721) );
  XNOR2_X1 U519 ( .A(n480), .B(n481), .ZN(n459) );
  NAND2_X1 U520 ( .A1(n395), .A2(n393), .ZN(n409) );
  NAND2_X1 U521 ( .A1(n423), .A2(n615), .ZN(n616) );
  XNOR2_X1 U522 ( .A(n610), .B(n611), .ZN(n422) );
  AND2_X1 U523 ( .A1(n369), .A2(n451), .ZN(n575) );
  NAND2_X1 U524 ( .A1(n370), .A2(n632), .ZN(n634) );
  NAND2_X1 U525 ( .A1(n371), .A2(n631), .ZN(n370) );
  NAND2_X1 U526 ( .A1(n375), .A2(n372), .ZN(n371) );
  INV_X1 U527 ( .A(n737), .ZN(n374) );
  NAND2_X1 U528 ( .A1(n752), .A2(KEYINPUT78), .ZN(n375) );
  NAND2_X1 U529 ( .A1(n378), .A2(n376), .ZN(n681) );
  NOR2_X1 U530 ( .A1(n648), .A2(n389), .ZN(n384) );
  INV_X1 U531 ( .A(n620), .ZN(n385) );
  NAND2_X1 U532 ( .A1(n648), .A2(n389), .ZN(n387) );
  NAND2_X1 U533 ( .A1(n620), .A2(n389), .ZN(n388) );
  XNOR2_X2 U534 ( .A(n390), .B(KEYINPUT73), .ZN(n705) );
  NAND2_X1 U535 ( .A1(n608), .A2(n607), .ZN(n390) );
  NAND2_X1 U536 ( .A1(n391), .A2(n437), .ZN(n436) );
  NAND2_X1 U537 ( .A1(n654), .A2(n391), .ZN(n576) );
  XNOR2_X2 U538 ( .A(n504), .B(KEYINPUT0), .ZN(n391) );
  NOR2_X2 U539 ( .A1(n392), .A2(KEYINPUT80), .ZN(n684) );
  NOR2_X1 U540 ( .A1(n392), .A2(KEYINPUT77), .ZN(n639) );
  XNOR2_X1 U541 ( .A(n392), .B(n631), .ZN(n685) );
  AND2_X2 U542 ( .A1(n638), .A2(n637), .ZN(n392) );
  INV_X1 U543 ( .A(n485), .ZN(n398) );
  NAND2_X1 U544 ( .A1(n585), .A2(n399), .ZN(n587) );
  NAND2_X1 U545 ( .A1(n421), .A2(n570), .ZN(n399) );
  AND2_X1 U546 ( .A1(n401), .A2(n400), .ZN(n454) );
  NAND2_X1 U547 ( .A1(n457), .A2(n643), .ZN(n401) );
  XOR2_X2 U548 ( .A(G119), .B(G110), .Z(n545) );
  NAND2_X1 U549 ( .A1(n426), .A2(n429), .ZN(n433) );
  NOR2_X1 U550 ( .A1(n403), .A2(n736), .ZN(G66) );
  NAND2_X1 U551 ( .A1(n472), .A2(n730), .ZN(n471) );
  NOR2_X1 U552 ( .A1(n404), .A2(n736), .ZN(G54) );
  XNOR2_X1 U553 ( .A(n717), .B(n473), .ZN(n472) );
  XNOR2_X1 U554 ( .A(n441), .B(n623), .ZN(n440) );
  XNOR2_X1 U555 ( .A(n516), .B(n550), .ZN(n405) );
  NAND2_X1 U556 ( .A1(n364), .A2(n644), .ZN(n450) );
  XNOR2_X1 U557 ( .A(n408), .B(n407), .ZN(G60) );
  NAND2_X1 U558 ( .A1(n415), .A2(n730), .ZN(n408) );
  XNOR2_X1 U559 ( .A(n410), .B(n444), .ZN(n443) );
  NAND2_X1 U560 ( .A1(n460), .A2(n461), .ZN(n410) );
  NOR2_X2 U561 ( .A1(n707), .A2(n710), .ZN(n664) );
  XNOR2_X2 U562 ( .A(n574), .B(KEYINPUT103), .ZN(n707) );
  NOR2_X1 U563 ( .A1(n412), .A2(n736), .ZN(G63) );
  BUF_X2 U564 ( .A(n377), .Z(n413) );
  NAND2_X1 U565 ( .A1(n727), .A2(G475), .ZN(n728) );
  AND2_X2 U566 ( .A1(n686), .A2(n685), .ZN(n727) );
  XNOR2_X1 U567 ( .A(n468), .B(n498), .ZN(n605) );
  XNOR2_X1 U568 ( .A(n728), .B(n729), .ZN(n415) );
  NAND2_X1 U569 ( .A1(n454), .A2(n453), .ZN(n458) );
  XNOR2_X1 U570 ( .A(n588), .B(n419), .ZN(n589) );
  NAND2_X1 U571 ( .A1(n501), .A2(n500), .ZN(n588) );
  NAND2_X1 U572 ( .A1(n699), .A2(n763), .ZN(n562) );
  NOR2_X2 U573 ( .A1(n605), .A2(n503), .ZN(n504) );
  XNOR2_X1 U574 ( .A(n614), .B(n424), .ZN(n423) );
  NAND2_X1 U575 ( .A1(n596), .A2(n659), .ZN(n598) );
  INV_X1 U576 ( .A(n733), .ZN(n428) );
  NAND2_X1 U577 ( .A1(n727), .A2(n432), .ZN(n431) );
  AND2_X1 U578 ( .A1(n687), .A2(G472), .ZN(n432) );
  XNOR2_X1 U579 ( .A(n433), .B(n689), .ZN(G57) );
  NAND2_X1 U580 ( .A1(n435), .A2(n659), .ZN(n468) );
  XNOR2_X2 U581 ( .A(n495), .B(n362), .ZN(n435) );
  NOR2_X1 U582 ( .A1(n662), .A2(n438), .ZN(n437) );
  NAND2_X1 U583 ( .A1(n443), .A2(n442), .ZN(n441) );
  INV_X1 U584 ( .A(KEYINPUT66), .ZN(n444) );
  XNOR2_X1 U585 ( .A(n446), .B(n445), .ZN(n615) );
  INV_X1 U586 ( .A(KEYINPUT76), .ZN(n445) );
  NAND2_X1 U587 ( .A1(n542), .A2(G221), .ZN(n543) );
  INV_X1 U588 ( .A(KEYINPUT71), .ZN(n452) );
  OR2_X1 U589 ( .A1(n643), .A2(n567), .ZN(n453) );
  NOR2_X1 U590 ( .A1(n578), .A2(n567), .ZN(n456) );
  AND2_X1 U591 ( .A1(n578), .A2(n567), .ZN(n457) );
  XNOR2_X1 U592 ( .A(n616), .B(KEYINPUT75), .ZN(n460) );
  XNOR2_X1 U593 ( .A(n621), .B(KEYINPUT36), .ZN(n462) );
  NOR2_X1 U594 ( .A1(n620), .A2(n464), .ZN(n463) );
  XNOR2_X1 U595 ( .A(n471), .B(n720), .ZN(G51) );
  XNOR2_X1 U596 ( .A(n719), .B(n718), .ZN(n473) );
  INV_X1 U597 ( .A(KEYINPUT48), .ZN(n622) );
  INV_X1 U598 ( .A(KEYINPUT4), .ZN(n474) );
  XNOR2_X1 U599 ( .A(n622), .B(KEYINPUT82), .ZN(n623) );
  XNOR2_X1 U600 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U601 ( .A(n587), .B(n586), .ZN(n636) );
  INV_X1 U602 ( .A(n411), .ZN(n558) );
  XNOR2_X1 U603 ( .A(n547), .B(n546), .ZN(n548) );
  INV_X1 U604 ( .A(KEYINPUT87), .ZN(n496) );
  INV_X1 U605 ( .A(G472), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n548), .B(n549), .ZN(n552) );
  XNOR2_X1 U607 ( .A(KEYINPUT53), .B(KEYINPUT119), .ZN(n680) );
  XNOR2_X1 U608 ( .A(n681), .B(n680), .ZN(G75) );
  NOR2_X1 U609 ( .A1(KEYINPUT44), .A2(KEYINPUT83), .ZN(n563) );
  XNOR2_X1 U610 ( .A(G134), .B(KEYINPUT65), .ZN(n475) );
  XNOR2_X1 U611 ( .A(n475), .B(G131), .ZN(n476) );
  XOR2_X1 U612 ( .A(n551), .B(G110), .Z(n477) );
  NAND2_X1 U613 ( .A1(G227), .A2(n377), .ZN(n479) );
  XNOR2_X1 U614 ( .A(KEYINPUT1), .B(KEYINPUT64), .ZN(n483) );
  NAND2_X1 U615 ( .A1(G224), .A2(n413), .ZN(n488) );
  XOR2_X1 U616 ( .A(G113), .B(n490), .Z(n539) );
  XOR2_X1 U617 ( .A(KEYINPUT16), .B(n545), .Z(n492) );
  XNOR2_X1 U618 ( .A(n507), .B(n521), .ZN(n491) );
  XNOR2_X1 U619 ( .A(n492), .B(n491), .ZN(n493) );
  NAND2_X1 U620 ( .A1(n719), .A2(n683), .ZN(n495) );
  AND2_X1 U621 ( .A1(G210), .A2(n497), .ZN(n494) );
  INV_X1 U622 ( .A(KEYINPUT19), .ZN(n498) );
  NAND2_X1 U623 ( .A1(G952), .A2(n501), .ZN(n675) );
  NOR2_X1 U624 ( .A1(G953), .A2(n675), .ZN(n592) );
  NOR2_X1 U625 ( .A1(G898), .A2(n588), .ZN(n502) );
  NOR2_X1 U626 ( .A1(n592), .A2(n502), .ZN(n503) );
  XNOR2_X1 U627 ( .A(KEYINPUT10), .B(n506), .ZN(n550) );
  XNOR2_X1 U628 ( .A(n507), .B(KEYINPUT12), .ZN(n511) );
  XOR2_X1 U629 ( .A(KEYINPUT11), .B(KEYINPUT98), .Z(n509) );
  XNOR2_X1 U630 ( .A(KEYINPUT96), .B(KEYINPUT97), .ZN(n508) );
  XNOR2_X1 U631 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U632 ( .A(n513), .B(n512), .ZN(n515) );
  NOR2_X1 U633 ( .A1(G953), .A2(G237), .ZN(n531) );
  NAND2_X1 U634 ( .A1(G214), .A2(n531), .ZN(n514) );
  XNOR2_X1 U635 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U636 ( .A(KEYINPUT13), .B(KEYINPUT99), .ZN(n517) );
  XOR2_X1 U637 ( .A(n518), .B(KEYINPUT9), .Z(n520) );
  NAND2_X1 U638 ( .A1(G217), .A2(n542), .ZN(n519) );
  XNOR2_X1 U639 ( .A(n520), .B(n519), .ZN(n522) );
  XOR2_X1 U640 ( .A(KEYINPUT7), .B(KEYINPUT101), .Z(n523) );
  XNOR2_X1 U641 ( .A(n524), .B(n523), .ZN(n732) );
  NOR2_X1 U642 ( .A1(G902), .A2(n732), .ZN(n526) );
  XNOR2_X1 U643 ( .A(KEYINPUT102), .B(G478), .ZN(n525) );
  NAND2_X1 U644 ( .A1(n571), .A2(n572), .ZN(n527) );
  XNOR2_X1 U645 ( .A(n527), .B(KEYINPUT104), .ZN(n662) );
  XOR2_X1 U646 ( .A(KEYINPUT92), .B(KEYINPUT21), .Z(n530) );
  NAND2_X1 U647 ( .A1(n683), .A2(G234), .ZN(n528) );
  XNOR2_X1 U648 ( .A(n528), .B(KEYINPUT20), .ZN(n553) );
  NAND2_X1 U649 ( .A1(G221), .A2(n553), .ZN(n529) );
  XNOR2_X1 U650 ( .A(n530), .B(n529), .ZN(n644) );
  XOR2_X1 U651 ( .A(G116), .B(KEYINPUT93), .Z(n533) );
  NAND2_X1 U652 ( .A1(G210), .A2(n531), .ZN(n532) );
  XNOR2_X1 U653 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U654 ( .A(n534), .B(KEYINPUT5), .Z(n536) );
  XNOR2_X1 U655 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U656 ( .A(G128), .B(KEYINPUT24), .Z(n544) );
  XNOR2_X1 U657 ( .A(n544), .B(n543), .ZN(n549) );
  XNOR2_X1 U658 ( .A(n545), .B(KEYINPUT90), .ZN(n547) );
  XNOR2_X1 U659 ( .A(n551), .B(n550), .ZN(n749) );
  NAND2_X1 U660 ( .A1(G217), .A2(n553), .ZN(n554) );
  XNOR2_X1 U661 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U662 ( .A(KEYINPUT91), .B(n556), .ZN(n557) );
  XNOR2_X1 U663 ( .A(n563), .B(n562), .ZN(n569) );
  NAND2_X1 U664 ( .A1(n644), .A2(n645), .ZN(n650) );
  NOR2_X1 U665 ( .A1(n649), .A2(n650), .ZN(n564) );
  XOR2_X1 U666 ( .A(KEYINPUT84), .B(KEYINPUT33), .Z(n565) );
  NOR2_X1 U667 ( .A1(n572), .A2(n571), .ZN(n612) );
  INV_X1 U668 ( .A(KEYINPUT35), .ZN(n568) );
  NAND2_X1 U669 ( .A1(n569), .A2(n762), .ZN(n570) );
  NOR2_X1 U670 ( .A1(n572), .A2(n573), .ZN(n710) );
  NAND2_X1 U671 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U672 ( .A(KEYINPUT31), .B(KEYINPUT95), .Z(n577) );
  XNOR2_X1 U673 ( .A(n575), .B(KEYINPUT94), .ZN(n654) );
  XNOR2_X1 U674 ( .A(n577), .B(n576), .ZN(n711) );
  INV_X1 U675 ( .A(n606), .ZN(n600) );
  INV_X1 U676 ( .A(n650), .ZN(n599) );
  AND2_X1 U677 ( .A1(n600), .A2(n599), .ZN(n579) );
  NAND2_X1 U678 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U679 ( .A1(n451), .A2(n580), .ZN(n696) );
  NOR2_X1 U680 ( .A1(n711), .A2(n696), .ZN(n581) );
  NOR2_X1 U681 ( .A1(n664), .A2(n581), .ZN(n584) );
  INV_X1 U682 ( .A(n582), .ZN(n619) );
  NAND2_X1 U683 ( .A1(n411), .A2(n363), .ZN(n583) );
  NOR2_X1 U684 ( .A1(n619), .A2(n583), .ZN(n690) );
  NOR2_X1 U685 ( .A1(n584), .A2(n690), .ZN(n585) );
  INV_X1 U686 ( .A(n636), .ZN(n737) );
  NAND2_X1 U687 ( .A1(KEYINPUT77), .A2(n737), .ZN(n632) );
  NOR2_X1 U688 ( .A1(G900), .A2(n589), .ZN(n590) );
  XNOR2_X1 U689 ( .A(n590), .B(KEYINPUT106), .ZN(n591) );
  NAND2_X1 U690 ( .A1(n608), .A2(n600), .ZN(n594) );
  NAND2_X1 U691 ( .A1(n660), .A2(n659), .ZN(n665) );
  XNOR2_X1 U692 ( .A(n593), .B(KEYINPUT41), .ZN(n658) );
  NOR2_X1 U693 ( .A1(n594), .A2(n658), .ZN(n595) );
  XNOR2_X1 U694 ( .A(KEYINPUT42), .B(n595), .ZN(n765) );
  XNOR2_X1 U695 ( .A(KEYINPUT30), .B(KEYINPUT107), .ZN(n597) );
  XNOR2_X1 U696 ( .A(n598), .B(n597), .ZN(n601) );
  NAND2_X1 U697 ( .A1(n609), .A2(n660), .ZN(n602) );
  XNOR2_X1 U698 ( .A(n602), .B(KEYINPUT39), .ZN(n624) );
  AND2_X1 U699 ( .A1(n624), .A2(n707), .ZN(n603) );
  XNOR2_X1 U700 ( .A(KEYINPUT40), .B(n603), .ZN(n764) );
  NOR2_X1 U701 ( .A1(n765), .A2(n764), .ZN(n604) );
  NOR2_X1 U702 ( .A1(n606), .A2(n605), .ZN(n607) );
  NAND2_X1 U703 ( .A1(KEYINPUT47), .A2(n664), .ZN(n613) );
  INV_X1 U704 ( .A(KEYINPUT108), .ZN(n611) );
  NOR2_X1 U705 ( .A1(n664), .A2(KEYINPUT47), .ZN(n617) );
  NAND2_X1 U706 ( .A1(n705), .A2(n617), .ZN(n618) );
  NOR2_X1 U707 ( .A1(n629), .A2(n627), .ZN(n621) );
  NAND2_X1 U708 ( .A1(n710), .A2(n624), .ZN(n625) );
  XNOR2_X1 U709 ( .A(n625), .B(KEYINPUT109), .ZN(n761) );
  OR2_X1 U710 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U711 ( .A(n628), .B(KEYINPUT43), .ZN(n630) );
  NAND2_X1 U712 ( .A1(n630), .A2(n629), .ZN(n716) );
  NAND2_X1 U713 ( .A1(n637), .A2(n716), .ZN(n752) );
  INV_X1 U714 ( .A(KEYINPUT2), .ZN(n631) );
  NOR2_X1 U715 ( .A1(KEYINPUT78), .A2(n752), .ZN(n633) );
  INV_X1 U716 ( .A(n716), .ZN(n635) );
  NOR2_X1 U717 ( .A1(n636), .A2(n635), .ZN(n638) );
  NAND2_X1 U718 ( .A1(KEYINPUT78), .A2(n639), .ZN(n640) );
  NAND2_X1 U719 ( .A1(KEYINPUT2), .A2(n640), .ZN(n641) );
  INV_X1 U720 ( .A(n643), .ZN(n669) );
  NOR2_X1 U721 ( .A1(n669), .A2(n658), .ZN(n678) );
  XOR2_X1 U722 ( .A(KEYINPUT52), .B(KEYINPUT117), .Z(n673) );
  NOR2_X1 U723 ( .A1(n411), .A2(n644), .ZN(n646) );
  XNOR2_X1 U724 ( .A(n646), .B(KEYINPUT49), .ZN(n647) );
  NAND2_X1 U725 ( .A1(n416), .A2(n647), .ZN(n653) );
  NAND2_X1 U726 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U727 ( .A(KEYINPUT50), .B(n651), .Z(n652) );
  NOR2_X1 U728 ( .A1(n653), .A2(n652), .ZN(n655) );
  NOR2_X1 U729 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U730 ( .A(KEYINPUT51), .B(n656), .Z(n657) );
  NOR2_X1 U731 ( .A1(n658), .A2(n657), .ZN(n671) );
  NOR2_X1 U732 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U733 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U734 ( .A(n663), .B(KEYINPUT116), .ZN(n667) );
  NOR2_X1 U735 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U736 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U737 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U738 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U739 ( .A(n673), .B(n672), .ZN(n674) );
  NOR2_X1 U740 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U741 ( .A(n676), .B(KEYINPUT118), .ZN(n677) );
  NOR2_X1 U742 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U743 ( .A(KEYINPUT63), .B(KEYINPUT85), .Z(n689) );
  XOR2_X1 U744 ( .A(n682), .B(KEYINPUT62), .Z(n687) );
  XNOR2_X1 U745 ( .A(n684), .B(n683), .ZN(n686) );
  NOR2_X1 U746 ( .A1(G952), .A2(n413), .ZN(n688) );
  XOR2_X1 U747 ( .A(G101), .B(n690), .Z(G3) );
  NAND2_X1 U748 ( .A1(n696), .A2(n707), .ZN(n691) );
  XNOR2_X1 U749 ( .A(n691), .B(KEYINPUT110), .ZN(n692) );
  XNOR2_X1 U750 ( .A(G104), .B(n692), .ZN(G6) );
  XOR2_X1 U751 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n694) );
  XNOR2_X1 U752 ( .A(G107), .B(KEYINPUT26), .ZN(n693) );
  XNOR2_X1 U753 ( .A(n694), .B(n693), .ZN(n695) );
  XOR2_X1 U754 ( .A(KEYINPUT27), .B(n695), .Z(n698) );
  NAND2_X1 U755 ( .A1(n696), .A2(n710), .ZN(n697) );
  XNOR2_X1 U756 ( .A(n698), .B(n697), .ZN(G9) );
  XNOR2_X1 U757 ( .A(n699), .B(G110), .ZN(G12) );
  XOR2_X1 U758 ( .A(KEYINPUT113), .B(KEYINPUT29), .Z(n701) );
  NAND2_X1 U759 ( .A1(n705), .A2(n710), .ZN(n700) );
  XNOR2_X1 U760 ( .A(n701), .B(n700), .ZN(n702) );
  XOR2_X1 U761 ( .A(G128), .B(n702), .Z(G30) );
  BUF_X1 U762 ( .A(n703), .Z(n704) );
  XNOR2_X1 U763 ( .A(G143), .B(n704), .ZN(G45) );
  NAND2_X1 U764 ( .A1(n705), .A2(n707), .ZN(n706) );
  XNOR2_X1 U765 ( .A(n706), .B(G146), .ZN(G48) );
  NAND2_X1 U766 ( .A1(n711), .A2(n707), .ZN(n708) );
  XNOR2_X1 U767 ( .A(n708), .B(KEYINPUT114), .ZN(n709) );
  XNOR2_X1 U768 ( .A(G113), .B(n709), .ZN(G15) );
  XOR2_X1 U769 ( .A(G116), .B(KEYINPUT115), .Z(n713) );
  NAND2_X1 U770 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U771 ( .A(n713), .B(n712), .ZN(G18) );
  XNOR2_X1 U772 ( .A(G125), .B(n714), .ZN(n715) );
  XNOR2_X1 U773 ( .A(n715), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U774 ( .A(G140), .B(n716), .ZN(G42) );
  XOR2_X1 U775 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n718) );
  NAND2_X1 U776 ( .A1(n727), .A2(G210), .ZN(n717) );
  XOR2_X1 U777 ( .A(KEYINPUT56), .B(KEYINPUT120), .Z(n720) );
  INV_X1 U778 ( .A(n730), .ZN(n736) );
  XNOR2_X1 U779 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n723) );
  XNOR2_X1 U780 ( .A(n721), .B(KEYINPUT57), .ZN(n722) );
  XNOR2_X1 U781 ( .A(n723), .B(n722), .ZN(n725) );
  NAND2_X1 U782 ( .A1(n733), .A2(G469), .ZN(n724) );
  NAND2_X1 U783 ( .A1(G478), .A2(n733), .ZN(n731) );
  NAND2_X1 U784 ( .A1(G217), .A2(n733), .ZN(n734) );
  NAND2_X1 U785 ( .A1(n737), .A2(n413), .ZN(n738) );
  XNOR2_X1 U786 ( .A(n738), .B(KEYINPUT122), .ZN(n742) );
  NAND2_X1 U787 ( .A1(G953), .A2(G224), .ZN(n739) );
  XNOR2_X1 U788 ( .A(KEYINPUT61), .B(n739), .ZN(n740) );
  NAND2_X1 U789 ( .A1(n740), .A2(G898), .ZN(n741) );
  NAND2_X1 U790 ( .A1(n742), .A2(n741), .ZN(n747) );
  NOR2_X1 U791 ( .A1(G898), .A2(n413), .ZN(n743) );
  NOR2_X1 U792 ( .A1(n744), .A2(n743), .ZN(n745) );
  XOR2_X1 U793 ( .A(KEYINPUT123), .B(n745), .Z(n746) );
  XNOR2_X1 U794 ( .A(n747), .B(n746), .ZN(G69) );
  XNOR2_X1 U795 ( .A(KEYINPUT124), .B(n748), .ZN(n750) );
  XOR2_X1 U796 ( .A(n750), .B(n749), .Z(n755) );
  XOR2_X1 U797 ( .A(n755), .B(KEYINPUT125), .Z(n751) );
  XNOR2_X1 U798 ( .A(n752), .B(n751), .ZN(n753) );
  NAND2_X1 U799 ( .A1(n413), .A2(n753), .ZN(n754) );
  XNOR2_X1 U800 ( .A(n754), .B(KEYINPUT126), .ZN(n759) );
  XNOR2_X1 U801 ( .A(G227), .B(n755), .ZN(n756) );
  NAND2_X1 U802 ( .A1(n756), .A2(G900), .ZN(n757) );
  NAND2_X1 U803 ( .A1(G953), .A2(n757), .ZN(n758) );
  NAND2_X1 U804 ( .A1(n759), .A2(n758), .ZN(n760) );
  XOR2_X1 U805 ( .A(KEYINPUT127), .B(n760), .Z(G72) );
  XOR2_X1 U806 ( .A(G134), .B(n761), .Z(G36) );
  XNOR2_X1 U807 ( .A(n762), .B(G122), .ZN(G24) );
  XNOR2_X1 U808 ( .A(G119), .B(n763), .ZN(G21) );
  XOR2_X1 U809 ( .A(G131), .B(n764), .Z(G33) );
  XOR2_X1 U810 ( .A(G137), .B(n765), .Z(G39) );
endmodule

