

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579;

  XNOR2_X1 U322 ( .A(n327), .B(n326), .ZN(n555) );
  XOR2_X1 U323 ( .A(G92GAT), .B(G85GAT), .Z(n290) );
  XOR2_X1 U324 ( .A(n366), .B(n431), .Z(n291) );
  XOR2_X1 U325 ( .A(KEYINPUT36), .B(n540), .Z(n576) );
  XNOR2_X1 U326 ( .A(n325), .B(n324), .ZN(n326) );
  NOR2_X1 U327 ( .A1(n529), .A2(n444), .ZN(n559) );
  XNOR2_X1 U328 ( .A(n449), .B(G190GAT), .ZN(n450) );
  XNOR2_X1 U329 ( .A(n451), .B(n450), .ZN(G1351GAT) );
  XOR2_X1 U330 ( .A(G127GAT), .B(G134GAT), .Z(n293) );
  XNOR2_X1 U331 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n292) );
  XNOR2_X1 U332 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U333 ( .A(G113GAT), .B(n294), .Z(n413) );
  XOR2_X1 U334 ( .A(G15GAT), .B(G183GAT), .Z(n296) );
  NAND2_X1 U335 ( .A1(G227GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U336 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U337 ( .A(n297), .B(G190GAT), .Z(n302) );
  XOR2_X1 U338 ( .A(KEYINPUT82), .B(KEYINPUT17), .Z(n299) );
  XNOR2_X1 U339 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n298) );
  XNOR2_X1 U340 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U341 ( .A(G169GAT), .B(n300), .Z(n396) );
  XNOR2_X1 U342 ( .A(G43GAT), .B(n396), .ZN(n301) );
  XNOR2_X1 U343 ( .A(n302), .B(n301), .ZN(n310) );
  XOR2_X1 U344 ( .A(G71GAT), .B(G176GAT), .Z(n304) );
  XNOR2_X1 U345 ( .A(KEYINPUT20), .B(KEYINPUT81), .ZN(n303) );
  XNOR2_X1 U346 ( .A(n304), .B(n303), .ZN(n308) );
  XOR2_X1 U347 ( .A(KEYINPUT65), .B(KEYINPUT80), .Z(n306) );
  XNOR2_X1 U348 ( .A(G99GAT), .B(KEYINPUT83), .ZN(n305) );
  XNOR2_X1 U349 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U350 ( .A(n308), .B(n307), .Z(n309) );
  XNOR2_X1 U351 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U352 ( .A(n413), .B(n311), .ZN(n529) );
  XNOR2_X1 U353 ( .A(G99GAT), .B(G106GAT), .ZN(n312) );
  XNOR2_X1 U354 ( .A(n290), .B(n312), .ZN(n366) );
  XOR2_X1 U355 ( .A(G50GAT), .B(G162GAT), .Z(n431) );
  NAND2_X1 U356 ( .A1(G232GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U357 ( .A(n291), .B(n313), .ZN(n317) );
  XOR2_X1 U358 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n315) );
  XNOR2_X1 U359 ( .A(KEYINPUT11), .B(KEYINPUT75), .ZN(n314) );
  XNOR2_X1 U360 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U361 ( .A(n317), .B(n316), .Z(n327) );
  XOR2_X1 U362 ( .A(G29GAT), .B(G43GAT), .Z(n319) );
  XNOR2_X1 U363 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n318) );
  XNOR2_X1 U364 ( .A(n319), .B(n318), .ZN(n348) );
  XOR2_X1 U365 ( .A(KEYINPUT74), .B(G218GAT), .Z(n321) );
  XNOR2_X1 U366 ( .A(G36GAT), .B(G190GAT), .ZN(n320) );
  XNOR2_X1 U367 ( .A(n321), .B(n320), .ZN(n393) );
  XNOR2_X1 U368 ( .A(n348), .B(n393), .ZN(n325) );
  XOR2_X1 U369 ( .A(KEYINPUT73), .B(KEYINPUT64), .Z(n323) );
  XNOR2_X1 U370 ( .A(G134GAT), .B(KEYINPUT72), .ZN(n322) );
  XNOR2_X1 U371 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U372 ( .A(G15GAT), .B(G1GAT), .Z(n328) );
  XNOR2_X1 U373 ( .A(KEYINPUT67), .B(n328), .ZN(n347) );
  INV_X1 U374 ( .A(n347), .ZN(n330) );
  XNOR2_X1 U375 ( .A(G8GAT), .B(G183GAT), .ZN(n329) );
  XNOR2_X1 U376 ( .A(n329), .B(G211GAT), .ZN(n388) );
  XNOR2_X1 U377 ( .A(n330), .B(n388), .ZN(n346) );
  XOR2_X1 U378 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n332) );
  XNOR2_X1 U379 ( .A(G64GAT), .B(KEYINPUT15), .ZN(n331) );
  XNOR2_X1 U380 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U381 ( .A(n333), .B(G78GAT), .Z(n335) );
  XOR2_X1 U382 ( .A(G22GAT), .B(G155GAT), .Z(n428) );
  XNOR2_X1 U383 ( .A(G127GAT), .B(n428), .ZN(n334) );
  XNOR2_X1 U384 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U385 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n337) );
  NAND2_X1 U386 ( .A1(G231GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U387 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U388 ( .A(n339), .B(n338), .Z(n344) );
  XOR2_X1 U389 ( .A(KEYINPUT70), .B(KEYINPUT13), .Z(n341) );
  XNOR2_X1 U390 ( .A(G71GAT), .B(G57GAT), .ZN(n340) );
  XNOR2_X1 U391 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U392 ( .A(KEYINPUT69), .B(n342), .ZN(n372) );
  XOR2_X1 U393 ( .A(n372), .B(KEYINPUT77), .Z(n343) );
  XNOR2_X1 U394 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U395 ( .A(n346), .B(n345), .ZN(n571) );
  XNOR2_X1 U396 ( .A(n571), .B(KEYINPUT112), .ZN(n560) );
  XNOR2_X1 U397 ( .A(n348), .B(n347), .ZN(n361) );
  XOR2_X1 U398 ( .A(KEYINPUT68), .B(KEYINPUT29), .Z(n350) );
  NAND2_X1 U399 ( .A1(G229GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U400 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U401 ( .A(n351), .B(KEYINPUT30), .Z(n359) );
  XOR2_X1 U402 ( .A(G141GAT), .B(G197GAT), .Z(n353) );
  XNOR2_X1 U403 ( .A(G36GAT), .B(G50GAT), .ZN(n352) );
  XNOR2_X1 U404 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U405 ( .A(G8GAT), .B(G113GAT), .Z(n355) );
  XNOR2_X1 U406 ( .A(G169GAT), .B(G22GAT), .ZN(n354) );
  XNOR2_X1 U407 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U408 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U409 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U410 ( .A(n361), .B(n360), .ZN(n564) );
  INV_X1 U411 ( .A(n564), .ZN(n452) );
  XOR2_X1 U412 ( .A(KEYINPUT71), .B(KEYINPUT32), .Z(n363) );
  NAND2_X1 U413 ( .A1(G230GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U414 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U415 ( .A(n364), .B(KEYINPUT33), .Z(n368) );
  XNOR2_X1 U416 ( .A(G176GAT), .B(G204GAT), .ZN(n365) );
  XNOR2_X1 U417 ( .A(n365), .B(G64GAT), .ZN(n390) );
  XNOR2_X1 U418 ( .A(n366), .B(n390), .ZN(n367) );
  XNOR2_X1 U419 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U420 ( .A(n369), .B(KEYINPUT31), .Z(n371) );
  XOR2_X1 U421 ( .A(G148GAT), .B(G78GAT), .Z(n427) );
  XNOR2_X1 U422 ( .A(G120GAT), .B(n427), .ZN(n370) );
  XNOR2_X1 U423 ( .A(n371), .B(n370), .ZN(n373) );
  XNOR2_X1 U424 ( .A(n373), .B(n372), .ZN(n568) );
  XNOR2_X1 U425 ( .A(n568), .B(KEYINPUT41), .ZN(n503) );
  NOR2_X1 U426 ( .A1(n452), .A2(n503), .ZN(n374) );
  XNOR2_X1 U427 ( .A(n374), .B(KEYINPUT46), .ZN(n375) );
  NOR2_X1 U428 ( .A1(n560), .A2(n375), .ZN(n376) );
  XNOR2_X1 U429 ( .A(n376), .B(KEYINPUT113), .ZN(n377) );
  NOR2_X1 U430 ( .A1(n555), .A2(n377), .ZN(n378) );
  XNOR2_X1 U431 ( .A(n378), .B(KEYINPUT47), .ZN(n383) );
  XNOR2_X1 U432 ( .A(KEYINPUT76), .B(n555), .ZN(n540) );
  INV_X1 U433 ( .A(n571), .ZN(n486) );
  NOR2_X1 U434 ( .A1(n576), .A2(n486), .ZN(n379) );
  XOR2_X1 U435 ( .A(KEYINPUT45), .B(n379), .Z(n380) );
  NOR2_X1 U436 ( .A1(n568), .A2(n380), .ZN(n381) );
  NAND2_X1 U437 ( .A1(n381), .A2(n452), .ZN(n382) );
  NAND2_X1 U438 ( .A1(n383), .A2(n382), .ZN(n385) );
  XNOR2_X1 U439 ( .A(KEYINPUT114), .B(KEYINPUT48), .ZN(n384) );
  XNOR2_X1 U440 ( .A(n385), .B(n384), .ZN(n527) );
  XOR2_X1 U441 ( .A(KEYINPUT94), .B(KEYINPUT93), .Z(n387) );
  NAND2_X1 U442 ( .A1(G226GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U443 ( .A(n387), .B(n386), .ZN(n389) );
  XOR2_X1 U444 ( .A(n389), .B(n388), .Z(n392) );
  XNOR2_X1 U445 ( .A(G92GAT), .B(n390), .ZN(n391) );
  XNOR2_X1 U446 ( .A(n392), .B(n391), .ZN(n394) );
  XOR2_X1 U447 ( .A(n394), .B(n393), .Z(n398) );
  XOR2_X1 U448 ( .A(G197GAT), .B(KEYINPUT21), .Z(n395) );
  XOR2_X1 U449 ( .A(KEYINPUT85), .B(n395), .Z(n425) );
  XNOR2_X1 U450 ( .A(n396), .B(n425), .ZN(n397) );
  XNOR2_X1 U451 ( .A(n398), .B(n397), .ZN(n475) );
  NAND2_X1 U452 ( .A1(n527), .A2(n475), .ZN(n401) );
  XNOR2_X1 U453 ( .A(KEYINPUT122), .B(KEYINPUT54), .ZN(n399) );
  XNOR2_X1 U454 ( .A(n399), .B(KEYINPUT121), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n401), .B(n400), .ZN(n424) );
  XOR2_X1 U456 ( .A(G57GAT), .B(KEYINPUT6), .Z(n403) );
  XNOR2_X1 U457 ( .A(KEYINPUT92), .B(KEYINPUT1), .ZN(n402) );
  XNOR2_X1 U458 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U459 ( .A(KEYINPUT5), .B(KEYINPUT90), .Z(n405) );
  XNOR2_X1 U460 ( .A(KEYINPUT91), .B(KEYINPUT89), .ZN(n404) );
  XNOR2_X1 U461 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U462 ( .A(n407), .B(n406), .Z(n415) );
  XOR2_X1 U463 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n409) );
  XNOR2_X1 U464 ( .A(G141GAT), .B(KEYINPUT86), .ZN(n408) );
  XNOR2_X1 U465 ( .A(n409), .B(n408), .ZN(n426) );
  XOR2_X1 U466 ( .A(n426), .B(KEYINPUT4), .Z(n411) );
  NAND2_X1 U467 ( .A1(G225GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U469 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U470 ( .A(n415), .B(n414), .ZN(n423) );
  XOR2_X1 U471 ( .A(KEYINPUT87), .B(KEYINPUT88), .Z(n417) );
  XNOR2_X1 U472 ( .A(G1GAT), .B(G148GAT), .ZN(n416) );
  XNOR2_X1 U473 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U474 ( .A(G85GAT), .B(G155GAT), .Z(n419) );
  XNOR2_X1 U475 ( .A(G29GAT), .B(G162GAT), .ZN(n418) );
  XNOR2_X1 U476 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U477 ( .A(n421), .B(n420), .Z(n422) );
  XNOR2_X1 U478 ( .A(n423), .B(n422), .ZN(n515) );
  NAND2_X1 U479 ( .A1(n424), .A2(n515), .ZN(n562) );
  XOR2_X1 U480 ( .A(n426), .B(n425), .Z(n442) );
  XOR2_X1 U481 ( .A(n428), .B(n427), .Z(n430) );
  NAND2_X1 U482 ( .A1(G228GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U483 ( .A(n430), .B(n429), .ZN(n432) );
  XOR2_X1 U484 ( .A(n432), .B(n431), .Z(n440) );
  XOR2_X1 U485 ( .A(KEYINPUT23), .B(KEYINPUT84), .Z(n434) );
  XNOR2_X1 U486 ( .A(G218GAT), .B(G106GAT), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U488 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n436) );
  XNOR2_X1 U489 ( .A(G211GAT), .B(G204GAT), .ZN(n435) );
  XNOR2_X1 U490 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U491 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U492 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U493 ( .A(n442), .B(n441), .ZN(n461) );
  NOR2_X1 U494 ( .A1(n562), .A2(n461), .ZN(n443) );
  XNOR2_X1 U495 ( .A(n443), .B(KEYINPUT55), .ZN(n444) );
  INV_X1 U496 ( .A(n503), .ZN(n546) );
  NAND2_X1 U497 ( .A1(n559), .A2(n546), .ZN(n448) );
  XOR2_X1 U498 ( .A(G176GAT), .B(KEYINPUT56), .Z(n446) );
  XNOR2_X1 U499 ( .A(KEYINPUT57), .B(KEYINPUT124), .ZN(n445) );
  XNOR2_X1 U500 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U501 ( .A(n448), .B(n447), .ZN(G1349GAT) );
  NAND2_X1 U502 ( .A1(n559), .A2(n540), .ZN(n451) );
  XOR2_X1 U503 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n449) );
  NOR2_X1 U504 ( .A1(n452), .A2(n568), .ZN(n488) );
  INV_X1 U505 ( .A(n515), .ZN(n472) );
  INV_X1 U506 ( .A(n475), .ZN(n517) );
  NOR2_X1 U507 ( .A1(n529), .A2(n517), .ZN(n453) );
  NOR2_X1 U508 ( .A1(n461), .A2(n453), .ZN(n454) );
  XOR2_X1 U509 ( .A(n454), .B(KEYINPUT98), .Z(n455) );
  XNOR2_X1 U510 ( .A(KEYINPUT25), .B(n455), .ZN(n459) );
  XOR2_X1 U511 ( .A(n475), .B(KEYINPUT27), .Z(n463) );
  XOR2_X1 U512 ( .A(KEYINPUT97), .B(KEYINPUT26), .Z(n457) );
  NAND2_X1 U513 ( .A1(n529), .A2(n461), .ZN(n456) );
  XNOR2_X1 U514 ( .A(n457), .B(n456), .ZN(n563) );
  NOR2_X1 U515 ( .A1(n463), .A2(n563), .ZN(n458) );
  NOR2_X1 U516 ( .A1(n459), .A2(n458), .ZN(n460) );
  NOR2_X1 U517 ( .A1(n472), .A2(n460), .ZN(n468) );
  XNOR2_X1 U518 ( .A(KEYINPUT28), .B(KEYINPUT66), .ZN(n462) );
  XNOR2_X1 U519 ( .A(n462), .B(n461), .ZN(n532) );
  NOR2_X1 U520 ( .A1(n463), .A2(n515), .ZN(n464) );
  XOR2_X1 U521 ( .A(KEYINPUT95), .B(n464), .Z(n528) );
  NAND2_X1 U522 ( .A1(n529), .A2(n528), .ZN(n465) );
  NOR2_X1 U523 ( .A1(n532), .A2(n465), .ZN(n466) );
  XNOR2_X1 U524 ( .A(n466), .B(KEYINPUT96), .ZN(n467) );
  NOR2_X1 U525 ( .A1(n468), .A2(n467), .ZN(n484) );
  NOR2_X1 U526 ( .A1(n540), .A2(n486), .ZN(n469) );
  XOR2_X1 U527 ( .A(KEYINPUT16), .B(n469), .Z(n470) );
  NOR2_X1 U528 ( .A1(n484), .A2(n470), .ZN(n504) );
  NAND2_X1 U529 ( .A1(n488), .A2(n504), .ZN(n471) );
  XNOR2_X1 U530 ( .A(KEYINPUT99), .B(n471), .ZN(n482) );
  NAND2_X1 U531 ( .A1(n482), .A2(n472), .ZN(n473) );
  XNOR2_X1 U532 ( .A(n473), .B(KEYINPUT34), .ZN(n474) );
  XNOR2_X1 U533 ( .A(G1GAT), .B(n474), .ZN(G1324GAT) );
  NAND2_X1 U534 ( .A1(n482), .A2(n475), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n476), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U536 ( .A(G15GAT), .B(KEYINPUT100), .Z(n479) );
  INV_X1 U537 ( .A(n529), .ZN(n477) );
  NAND2_X1 U538 ( .A1(n482), .A2(n477), .ZN(n478) );
  XNOR2_X1 U539 ( .A(n479), .B(n478), .ZN(n481) );
  XOR2_X1 U540 ( .A(KEYINPUT35), .B(KEYINPUT101), .Z(n480) );
  XNOR2_X1 U541 ( .A(n481), .B(n480), .ZN(G1326GAT) );
  NAND2_X1 U542 ( .A1(n532), .A2(n482), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n483), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U544 ( .A1(n576), .A2(n484), .ZN(n485) );
  NAND2_X1 U545 ( .A1(n486), .A2(n485), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n487), .B(KEYINPUT37), .ZN(n514) );
  NAND2_X1 U547 ( .A1(n488), .A2(n514), .ZN(n489) );
  XNOR2_X1 U548 ( .A(n489), .B(KEYINPUT38), .ZN(n498) );
  NOR2_X1 U549 ( .A1(n498), .A2(n515), .ZN(n491) );
  XNOR2_X1 U550 ( .A(KEYINPUT39), .B(KEYINPUT102), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U552 ( .A(G29GAT), .B(n492), .ZN(G1328GAT) );
  NOR2_X1 U553 ( .A1(n498), .A2(n517), .ZN(n493) );
  XOR2_X1 U554 ( .A(G36GAT), .B(n493), .Z(G1329GAT) );
  XOR2_X1 U555 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n495) );
  XNOR2_X1 U556 ( .A(G43GAT), .B(KEYINPUT103), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n495), .B(n494), .ZN(n497) );
  NOR2_X1 U558 ( .A1(n529), .A2(n498), .ZN(n496) );
  XOR2_X1 U559 ( .A(n497), .B(n496), .Z(G1330GAT) );
  XNOR2_X1 U560 ( .A(G50GAT), .B(KEYINPUT105), .ZN(n500) );
  INV_X1 U561 ( .A(n532), .ZN(n523) );
  NOR2_X1 U562 ( .A1(n523), .A2(n498), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n500), .B(n499), .ZN(G1331GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT107), .B(KEYINPUT42), .Z(n502) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(KEYINPUT106), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n502), .B(n501), .ZN(n506) );
  NOR2_X1 U567 ( .A1(n564), .A2(n503), .ZN(n513) );
  NAND2_X1 U568 ( .A1(n504), .A2(n513), .ZN(n510) );
  NOR2_X1 U569 ( .A1(n515), .A2(n510), .ZN(n505) );
  XOR2_X1 U570 ( .A(n506), .B(n505), .Z(G1332GAT) );
  NOR2_X1 U571 ( .A1(n517), .A2(n510), .ZN(n507) );
  XOR2_X1 U572 ( .A(KEYINPUT108), .B(n507), .Z(n508) );
  XNOR2_X1 U573 ( .A(G64GAT), .B(n508), .ZN(G1333GAT) );
  NOR2_X1 U574 ( .A1(n529), .A2(n510), .ZN(n509) );
  XOR2_X1 U575 ( .A(G71GAT), .B(n509), .Z(G1334GAT) );
  NOR2_X1 U576 ( .A1(n523), .A2(n510), .ZN(n512) );
  XNOR2_X1 U577 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n512), .B(n511), .ZN(G1335GAT) );
  NAND2_X1 U579 ( .A1(n514), .A2(n513), .ZN(n522) );
  NOR2_X1 U580 ( .A1(n515), .A2(n522), .ZN(n516) );
  XOR2_X1 U581 ( .A(G85GAT), .B(n516), .Z(G1336GAT) );
  NOR2_X1 U582 ( .A1(n517), .A2(n522), .ZN(n518) );
  XOR2_X1 U583 ( .A(G92GAT), .B(n518), .Z(G1337GAT) );
  NOR2_X1 U584 ( .A1(n529), .A2(n522), .ZN(n520) );
  XNOR2_X1 U585 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U587 ( .A(G99GAT), .B(n521), .ZN(G1338GAT) );
  NOR2_X1 U588 ( .A1(n523), .A2(n522), .ZN(n525) );
  XNOR2_X1 U589 ( .A(KEYINPUT111), .B(KEYINPUT44), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  NAND2_X1 U592 ( .A1(n528), .A2(n527), .ZN(n544) );
  NOR2_X1 U593 ( .A1(n529), .A2(n544), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n530), .B(KEYINPUT115), .ZN(n531) );
  NOR2_X1 U595 ( .A1(n532), .A2(n531), .ZN(n541) );
  NAND2_X1 U596 ( .A1(n564), .A2(n541), .ZN(n533) );
  XNOR2_X1 U597 ( .A(n533), .B(KEYINPUT116), .ZN(n534) );
  XNOR2_X1 U598 ( .A(G113GAT), .B(n534), .ZN(G1340GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n536) );
  NAND2_X1 U600 ( .A1(n541), .A2(n546), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U602 ( .A(G120GAT), .B(n537), .Z(G1341GAT) );
  NAND2_X1 U603 ( .A1(n560), .A2(n541), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n538), .B(KEYINPUT50), .ZN(n539) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(n539), .ZN(G1342GAT) );
  XOR2_X1 U606 ( .A(G134GAT), .B(KEYINPUT51), .Z(n543) );
  NAND2_X1 U607 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(G1343GAT) );
  NOR2_X1 U609 ( .A1(n563), .A2(n544), .ZN(n554) );
  NAND2_X1 U610 ( .A1(n554), .A2(n564), .ZN(n545) );
  XNOR2_X1 U611 ( .A(G141GAT), .B(n545), .ZN(G1344GAT) );
  NAND2_X1 U612 ( .A1(n554), .A2(n546), .ZN(n552) );
  XOR2_X1 U613 ( .A(KEYINPUT120), .B(KEYINPUT119), .Z(n548) );
  XNOR2_X1 U614 ( .A(KEYINPUT118), .B(KEYINPUT53), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n550) );
  XOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT52), .Z(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(G1345GAT) );
  NAND2_X1 U619 ( .A1(n554), .A2(n571), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U623 ( .A(G169GAT), .B(KEYINPUT123), .Z(n558) );
  NAND2_X1 U624 ( .A1(n559), .A2(n564), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(G1348GAT) );
  NAND2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n566) );
  NOR2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n574) );
  NAND2_X1 U630 ( .A1(n574), .A2(n564), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(n567), .ZN(G1352GAT) );
  XOR2_X1 U633 ( .A(G204GAT), .B(KEYINPUT61), .Z(n570) );
  NAND2_X1 U634 ( .A1(n574), .A2(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1353GAT) );
  NAND2_X1 U636 ( .A1(n574), .A2(n571), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n572), .B(KEYINPUT126), .ZN(n573) );
  XNOR2_X1 U638 ( .A(G211GAT), .B(n573), .ZN(G1354GAT) );
  INV_X1 U639 ( .A(n574), .ZN(n575) );
  NOR2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n578) );
  XNOR2_X1 U641 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(n579), .ZN(G1355GAT) );
endmodule

