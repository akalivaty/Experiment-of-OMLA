//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0 1 0 1 1 1 1 1 1 1 0 0 0 1 1 0 0 1 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 1 0 1 1 1 1 0 1 0 0 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n557,
    new_n558, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  NAND2_X1  g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI211_X1 g036(.A(G137), .B(new_n458), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  AOI21_X1  g040(.A(KEYINPUT68), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n462), .A2(KEYINPUT68), .A3(new_n465), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(new_n463), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(new_n459), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n469), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n467), .A2(new_n468), .B1(G2105), .B2(new_n475), .ZN(G160));
  NOR2_X1   g051(.A1(new_n473), .A2(new_n458), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n472), .A2(new_n458), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n458), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n478), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  INV_X1    g061(.A(G138), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n486), .B1(new_n479), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(KEYINPUT4), .A2(G138), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n489), .B1(new_n471), .B2(new_n459), .ZN(new_n490));
  AND2_X1   g065(.A1(G102), .A2(G2104), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n458), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G126), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n493), .B1(new_n471), .B2(new_n459), .ZN(new_n494));
  AND2_X1   g069(.A1(G114), .A2(G2104), .ZN(new_n495));
  OAI21_X1  g070(.A(G2105), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n488), .A2(new_n492), .A3(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  OAI21_X1  g074(.A(KEYINPUT70), .B1(new_n499), .B2(KEYINPUT5), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n501), .A2(new_n502), .A3(G543), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n504), .B1(new_n502), .B2(G543), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n499), .A2(KEYINPUT69), .A3(KEYINPUT5), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n500), .A2(new_n503), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n508));
  OR2_X1    g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n507), .A2(G62), .ZN(new_n515));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  XOR2_X1   g091(.A(new_n516), .B(KEYINPUT71), .Z(new_n517));
  AOI21_X1  g092(.A(new_n514), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n513), .A2(new_n518), .ZN(G166));
  INV_X1    g094(.A(G51), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n509), .A2(KEYINPUT72), .A3(new_n510), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n522));
  AND2_X1   g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n521), .A2(new_n525), .A3(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT73), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT73), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n521), .A2(new_n525), .A3(new_n528), .A4(G543), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n520), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n507), .A2(G89), .A3(new_n511), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n530), .A2(new_n535), .ZN(G168));
  NAND2_X1  g111(.A1(new_n500), .A2(new_n503), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n505), .A2(new_n506), .ZN(new_n538));
  AND3_X1   g113(.A1(new_n537), .A2(new_n538), .A3(new_n511), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G90), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n541), .B2(new_n514), .ZN(new_n542));
  INV_X1    g117(.A(G52), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n543), .B1(new_n527), .B2(new_n529), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n542), .A2(new_n544), .ZN(G171));
  NAND2_X1  g120(.A1(new_n527), .A2(new_n529), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G43), .ZN(new_n547));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n537), .A2(new_n538), .ZN(new_n549));
  INV_X1    g124(.A(G56), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n551), .A2(G651), .B1(G81), .B2(new_n539), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n547), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  INV_X1    g134(.A(G53), .ZN(new_n560));
  OR3_X1    g135(.A1(new_n526), .A2(KEYINPUT9), .A3(new_n560), .ZN(new_n561));
  OAI21_X1  g136(.A(KEYINPUT9), .B1(new_n526), .B2(new_n560), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n539), .A2(G91), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n549), .A2(KEYINPUT74), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT74), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n537), .A2(new_n538), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n568), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n563), .B(new_n564), .C1(new_n569), .C2(new_n514), .ZN(G299));
  INV_X1    g145(.A(G171), .ZN(G301));
  INV_X1    g146(.A(G168), .ZN(G286));
  INV_X1    g147(.A(G166), .ZN(G303));
  NAND2_X1  g148(.A1(new_n539), .A2(G87), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n499), .B1(new_n511), .B2(new_n522), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n575), .A2(G49), .A3(new_n521), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(G288));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n549), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G651), .ZN(new_n582));
  NAND2_X1  g157(.A1(G48), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G86), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n549), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(new_n511), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n582), .A2(new_n586), .ZN(G305));
  NAND2_X1  g162(.A1(new_n546), .A2(G47), .ZN(new_n588));
  NAND2_X1  g163(.A1(G72), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G60), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n549), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n591), .A2(G651), .B1(G85), .B2(new_n539), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n588), .A2(new_n592), .ZN(G290));
  AOI21_X1  g168(.A(new_n528), .B1(new_n575), .B2(new_n521), .ZN(new_n594));
  INV_X1    g169(.A(new_n529), .ZN(new_n595));
  OAI21_X1  g170(.A(G54), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n537), .A2(new_n538), .A3(G92), .A4(new_n511), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g174(.A1(new_n507), .A2(KEYINPUT10), .A3(G92), .A4(new_n511), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n596), .A2(new_n601), .ZN(new_n602));
  AND3_X1   g177(.A1(new_n537), .A2(new_n538), .A3(new_n566), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n566), .B1(new_n537), .B2(new_n538), .ZN(new_n604));
  OAI21_X1  g179(.A(G66), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(G79), .A2(G543), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n514), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT75), .ZN(new_n608));
  NOR3_X1   g183(.A1(new_n602), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(G66), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n610), .B1(new_n565), .B2(new_n567), .ZN(new_n611));
  INV_X1    g186(.A(new_n606), .ZN(new_n612));
  OAI21_X1  g187(.A(G651), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n546), .A2(G54), .B1(new_n599), .B2(new_n600), .ZN(new_n614));
  AOI21_X1  g189(.A(KEYINPUT75), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NOR3_X1   g190(.A1(new_n609), .A2(new_n615), .A3(G868), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(G868), .B2(G171), .ZN(G284));
  AOI21_X1  g192(.A(new_n616), .B1(G868), .B2(G171), .ZN(G321));
  NAND2_X1  g193(.A1(G286), .A2(G868), .ZN(new_n619));
  INV_X1    g194(.A(G299), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G868), .ZN(G297));
  XNOR2_X1  g196(.A(G297), .B(KEYINPUT76), .ZN(G280));
  NOR2_X1   g197(.A1(new_n609), .A2(new_n615), .ZN(new_n623));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(G860), .ZN(G148));
  NAND2_X1  g200(.A1(new_n613), .A2(new_n614), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(new_n608), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n613), .A2(new_n614), .A3(KEYINPUT75), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n627), .A2(new_n624), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G868), .ZN(new_n630));
  OAI22_X1  g205(.A1(new_n630), .A2(KEYINPUT77), .B1(G868), .B2(new_n554), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n631), .B1(KEYINPUT77), .B2(new_n630), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT78), .Z(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g209(.A1(new_n472), .A2(new_n464), .ZN(new_n635));
  XOR2_X1   g210(.A(KEYINPUT79), .B(KEYINPUT12), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  INV_X1    g213(.A(G2100), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n477), .A2(G123), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n480), .A2(G135), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n458), .A2(G111), .ZN(new_n643));
  OAI21_X1  g218(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n641), .B(new_n642), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(G2096), .Z(new_n646));
  NAND2_X1  g221(.A1(new_n638), .A2(new_n639), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n640), .A2(new_n646), .A3(new_n647), .ZN(G156));
  XNOR2_X1  g223(.A(G2427), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2430), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(KEYINPUT14), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G1341), .B(G1348), .Z(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n654), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2451), .B(G2454), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n659), .B(new_n660), .Z(new_n661));
  OR2_X1    g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n658), .A2(new_n661), .ZN(new_n663));
  AND3_X1   g238(.A1(new_n662), .A2(G14), .A3(new_n663), .ZN(G401));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  XNOR2_X1  g240(.A(G2072), .B(G2078), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT18), .Z(new_n669));
  AOI21_X1  g244(.A(new_n667), .B1(new_n666), .B2(KEYINPUT81), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n670), .B1(KEYINPUT81), .B2(new_n666), .ZN(new_n671));
  INV_X1    g246(.A(new_n665), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n666), .B(KEYINPUT17), .Z(new_n673));
  INV_X1    g248(.A(new_n667), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n671), .B(new_n672), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n673), .A2(new_n674), .A3(new_n665), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n669), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2096), .B(G2100), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G227));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT82), .ZN(new_n681));
  XOR2_X1   g256(.A(G1961), .B(G1966), .Z(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n683), .A2(KEYINPUT83), .ZN(new_n684));
  XOR2_X1   g259(.A(G1971), .B(G1976), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT19), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(KEYINPUT83), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n684), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT20), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n681), .A2(new_n682), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(new_n683), .B2(new_n686), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT84), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n686), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n691), .B(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n689), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(G1991), .B(G1996), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1981), .B(G1986), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(G229));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G33), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT25), .ZN(new_n706));
  AOI22_X1  g281(.A1(new_n472), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n707), .A2(new_n458), .ZN(new_n708));
  AOI211_X1 g283(.A(new_n706), .B(new_n708), .C1(G139), .C2(new_n480), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n704), .B1(new_n709), .B2(new_n703), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G2072), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT91), .Z(new_n712));
  NAND2_X1  g287(.A1(new_n703), .A2(G35), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G162), .B2(new_n703), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT97), .B(KEYINPUT29), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G2090), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n714), .B(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT30), .B(G28), .ZN(new_n718));
  OR2_X1    g293(.A1(KEYINPUT31), .A2(G11), .ZN(new_n719));
  NAND2_X1  g294(.A1(KEYINPUT31), .A2(G11), .ZN(new_n720));
  AOI22_X1  g295(.A1(new_n718), .A2(new_n703), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OAI221_X1 g296(.A(new_n721), .B1(new_n703), .B2(new_n645), .C1(new_n710), .C2(G2072), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT24), .B(G34), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(new_n703), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT90), .ZN(new_n725));
  INV_X1    g300(.A(G160), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(new_n703), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(G2084), .Z(new_n728));
  OR4_X1    g303(.A1(new_n712), .A2(new_n717), .A3(new_n722), .A4(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(G29), .A2(G32), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n477), .A2(G129), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n464), .A2(G105), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G141), .B2(new_n480), .ZN(new_n734));
  NAND3_X1  g309(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT92), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT26), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT93), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n730), .B1(new_n739), .B2(G29), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT27), .B(G1996), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G1966), .ZN(new_n743));
  INV_X1    g318(.A(G16), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G21), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G168), .B2(new_n744), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n740), .A2(new_n742), .B1(new_n743), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(G171), .A2(new_n744), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G5), .B2(new_n744), .ZN(new_n750));
  INV_X1    g325(.A(G1961), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n703), .A2(G27), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G164), .B2(new_n703), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT96), .ZN(new_n754));
  INV_X1    g329(.A(G2078), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n750), .A2(new_n751), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n748), .A2(new_n756), .ZN(new_n757));
  OAI22_X1  g332(.A1(new_n740), .A2(new_n742), .B1(new_n755), .B2(new_n754), .ZN(new_n758));
  NOR3_X1   g333(.A1(new_n729), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n746), .A2(G1966), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT94), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n750), .A2(new_n751), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT95), .ZN(new_n763));
  AND3_X1   g338(.A1(new_n759), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n744), .A2(G19), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n554), .B2(new_n744), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT87), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G1341), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n703), .A2(G26), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT28), .ZN(new_n770));
  AOI22_X1  g345(.A1(G128), .A2(new_n477), .B1(new_n480), .B2(G140), .ZN(new_n771));
  OAI21_X1  g346(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n772));
  INV_X1    g347(.A(G116), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(G2105), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT88), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n770), .B1(new_n776), .B2(new_n703), .ZN(new_n777));
  INV_X1    g352(.A(G2067), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n744), .A2(G4), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n623), .B2(new_n744), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(G1348), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n781), .A2(G1348), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n768), .A2(new_n779), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT89), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n744), .A2(G20), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT23), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n620), .B2(new_n744), .ZN(new_n790));
  INV_X1    g365(.A(G1956), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n764), .A2(new_n786), .A3(new_n787), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n744), .A2(G6), .ZN(new_n794));
  INV_X1    g369(.A(G305), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(new_n744), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT86), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT32), .B(G1981), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n744), .A2(G22), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G166), .B2(new_n744), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(G1971), .Z(new_n803));
  NAND2_X1  g378(.A1(new_n744), .A2(G23), .ZN(new_n804));
  INV_X1    g379(.A(G288), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n805), .B2(new_n744), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT33), .B(G1976), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n799), .A2(new_n800), .A3(new_n803), .A4(new_n808), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n809), .A2(KEYINPUT34), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(KEYINPUT34), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n744), .A2(G24), .ZN(new_n812));
  INV_X1    g387(.A(G290), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n812), .B1(new_n813), .B2(new_n744), .ZN(new_n814));
  INV_X1    g389(.A(G1986), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n477), .A2(G119), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n480), .A2(G131), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n458), .A2(G107), .ZN(new_n819));
  OAI21_X1  g394(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n817), .B(new_n818), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G29), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n703), .A2(G25), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT85), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT35), .B(G1991), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n810), .A2(new_n811), .A3(new_n816), .A4(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT36), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n793), .A2(new_n830), .ZN(G311));
  INV_X1    g406(.A(G311), .ZN(G150));
  INV_X1    g407(.A(G860), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n623), .A2(G559), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT38), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n539), .A2(G81), .ZN(new_n836));
  AOI22_X1  g411(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n836), .B1(new_n837), .B2(new_n514), .ZN(new_n838));
  INV_X1    g413(.A(G43), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(new_n527), .B2(new_n529), .ZN(new_n840));
  XNOR2_X1  g415(.A(KEYINPUT98), .B(G93), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n507), .A2(new_n511), .A3(new_n841), .ZN(new_n842));
  AOI22_X1  g417(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n842), .B1(new_n843), .B2(new_n514), .ZN(new_n844));
  INV_X1    g419(.A(G55), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(new_n527), .B2(new_n529), .ZN(new_n846));
  OAI22_X1  g421(.A1(new_n838), .A2(new_n840), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(G55), .B1(new_n594), .B2(new_n595), .ZN(new_n848));
  AND4_X1   g423(.A1(new_n538), .A2(new_n537), .A3(new_n511), .A4(new_n841), .ZN(new_n849));
  NAND2_X1  g424(.A1(G80), .A2(G543), .ZN(new_n850));
  INV_X1    g425(.A(G67), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n850), .B1(new_n549), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n849), .B1(new_n852), .B2(G651), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n547), .A2(new_n552), .A3(new_n848), .A4(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n847), .A2(new_n854), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n835), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n835), .A2(new_n855), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n833), .B1(new_n858), .B2(KEYINPUT39), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n856), .A2(new_n857), .A3(KEYINPUT39), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT99), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n860), .A2(new_n861), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n859), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(G860), .B1(new_n844), .B2(new_n846), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT37), .ZN(new_n867));
  OAI21_X1  g442(.A(KEYINPUT100), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT100), .ZN(new_n869));
  INV_X1    g444(.A(new_n867), .ZN(new_n870));
  INV_X1    g445(.A(new_n864), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n871), .A2(new_n862), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n869), .B(new_n870), .C1(new_n872), .C2(new_n859), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n868), .A2(new_n873), .ZN(G145));
  XNOR2_X1  g449(.A(new_n776), .B(new_n497), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n477), .A2(G130), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n458), .A2(G118), .ZN(new_n877));
  OAI21_X1  g452(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n480), .A2(KEYINPUT101), .A3(G142), .ZN(new_n879));
  AOI21_X1  g454(.A(KEYINPUT101), .B1(new_n480), .B2(G142), .ZN(new_n880));
  OAI221_X1 g455(.A(new_n876), .B1(new_n877), .B2(new_n878), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n875), .B(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n821), .B(new_n637), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n882), .B(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n739), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n709), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n886), .B1(new_n738), .B2(new_n709), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n884), .B(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(G162), .B(G160), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(new_n645), .ZN(new_n890));
  AOI21_X1  g465(.A(G37), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n891), .B1(new_n890), .B2(new_n888), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g468(.A1(new_n844), .A2(new_n846), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n894), .A2(G868), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT104), .ZN(new_n896));
  NAND2_X1  g471(.A1(G288), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n574), .A2(KEYINPUT104), .A3(new_n576), .A4(new_n577), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n897), .A2(G305), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(G305), .B1(new_n897), .B2(new_n898), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(G290), .A2(G166), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n813), .A2(G303), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n602), .A2(new_n607), .ZN(new_n908));
  NAND2_X1  g483(.A1(G299), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n564), .ZN(new_n910));
  OAI21_X1  g485(.A(G65), .B1(new_n603), .B2(new_n604), .ZN(new_n911));
  NAND2_X1  g486(.A1(G78), .A2(G543), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n910), .B1(new_n913), .B2(G651), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n626), .A2(new_n914), .A3(new_n563), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT103), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n909), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(G299), .A2(new_n908), .A3(KEYINPUT103), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(KEYINPUT41), .A3(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT41), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n909), .A2(new_n915), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n855), .A2(KEYINPUT102), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT102), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n847), .A2(new_n854), .A3(new_n923), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n623), .A2(new_n922), .A3(new_n624), .A4(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n923), .B1(new_n847), .B2(new_n854), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n847), .A2(new_n854), .A3(new_n923), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n629), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AOI22_X1  g503(.A1(new_n919), .A2(new_n921), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n917), .A2(new_n918), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n930), .A2(new_n925), .A3(new_n928), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n929), .A2(new_n931), .A3(KEYINPUT42), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT42), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n919), .A2(new_n921), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n925), .A2(new_n928), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n930), .A2(new_n925), .A3(new_n928), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n933), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n907), .B1(new_n932), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(KEYINPUT42), .B1(new_n929), .B2(new_n931), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n936), .A2(new_n933), .A3(new_n937), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(new_n941), .A3(new_n906), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n939), .A2(G868), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n895), .B1(new_n943), .B2(KEYINPUT105), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT105), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n939), .A2(new_n945), .A3(G868), .A4(new_n942), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n944), .A2(new_n946), .ZN(G295));
  INV_X1    g522(.A(KEYINPUT106), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n943), .A2(KEYINPUT105), .ZN(new_n949));
  INV_X1    g524(.A(new_n895), .ZN(new_n950));
  AND4_X1   g525(.A1(new_n948), .A2(new_n949), .A3(new_n946), .A4(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n948), .B1(new_n944), .B2(new_n946), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(G331));
  INV_X1    g528(.A(KEYINPUT111), .ZN(new_n954));
  NAND2_X1  g529(.A1(G77), .A2(G543), .ZN(new_n955));
  INV_X1    g530(.A(G64), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n955), .B1(new_n549), .B2(new_n956), .ZN(new_n957));
  AOI22_X1  g532(.A1(new_n957), .A2(G651), .B1(G90), .B2(new_n539), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n546), .A2(G51), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(new_n960));
  OAI21_X1  g535(.A(G52), .B1(new_n594), .B2(new_n595), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n958), .A2(new_n959), .A3(new_n960), .A4(new_n961), .ZN(new_n962));
  OAI22_X1  g537(.A1(new_n542), .A2(new_n544), .B1(new_n530), .B2(new_n535), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n965));
  OR3_X1    g540(.A1(new_n855), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n855), .A2(new_n964), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n847), .A2(new_n962), .A3(new_n854), .A4(new_n963), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n967), .A2(new_n965), .A3(new_n968), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n919), .A2(new_n921), .A3(new_n966), .A4(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT108), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n967), .A2(new_n971), .A3(new_n968), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n855), .A2(new_n964), .A3(KEYINPUT108), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n917), .A2(new_n918), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n970), .A2(new_n976), .A3(new_n906), .ZN(new_n977));
  INV_X1    g552(.A(G37), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n966), .A2(new_n969), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n975), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT109), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT109), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n980), .A2(new_n975), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n930), .A2(new_n920), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n909), .A2(new_n915), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT41), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n985), .A2(new_n973), .A3(new_n972), .A4(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n982), .A2(new_n984), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n979), .B1(new_n907), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT43), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n989), .A2(new_n907), .ZN(new_n993));
  INV_X1    g568(.A(new_n979), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n993), .A2(new_n994), .A3(new_n991), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n954), .B1(new_n992), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT43), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n993), .A2(new_n994), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n997), .B1(new_n998), .B2(KEYINPUT110), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n990), .A2(new_n991), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n999), .A2(KEYINPUT111), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT44), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n906), .B1(new_n970), .B2(new_n976), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n979), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1002), .B1(new_n1004), .B2(new_n997), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n996), .A2(new_n1001), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n990), .A2(new_n997), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(new_n997), .B2(new_n1004), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n1002), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1006), .A2(new_n1009), .ZN(G397));
  INV_X1    g585(.A(G1384), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT45), .B1(new_n497), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n475), .A2(G2105), .ZN(new_n1014));
  INV_X1    g589(.A(new_n468), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1014), .B(G40), .C1(new_n466), .C2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n776), .B(G2067), .ZN(new_n1018));
  INV_X1    g593(.A(new_n738), .ZN(new_n1019));
  INV_X1    g594(.A(G1996), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1018), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1021), .B1(new_n739), .B2(new_n1020), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n821), .B(new_n826), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1022), .B(new_n1023), .C1(new_n815), .C2(new_n813), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n813), .A2(new_n815), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n1025), .B(KEYINPUT112), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1017), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT119), .ZN(new_n1028));
  NAND2_X1  g603(.A1(G305), .A2(G1981), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT49), .ZN(new_n1030));
  INV_X1    g605(.A(G1981), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n582), .A2(new_n586), .A3(new_n1031), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n1029), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1030), .B1(new_n1029), .B2(new_n1032), .ZN(new_n1034));
  NAND4_X1  g609(.A1(G160), .A2(G40), .A3(new_n1011), .A4(new_n497), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT115), .B1(new_n1035), .B2(G8), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n497), .A2(new_n1011), .ZN(new_n1037));
  OAI211_X1 g612(.A(KEYINPUT115), .B(G8), .C1(new_n1016), .C2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  OAI22_X1  g614(.A1(new_n1033), .A2(new_n1034), .B1(new_n1036), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n805), .A2(G1976), .ZN(new_n1041));
  INV_X1    g616(.A(G1976), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT52), .B1(G288), .B2(new_n1042), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1041), .B(new_n1043), .C1(new_n1036), .C2(new_n1039), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1016), .A2(new_n1037), .ZN(new_n1046));
  INV_X1    g621(.A(G8), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1045), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n1048), .A2(new_n1038), .B1(G1976), .B2(new_n805), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1040), .B(new_n1044), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n1011), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT113), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n1013), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1016), .B1(new_n1012), .B2(KEYINPUT113), .ZN(new_n1056));
  AOI21_X1  g631(.A(G1971), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1037), .A2(KEYINPUT50), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1016), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n497), .A2(new_n1060), .A3(new_n1011), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1058), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1062), .A2(G2090), .ZN(new_n1063));
  OAI21_X1  g638(.A(G8), .B1(new_n1057), .B2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(G166), .A2(new_n1047), .ZN(new_n1065));
  AND2_X1   g640(.A1(KEYINPUT114), .A2(KEYINPUT55), .ZN(new_n1066));
  OR2_X1    g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(KEYINPUT114), .A2(KEYINPUT55), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1065), .B1(new_n1068), .B2(new_n1066), .ZN(new_n1069));
  AND2_X1   g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1064), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1051), .B1(new_n1052), .B2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1064), .A2(new_n1070), .A3(KEYINPUT116), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1074), .B(G8), .C1(new_n1057), .C2(new_n1063), .ZN(new_n1075));
  AND2_X1   g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1013), .A2(new_n1059), .A3(new_n1053), .ZN(new_n1077));
  XNOR2_X1  g652(.A(KEYINPUT117), .B(G2084), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  OAI22_X1  g654(.A1(new_n1077), .A2(G1966), .B1(new_n1062), .B2(new_n1079), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1080), .A2(G8), .A3(G168), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1072), .A2(new_n1076), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT63), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT118), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1064), .A2(new_n1070), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1084), .B1(new_n1085), .B2(new_n1051), .ZN(new_n1086));
  AND2_X1   g661(.A1(new_n1040), .A2(new_n1044), .ZN(new_n1087));
  OR2_X1    g662(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1087), .A2(new_n1071), .A3(new_n1088), .A4(KEYINPUT118), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1081), .A2(new_n1075), .A3(KEYINPUT63), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1082), .A2(new_n1083), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1051), .A2(new_n1075), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1048), .A2(new_n1038), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1040), .A2(new_n1042), .A3(new_n805), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n1032), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1093), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1028), .B1(new_n1092), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1102), .A2(KEYINPUT119), .A3(new_n1097), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1099), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1105), .B1(new_n1106), .B2(G2078), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1105), .A2(G2078), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1077), .A2(new_n1108), .B1(new_n1062), .B2(new_n751), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(G171), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1080), .B(G168), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT51), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1113), .A2(new_n1047), .ZN(new_n1114));
  OAI21_X1  g689(.A(G8), .B1(new_n1080), .B2(G286), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1112), .A2(new_n1114), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1111), .B1(new_n1116), .B2(KEYINPUT62), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1072), .A2(new_n1076), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1117), .B(new_n1118), .C1(KEYINPUT62), .C2(new_n1116), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT56), .B(G2072), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1055), .A2(new_n1120), .A3(new_n1056), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT122), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1055), .A2(new_n1056), .A3(KEYINPUT122), .A4(new_n1120), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1062), .A2(new_n791), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  OR2_X1    g702(.A1(new_n914), .A2(KEYINPUT120), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n914), .A2(KEYINPUT120), .B1(new_n562), .B2(new_n561), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT57), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n620), .A2(KEYINPUT57), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1127), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT123), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1046), .A2(new_n778), .ZN(new_n1138));
  INV_X1    g713(.A(G1348), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1137), .A2(new_n1138), .B1(new_n1062), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1046), .A2(KEYINPUT123), .A3(new_n778), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n626), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1136), .A2(new_n1142), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1144));
  OAI21_X1  g719(.A(KEYINPUT121), .B1(new_n1144), .B2(KEYINPUT57), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1145), .A2(new_n1132), .A3(new_n1134), .A4(new_n1126), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(KEYINPUT61), .B1(new_n1136), .B2(new_n1146), .ZN(new_n1148));
  XNOR2_X1  g723(.A(KEYINPUT58), .B(G1341), .ZN(new_n1149));
  OAI22_X1  g724(.A1(new_n1106), .A2(G1996), .B1(new_n1046), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n554), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT59), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n626), .A2(KEYINPUT60), .ZN(new_n1154));
  AOI22_X1  g729(.A1(new_n1151), .A2(new_n1152), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n1140), .A2(new_n626), .A3(new_n1141), .ZN(new_n1156));
  OAI21_X1  g731(.A(KEYINPUT60), .B1(new_n1156), .B2(new_n1142), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1150), .A2(KEYINPUT59), .A3(new_n554), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1155), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1148), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1136), .A2(new_n1146), .A3(KEYINPUT61), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1147), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1110), .B(G171), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT54), .ZN(new_n1164));
  OR2_X1    g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1165), .A2(new_n1118), .A3(new_n1166), .A4(new_n1116), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1119), .B1(new_n1162), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1027), .B1(new_n1104), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT46), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n1172), .B(KEYINPUT124), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1174));
  AOI22_X1  g749(.A1(new_n1174), .A2(new_n1017), .B1(new_n1171), .B2(new_n1170), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  XOR2_X1   g751(.A(new_n1176), .B(KEYINPUT125), .Z(new_n1177));
  OR2_X1    g752(.A1(new_n1177), .A2(KEYINPUT47), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(KEYINPUT47), .ZN(new_n1179));
  AOI21_X1  g754(.A(KEYINPUT48), .B1(new_n1026), .B2(new_n1017), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1180), .B1(new_n1181), .B2(new_n1017), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1026), .A2(KEYINPUT48), .A3(new_n1017), .ZN(new_n1183));
  INV_X1    g758(.A(new_n826), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n821), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1022), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n776), .A2(new_n778), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  AOI22_X1  g763(.A1(new_n1182), .A2(new_n1183), .B1(new_n1188), .B2(new_n1017), .ZN(new_n1189));
  AND3_X1   g764(.A1(new_n1178), .A2(new_n1179), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1169), .A2(new_n1190), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g766(.A(G319), .ZN(new_n1193));
  NOR2_X1   g767(.A1(G227), .A2(new_n1193), .ZN(new_n1194));
  XOR2_X1   g768(.A(new_n1194), .B(KEYINPUT126), .Z(new_n1195));
  NOR2_X1   g769(.A1(new_n1195), .A2(G401), .ZN(new_n1196));
  XNOR2_X1  g770(.A(new_n1196), .B(KEYINPUT127), .ZN(new_n1197));
  NAND4_X1  g771(.A1(new_n892), .A2(new_n1008), .A3(new_n701), .A4(new_n1197), .ZN(G225));
  INV_X1    g772(.A(G225), .ZN(G308));
endmodule


