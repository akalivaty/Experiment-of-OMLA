//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 1 0 1 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n202), .A2(new_n203), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n210), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(KEYINPUT64), .B(G77), .ZN(new_n218));
  AND2_X1   g0018(.A1(new_n218), .A2(G244), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G58), .A2(G232), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n207), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n217), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT65), .Z(G361));
  XOR2_X1   g0029(.A(G250), .B(G257), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT66), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n233), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT67), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  XNOR2_X1  g0047(.A(KEYINPUT3), .B(G33), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n248), .A2(G223), .A3(G1698), .ZN(new_n249));
  INV_X1    g0049(.A(new_n218), .ZN(new_n250));
  INV_X1    g0050(.A(G222), .ZN(new_n251));
  INV_X1    g0051(.A(G1698), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  OAI221_X1 g0053(.A(new_n249), .B1(new_n250), .B2(new_n248), .C1(new_n251), .C2(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n211), .B1(G33), .B2(G41), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G274), .ZN(new_n257));
  AND2_X1   g0057(.A1(G1), .A2(G13), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT68), .B(G45), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n260), .B(new_n261), .C1(new_n262), .C2(G41), .ZN(new_n263));
  OR2_X1    g0063(.A1(KEYINPUT69), .A2(G1), .ZN(new_n264));
  NAND2_X1  g0064(.A1(KEYINPUT69), .A2(G1), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n264), .A2(G41), .A3(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n264), .A2(G45), .A3(new_n265), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n258), .A2(new_n259), .ZN(new_n268));
  AND3_X1   g0068(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G226), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n256), .A2(new_n263), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT70), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n256), .A2(KEYINPUT70), .A3(new_n263), .A4(new_n270), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(G190), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n264), .A2(G13), .A3(G20), .A4(new_n265), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n201), .ZN(new_n280));
  AND2_X1   g0080(.A1(KEYINPUT69), .A2(G1), .ZN(new_n281));
  NOR2_X1   g0081(.A1(KEYINPUT69), .A2(G1), .ZN(new_n282));
  NOR3_X1   g0082(.A1(new_n281), .A2(new_n282), .A3(new_n212), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n211), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n280), .B1(new_n287), .B2(new_n201), .ZN(new_n288));
  INV_X1    g0088(.A(new_n285), .ZN(new_n289));
  NAND2_X1  g0089(.A1(KEYINPUT71), .A2(G58), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n290), .B(KEYINPUT8), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(new_n212), .A3(G33), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G20), .A2(G33), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n289), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n288), .A2(new_n295), .ZN(new_n296));
  OR2_X1    g0096(.A1(new_n296), .A2(KEYINPUT9), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(KEYINPUT9), .ZN(new_n298));
  NAND2_X1  g0098(.A1(KEYINPUT74), .A2(KEYINPUT10), .ZN(new_n299));
  AND3_X1   g0099(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n273), .A2(G200), .A3(new_n275), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n277), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(KEYINPUT74), .A2(KEYINPUT10), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G169), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n273), .A2(new_n305), .A3(new_n275), .ZN(new_n306));
  INV_X1    g0106(.A(new_n296), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g0108(.A(KEYINPUT72), .B(G179), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n274), .A2(new_n276), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n308), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n303), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n277), .A2(new_n300), .A3(new_n313), .A4(new_n301), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n304), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT78), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT18), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n287), .A2(new_n291), .ZN(new_n318));
  INV_X1    g0118(.A(new_n291), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n278), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT7), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(new_n248), .B2(G20), .ZN(new_n324));
  INV_X1    g0124(.A(G33), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT3), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT3), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G33), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n329), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n203), .B1(new_n324), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(KEYINPUT77), .B1(new_n202), .B2(new_n203), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT77), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n333), .A2(G58), .A3(G68), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(new_n214), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G20), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n293), .A2(G159), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n331), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n289), .B1(new_n339), .B2(KEYINPUT16), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT16), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(new_n331), .B2(new_n338), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n322), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n326), .A2(new_n328), .A3(G223), .A4(new_n252), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n326), .A2(new_n328), .A3(G226), .A4(G1698), .ZN(new_n345));
  INV_X1    g0145(.A(G87), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n344), .B(new_n345), .C1(new_n325), .C2(new_n346), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n347), .A2(new_n255), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n266), .A2(new_n267), .A3(G232), .A4(new_n268), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n263), .ZN(new_n350));
  OAI21_X1  g0150(.A(G169), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n347), .A2(new_n255), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n352), .A2(new_n310), .A3(new_n263), .A4(new_n349), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n316), .B(new_n317), .C1(new_n343), .C2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n324), .A2(new_n330), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(G68), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n335), .A2(G20), .B1(G159), .B2(new_n293), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n358), .A2(KEYINPUT16), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n360), .A2(new_n342), .A3(new_n285), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n352), .A2(G190), .A3(new_n263), .A4(new_n349), .ZN(new_n362));
  OAI21_X1  g0162(.A(G200), .B1(new_n348), .B2(new_n350), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n361), .A2(new_n321), .A3(new_n362), .A4(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT17), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n343), .A2(KEYINPUT17), .A3(new_n362), .A4(new_n363), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n356), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(KEYINPUT18), .B1(new_n343), .B2(new_n355), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n361), .A2(new_n321), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n370), .A2(new_n317), .A3(new_n354), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n316), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  OR2_X1    g0172(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT75), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n212), .A2(G33), .A3(G77), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n203), .A2(G20), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n212), .A2(new_n325), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n375), .B(new_n376), .C1(new_n377), .C2(new_n201), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n378), .A2(KEYINPUT11), .A3(new_n285), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(KEYINPUT11), .B1(new_n378), .B2(new_n285), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n374), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n381), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n383), .A2(KEYINPUT75), .A3(new_n379), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT12), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n279), .A2(new_n385), .A3(new_n203), .ZN(new_n386));
  OAI21_X1  g0186(.A(KEYINPUT12), .B1(new_n278), .B2(G68), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n386), .A2(new_n387), .B1(new_n286), .B2(G68), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n382), .A2(new_n384), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT76), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n382), .A2(new_n384), .A3(new_n388), .A4(KEYINPUT76), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n266), .A2(new_n267), .A3(G238), .A4(new_n268), .ZN(new_n395));
  NOR2_X1   g0195(.A1(G226), .A2(G1698), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n396), .B1(new_n235), .B2(G1698), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n397), .A2(new_n248), .B1(G33), .B2(G97), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n263), .B(new_n395), .C1(new_n398), .C2(new_n268), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT13), .ZN(new_n400));
  NAND2_X1  g0200(.A1(G33), .A2(G97), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n235), .A2(G1698), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(G226), .B2(G1698), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n401), .B1(new_n403), .B2(new_n329), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n255), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT13), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n405), .A2(new_n406), .A3(new_n263), .A4(new_n395), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n305), .B1(new_n400), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT14), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n400), .A2(G179), .A3(new_n407), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n408), .A2(new_n409), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n394), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n400), .A2(new_n407), .ZN(new_n415));
  INV_X1    g0215(.A(G190), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n417), .B1(G200), .B2(new_n415), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n393), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n248), .A2(G238), .A3(G1698), .ZN(new_n420));
  INV_X1    g0220(.A(G107), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n420), .B1(new_n421), .B2(new_n248), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT73), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(new_n253), .B2(new_n235), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n248), .A2(KEYINPUT73), .A3(G232), .A4(new_n252), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n422), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n426), .A2(new_n268), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n269), .A2(G244), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n263), .ZN(new_n429));
  OAI21_X1  g0229(.A(G200), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n429), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n431), .B(G190), .C1(new_n268), .C2(new_n426), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n218), .A2(G20), .ZN(new_n433));
  XNOR2_X1  g0233(.A(KEYINPUT8), .B(G58), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n212), .A2(G33), .ZN(new_n435));
  XNOR2_X1  g0235(.A(KEYINPUT15), .B(G87), .ZN(new_n436));
  OAI221_X1 g0236(.A(new_n433), .B1(new_n377), .B2(new_n434), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n437), .A2(new_n285), .ZN(new_n438));
  INV_X1    g0238(.A(G77), .ZN(new_n439));
  OAI22_X1  g0239(.A1(new_n287), .A2(new_n439), .B1(new_n218), .B2(new_n278), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n430), .A2(new_n432), .A3(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n305), .B1(new_n427), .B2(new_n429), .ZN(new_n443));
  INV_X1    g0243(.A(new_n441), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n431), .B(new_n309), .C1(new_n268), .C2(new_n426), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n414), .A2(new_n419), .A3(new_n442), .A4(new_n446), .ZN(new_n447));
  NOR3_X1   g0247(.A1(new_n315), .A2(new_n373), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(KEYINPUT88), .A2(KEYINPUT25), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n421), .B1(KEYINPUT88), .B2(KEYINPUT25), .ZN(new_n450));
  OR3_X1    g0250(.A1(new_n278), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n449), .B1(new_n278), .B2(new_n450), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n264), .A2(G33), .A3(new_n265), .ZN(new_n453));
  AND3_X1   g0253(.A1(new_n278), .A2(new_n289), .A3(new_n453), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n451), .A2(new_n452), .B1(new_n454), .B2(G107), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G33), .A2(G116), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(G20), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT87), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n458), .B1(new_n212), .B2(G107), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT23), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT23), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n458), .B(new_n461), .C1(new_n212), .C2(G107), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n457), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g0263(.A1(KEYINPUT86), .A2(KEYINPUT22), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n248), .A2(new_n212), .A3(G87), .A4(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n326), .A2(new_n328), .A3(new_n212), .A4(G87), .ZN(new_n466));
  NOR2_X1   g0266(.A1(KEYINPUT86), .A2(KEYINPUT22), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n463), .A2(new_n465), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT24), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT24), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n463), .A2(new_n472), .A3(new_n469), .A4(new_n465), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n455), .B1(new_n474), .B2(new_n289), .ZN(new_n475));
  INV_X1    g0275(.A(G45), .ZN(new_n476));
  NOR3_X1   g0276(.A1(new_n281), .A2(new_n282), .A3(new_n476), .ZN(new_n477));
  XNOR2_X1  g0277(.A(KEYINPUT5), .B(G41), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n255), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(G264), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n326), .A2(new_n328), .A3(G250), .A4(new_n252), .ZN(new_n481));
  NAND2_X1  g0281(.A1(G33), .A2(G294), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n326), .A2(new_n328), .A3(G257), .A4(G1698), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT89), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n248), .A2(KEYINPUT89), .A3(G257), .A4(G1698), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n483), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n480), .B1(new_n488), .B2(new_n268), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n281), .A2(new_n282), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n260), .A2(new_n490), .A3(new_n478), .A4(G45), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT81), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n477), .A2(KEYINPUT81), .A3(new_n260), .A4(new_n478), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n489), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(G179), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n305), .B1(new_n489), .B2(new_n496), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n475), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n289), .B1(new_n471), .B2(new_n473), .ZN(new_n502));
  INV_X1    g0302(.A(new_n455), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n489), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(G190), .A3(new_n495), .ZN(new_n506));
  OAI21_X1  g0306(.A(G200), .B1(new_n489), .B2(new_n496), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n504), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n493), .A2(new_n494), .B1(G257), .B2(new_n479), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n326), .A2(new_n328), .A3(G250), .A4(G1698), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G283), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n326), .A2(new_n328), .A3(G244), .A4(new_n252), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT4), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n510), .B(new_n511), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n512), .A2(new_n513), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n255), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n509), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n305), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n509), .A2(new_n309), .A3(new_n516), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n357), .A2(G107), .ZN(new_n520));
  NOR4_X1   g0320(.A1(new_n439), .A2(KEYINPUT79), .A3(G20), .A4(G33), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT79), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n522), .B1(new_n293), .B2(G77), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n421), .A2(KEYINPUT6), .A3(G97), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT6), .ZN(new_n527));
  XNOR2_X1  g0327(.A(G97), .B(G107), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(KEYINPUT80), .B(new_n524), .C1(new_n529), .C2(new_n212), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT80), .ZN(new_n531));
  AND2_X1   g0331(.A1(G97), .A2(G107), .ZN(new_n532));
  NOR2_X1   g0332(.A1(G97), .A2(G107), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n527), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n212), .B1(new_n534), .B2(new_n525), .ZN(new_n535));
  OAI21_X1  g0335(.A(KEYINPUT79), .B1(new_n377), .B2(new_n439), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n293), .A2(new_n522), .A3(G77), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n531), .B1(new_n535), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n520), .A2(new_n530), .A3(new_n539), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n540), .A2(new_n285), .ZN(new_n541));
  INV_X1    g0341(.A(G97), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n279), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n278), .A2(new_n289), .A3(new_n453), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n543), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n518), .B(new_n519), .C1(new_n541), .C2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n517), .A2(G200), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n545), .B1(new_n540), .B2(new_n285), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n547), .B(new_n548), .C1(new_n416), .C2(new_n517), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n501), .A2(new_n508), .A3(new_n546), .A4(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n248), .A2(G244), .A3(G1698), .ZN(new_n551));
  INV_X1    g0351(.A(G238), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n551), .B(new_n456), .C1(new_n253), .C2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n255), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n477), .A2(new_n255), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n555), .A2(G250), .B1(new_n260), .B2(new_n477), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n554), .A2(new_n556), .A3(new_n309), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(KEYINPUT82), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT82), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n554), .A2(new_n556), .A3(new_n559), .A4(new_n309), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  XOR2_X1   g0361(.A(KEYINPUT15), .B(G87), .Z(new_n562));
  NOR2_X1   g0362(.A1(new_n278), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT19), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n212), .B1(new_n401), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n533), .A2(new_n346), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n326), .A2(new_n328), .A3(new_n212), .A4(G68), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n564), .B1(new_n435), .B2(new_n542), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT83), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n289), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n567), .A2(new_n568), .A3(KEYINPUT83), .A4(new_n569), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n563), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n278), .A2(new_n562), .A3(new_n289), .A4(new_n453), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT84), .ZN(new_n576));
  XNOR2_X1  g0376(.A(new_n575), .B(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n554), .A2(new_n556), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n574), .A2(new_n577), .B1(new_n578), .B2(new_n305), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n561), .A2(new_n579), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n554), .A2(new_n556), .A3(G190), .ZN(new_n581));
  INV_X1    g0381(.A(G200), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n582), .B1(new_n554), .B2(new_n556), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n454), .A2(G87), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n574), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n580), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT21), .ZN(new_n589));
  INV_X1    g0389(.A(G116), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n284), .A2(new_n211), .B1(G20), .B2(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n511), .B(new_n212), .C1(G33), .C2(new_n542), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(KEYINPUT20), .A3(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT20), .B1(new_n591), .B2(new_n592), .ZN(new_n595));
  OAI22_X1  g0395(.A1(new_n594), .A2(new_n595), .B1(G116), .B2(new_n278), .ZN(new_n596));
  NOR3_X1   g0396(.A1(new_n544), .A2(KEYINPUT85), .A3(new_n590), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(KEYINPUT85), .B1(new_n544), .B2(new_n590), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n596), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(G303), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n268), .B1(new_n329), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(G257), .A2(G1698), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n252), .A2(G264), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n248), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n479), .A2(G270), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n495), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(G169), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n589), .B1(new_n600), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(G200), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n610), .B(new_n600), .C1(new_n416), .C2(new_n607), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n495), .A2(new_n606), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n278), .A2(G116), .ZN(new_n613));
  INV_X1    g0413(.A(new_n595), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n613), .B1(new_n614), .B2(new_n593), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT85), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(new_n454), .B2(G116), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n615), .B1(new_n617), .B2(new_n597), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n612), .A2(new_n618), .A3(G179), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n618), .A2(KEYINPUT21), .A3(G169), .A4(new_n607), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n609), .A2(new_n611), .A3(new_n619), .A4(new_n620), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n550), .A2(new_n588), .A3(new_n621), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n448), .A2(new_n622), .ZN(G372));
  INV_X1    g0423(.A(new_n312), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n304), .A2(new_n314), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n367), .A2(new_n366), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n414), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n446), .B1(new_n418), .B2(new_n393), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT93), .ZN(new_n631));
  AOI221_X4 g0431(.A(KEYINPUT18), .B1(new_n351), .B2(new_n353), .C1(new_n361), .C2(new_n321), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n317), .B1(new_n370), .B2(new_n354), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n369), .A2(KEYINPUT93), .A3(new_n371), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n625), .B1(new_n637), .B2(KEYINPUT94), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT94), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n630), .A2(new_n639), .A3(new_n636), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n624), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n448), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n620), .A2(new_n619), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n501), .A2(new_n643), .A3(new_n609), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n546), .A2(new_n549), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n574), .A2(new_n577), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n578), .A2(new_n305), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n646), .A2(new_n647), .A3(new_n557), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n574), .A2(new_n585), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(KEYINPUT90), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT90), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n574), .A2(new_n651), .A3(new_n585), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n648), .B1(new_n653), .B2(new_n584), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n644), .A2(new_n645), .A3(new_n654), .A4(new_n508), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n648), .B(KEYINPUT91), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n572), .A2(new_n573), .ZN(new_n658));
  INV_X1    g0458(.A(new_n563), .ZN(new_n659));
  AND4_X1   g0459(.A1(new_n651), .A2(new_n658), .A3(new_n585), .A4(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n651), .B1(new_n574), .B2(new_n585), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n584), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n479), .A2(G257), .ZN(new_n663));
  AND4_X1   g0463(.A1(new_n309), .A2(new_n516), .A3(new_n495), .A4(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(G169), .B1(new_n509), .B2(new_n516), .ZN(new_n665));
  NOR3_X1   g0465(.A1(new_n548), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n646), .A2(new_n647), .A3(new_n557), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n662), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT26), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(KEYINPUT92), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT92), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n668), .A2(new_n672), .A3(new_n669), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n561), .A2(new_n579), .B1(new_n584), .B2(new_n586), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n674), .A2(KEYINPUT26), .A3(new_n666), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n671), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n657), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n641), .B1(new_n642), .B2(new_n678), .ZN(G369));
  NAND2_X1  g0479(.A1(new_n643), .A2(new_n609), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n212), .A2(G13), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n490), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(G213), .B1(new_n682), .B2(KEYINPUT27), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(KEYINPUT95), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT95), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n682), .A2(new_n686), .A3(KEYINPUT27), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n683), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n688), .A2(G343), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(new_n600), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n680), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n621), .B2(new_n691), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(G330), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n508), .B1(new_n504), .B2(new_n690), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n698), .A2(new_n501), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n501), .A2(new_n689), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n697), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n680), .A2(new_n690), .ZN(new_n705));
  OAI22_X1  g0505(.A1(new_n699), .A2(new_n705), .B1(new_n501), .B2(new_n689), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n704), .A2(new_n707), .ZN(G399));
  INV_X1    g0508(.A(new_n208), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G41), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n566), .A2(G116), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(G1), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n215), .B2(new_n711), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT28), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT29), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n668), .A2(KEYINPUT26), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n674), .A2(new_n669), .A3(new_n666), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n655), .A2(new_n656), .A3(new_n717), .A4(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n716), .B1(new_n719), .B2(new_n690), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n689), .B1(new_n657), .B2(new_n676), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n720), .B1(new_n716), .B2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT31), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n612), .A2(G179), .A3(new_n516), .A4(new_n509), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n505), .A2(KEYINPUT96), .A3(new_n554), .A4(new_n556), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT96), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(new_n578), .B2(new_n489), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n724), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n578), .A2(KEYINPUT97), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n310), .B1(new_n495), .B2(new_n606), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT97), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n554), .A2(new_n556), .A3(new_n731), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n729), .A2(new_n517), .A3(new_n730), .A4(new_n732), .ZN(new_n733));
  OAI22_X1  g0533(.A1(new_n728), .A2(KEYINPUT30), .B1(new_n497), .B2(new_n733), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n517), .A2(new_n607), .A3(new_n498), .ZN(new_n735));
  INV_X1    g0535(.A(new_n727), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n578), .A2(new_n489), .A3(new_n726), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT30), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n689), .B1(new_n734), .B2(new_n740), .ZN(new_n741));
  AOI22_X1  g0541(.A1(new_n723), .A2(new_n741), .B1(new_n622), .B2(new_n690), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n733), .A2(new_n497), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n743), .B1(new_n738), .B2(new_n739), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n728), .A2(KEYINPUT30), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n690), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(KEYINPUT31), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n695), .B1(new_n742), .B2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n722), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n715), .B1(new_n751), .B2(G1), .ZN(G364));
  AOI21_X1  g0552(.A(new_n261), .B1(new_n681), .B2(G45), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n710), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n696), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n756), .B1(G330), .B2(new_n693), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n755), .B(KEYINPUT98), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n248), .A2(new_n208), .ZN(new_n759));
  INV_X1    g0559(.A(G355), .ZN(new_n760));
  OAI22_X1  g0560(.A1(new_n759), .A2(new_n760), .B1(G116), .B2(new_n208), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n246), .A2(G45), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n709), .A2(new_n248), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n215), .A2(new_n262), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n761), .B1(new_n762), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G13), .A2(G33), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G20), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n211), .B1(G20), .B2(new_n305), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n758), .B1(new_n767), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n309), .A2(new_n212), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n416), .A2(G200), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G322), .ZN(new_n779));
  INV_X1    g0579(.A(G311), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G190), .A2(G200), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n775), .A2(new_n781), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n778), .A2(new_n779), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n781), .A2(G20), .A3(new_n498), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n248), .B1(new_n785), .B2(G329), .ZN(new_n786));
  INV_X1    g0586(.A(G283), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n212), .A2(new_n582), .A3(G179), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(new_n416), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n786), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n776), .A2(new_n498), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G20), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G294), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n788), .A2(G190), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n793), .A2(new_n794), .B1(new_n601), .B2(new_n795), .ZN(new_n796));
  NOR3_X1   g0596(.A1(new_n783), .A2(new_n790), .A3(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(G326), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n775), .A2(G190), .A3(G200), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT101), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n775), .A2(new_n416), .A3(G200), .ZN(new_n801));
  XOR2_X1   g0601(.A(KEYINPUT33), .B(G317), .Z(new_n802));
  OAI221_X1 g0602(.A(new_n797), .B1(new_n798), .B2(new_n800), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n803), .A2(KEYINPUT102), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n792), .A2(G97), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(new_n801), .B2(new_n203), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT100), .Z(new_n807));
  OAI221_X1 g0607(.A(new_n248), .B1(new_n346), .B2(new_n795), .C1(new_n782), .C2(new_n250), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(G58), .B2(new_n777), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n789), .A2(new_n421), .ZN(new_n810));
  INV_X1    g0610(.A(G159), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n784), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g0612(.A(KEYINPUT99), .B(KEYINPUT32), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n812), .B(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n799), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n810), .B(new_n814), .C1(G50), .C2(new_n815), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n807), .A2(new_n809), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n803), .A2(KEYINPUT102), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n804), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n774), .B1(new_n819), .B2(new_n771), .ZN(new_n820));
  INV_X1    g0620(.A(new_n770), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n820), .B1(new_n693), .B2(new_n821), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n757), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(G396));
  NOR2_X1   g0624(.A1(new_n446), .A2(new_n689), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT105), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n690), .B2(new_n441), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n444), .A2(KEYINPUT105), .A3(new_n689), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n827), .A2(new_n442), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n825), .B1(new_n829), .B2(new_n446), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n690), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  AND3_X1   g0632(.A1(new_n668), .A2(new_n672), .A3(new_n669), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n672), .B1(new_n668), .B2(new_n669), .ZN(new_n834));
  NOR3_X1   g0634(.A1(new_n588), .A2(new_n669), .A3(new_n546), .ZN(new_n835));
  NOR3_X1   g0635(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n655), .A2(new_n656), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n832), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n721), .B2(new_n830), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n755), .B1(new_n839), .B2(new_n749), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n749), .B2(new_n839), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n789), .A2(new_n346), .ZN(new_n842));
  INV_X1    g0642(.A(new_n795), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n842), .B1(G107), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n248), .B1(new_n785), .B2(G311), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n844), .A2(new_n805), .A3(new_n845), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n801), .A2(new_n787), .B1(new_n782), .B2(new_n590), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT103), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n847), .A2(new_n848), .B1(new_n601), .B2(new_n799), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(new_n848), .B2(new_n847), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(KEYINPUT104), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n846), .B(new_n851), .C1(G294), .C2(new_n777), .ZN(new_n852));
  INV_X1    g0652(.A(new_n782), .ZN(new_n853));
  AOI22_X1  g0653(.A1(G159), .A2(new_n853), .B1(new_n777), .B2(G143), .ZN(new_n854));
  INV_X1    g0654(.A(G137), .ZN(new_n855));
  INV_X1    g0655(.A(G150), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n854), .B1(new_n855), .B2(new_n799), .C1(new_n856), .C2(new_n801), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT34), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n857), .A2(new_n858), .ZN(new_n860));
  INV_X1    g0660(.A(G132), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n248), .B1(new_n784), .B2(new_n861), .C1(new_n793), .C2(new_n202), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n201), .A2(new_n795), .B1(new_n789), .B2(new_n203), .ZN(new_n863));
  NOR4_X1   g0663(.A1(new_n859), .A2(new_n860), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n771), .B1(new_n852), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n758), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n771), .A2(new_n768), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n866), .B1(new_n439), .B2(new_n867), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n865), .B(new_n868), .C1(new_n769), .C2(new_n830), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n841), .A2(new_n869), .ZN(G384));
  INV_X1    g0670(.A(new_n529), .ZN(new_n871));
  OR2_X1    g0671(.A1(new_n871), .A2(KEYINPUT35), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(KEYINPUT35), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n872), .A2(G116), .A3(new_n213), .A4(new_n873), .ZN(new_n874));
  XOR2_X1   g0674(.A(new_n874), .B(KEYINPUT36), .Z(new_n875));
  OR3_X1    g0675(.A1(new_n335), .A2(new_n250), .A3(new_n201), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n201), .A2(G68), .ZN(new_n877));
  AOI211_X1 g0677(.A(G13), .B(new_n490), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n339), .A2(KEYINPUT107), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT107), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n331), .B2(new_n338), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n880), .A2(new_n341), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n322), .B1(new_n883), .B2(new_n340), .ZN(new_n884));
  INV_X1    g0684(.A(new_n688), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n368), .B2(new_n372), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n351), .A2(new_n885), .A3(new_n353), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n364), .B1(new_n884), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n370), .A2(new_n888), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n364), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n891), .B1(KEYINPUT37), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT38), .B1(new_n887), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n887), .A2(new_n894), .A3(KEYINPUT38), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n391), .A2(new_n689), .A3(new_n392), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n414), .A2(new_n419), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n899), .B1(new_n412), .B2(new_n413), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT106), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT106), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n899), .B(new_n904), .C1(new_n412), .C2(new_n413), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n901), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n830), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n742), .B2(new_n747), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT40), .B1(new_n898), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT37), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT108), .B1(new_n370), .B2(new_n888), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n893), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n892), .A2(KEYINPUT108), .A3(new_n364), .A4(KEYINPUT37), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n632), .A2(new_n633), .A3(new_n631), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT93), .B1(new_n369), .B2(new_n371), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n627), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n370), .A2(new_n688), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n914), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n897), .B1(new_n920), .B2(KEYINPUT38), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n908), .A2(new_n921), .A3(KEYINPUT40), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT109), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT40), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT38), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n918), .B1(new_n636), .B2(new_n627), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n926), .B1(new_n927), .B2(new_n914), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n925), .B1(new_n928), .B2(new_n897), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n929), .A2(KEYINPUT109), .A3(new_n908), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n909), .B1(new_n924), .B2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n741), .A2(new_n723), .ZN(new_n933));
  INV_X1    g0733(.A(new_n550), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n621), .A2(new_n588), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n934), .A2(new_n935), .A3(new_n690), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n747), .A2(new_n933), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n448), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(G330), .B1(new_n932), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n938), .B2(new_n932), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT39), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n921), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n628), .A2(new_n690), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n942), .B(new_n944), .C1(new_n941), .C2(new_n898), .ZN(new_n945));
  INV_X1    g0745(.A(new_n906), .ZN(new_n946));
  INV_X1    g0746(.A(new_n825), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n946), .B1(new_n838), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n898), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n634), .A2(new_n635), .A3(new_n885), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n945), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n722), .A2(new_n642), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n641), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n951), .B(new_n953), .Z(new_n954));
  NAND2_X1  g0754(.A1(new_n940), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n940), .A2(new_n954), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT110), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n955), .B1(new_n490), .B2(new_n681), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n956), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n959), .A2(KEYINPUT110), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n879), .B1(new_n958), .B2(new_n960), .ZN(G367));
  NAND2_X1  g0761(.A1(new_n233), .A2(new_n763), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n773), .B1(new_n709), .B2(new_n562), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n866), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n650), .A2(new_n652), .A3(new_n689), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n656), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n654), .A2(new_n965), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT46), .ZN(new_n969));
  NOR3_X1   g0769(.A1(new_n795), .A2(new_n969), .A3(new_n590), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(new_n777), .B2(G303), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n969), .B1(new_n795), .B2(new_n590), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n971), .B(new_n972), .C1(new_n787), .C2(new_n782), .ZN(new_n973));
  INV_X1    g0773(.A(G317), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n329), .B1(new_n784), .B2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n789), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n975), .B1(new_n976), .B2(G97), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n977), .B1(new_n421), .B2(new_n793), .C1(new_n794), .C2(new_n801), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n973), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n780), .B2(new_n800), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT114), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n778), .A2(new_n856), .B1(new_n201), .B2(new_n782), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n792), .A2(G68), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n983), .B1(new_n202), .B2(new_n795), .C1(new_n855), .C2(new_n784), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT115), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n248), .B1(new_n789), .B2(new_n250), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n986), .A2(new_n987), .B1(new_n801), .B2(new_n811), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(new_n986), .B2(new_n987), .ZN(new_n989));
  INV_X1    g0789(.A(G143), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n985), .B(new_n989), .C1(new_n990), .C2(new_n800), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n981), .A2(new_n991), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT47), .Z(new_n993));
  INV_X1    g0793(.A(new_n771), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n964), .B1(new_n821), .B2(new_n968), .C1(new_n993), .C2(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT111), .Z(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(KEYINPUT113), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n645), .B1(new_n548), .B2(new_n690), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n666), .A2(new_n689), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n704), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n705), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n701), .A2(new_n1001), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(KEYINPUT42), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT42), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n701), .A2(new_n1001), .A3(new_n1007), .A4(new_n1004), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n546), .B1(new_n999), .B2(new_n501), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n690), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1006), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT112), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1006), .A2(KEYINPUT112), .A3(new_n1008), .A4(new_n1010), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n998), .A2(new_n1003), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1003), .B1(new_n998), .B2(new_n1016), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n1018), .A2(new_n1019), .B1(KEYINPUT113), .B2(new_n997), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1019), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n997), .A2(KEYINPUT113), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1021), .A2(new_n1022), .A3(new_n1017), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1002), .A2(new_n706), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT44), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1025), .B(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n707), .A2(KEYINPUT45), .A3(new_n1001), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT45), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n1002), .B2(new_n706), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1027), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n703), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1027), .A2(new_n704), .A3(new_n1031), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n701), .B(new_n1004), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(new_n696), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n751), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n751), .B1(new_n1035), .B2(new_n1038), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n710), .B(KEYINPUT41), .Z(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n754), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n995), .B1(new_n1024), .B2(new_n1042), .ZN(G387));
  NAND2_X1  g0843(.A1(new_n1037), .A2(new_n754), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(G303), .A2(new_n853), .B1(new_n777), .B2(G317), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n780), .B2(new_n801), .C1(new_n800), .C2(new_n779), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT48), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n843), .A2(G294), .B1(new_n792), .B2(G283), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT49), .ZN(new_n1052));
  AND2_X1   g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n329), .B1(new_n798), .B2(new_n784), .C1(new_n789), .C2(new_n590), .ZN(new_n1055));
  OR3_X1    g0855(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n778), .A2(new_n201), .B1(new_n203), .B2(new_n782), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n248), .B1(new_n856), .B2(new_n784), .C1(new_n789), .C2(new_n542), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n793), .A2(new_n436), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n795), .A2(new_n250), .ZN(new_n1060));
  NOR4_X1   g0860(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1061), .B1(new_n811), .B2(new_n799), .C1(new_n319), .C2(new_n801), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n994), .B1(new_n1056), .B2(new_n1062), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n759), .A2(new_n712), .B1(G107), .B2(new_n208), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n712), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n476), .B1(new_n203), .B2(new_n439), .C1(new_n1065), .C2(KEYINPUT116), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(KEYINPUT116), .B2(new_n1065), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n434), .A2(G50), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT50), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n764), .B1(new_n238), .B2(new_n262), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1064), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n758), .B1(new_n773), .B2(new_n1072), .C1(new_n701), .C2(new_n821), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1038), .A2(new_n710), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n751), .A2(new_n1037), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1044), .B1(new_n1063), .B2(new_n1073), .C1(new_n1074), .C2(new_n1075), .ZN(G393));
  INV_X1    g0876(.A(new_n1034), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n704), .B1(new_n1027), .B2(new_n1031), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1038), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n711), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1035), .A2(KEYINPUT118), .A3(new_n1038), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(KEYINPUT118), .B1(new_n1035), .B2(new_n1038), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1081), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1002), .A2(new_n770), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n243), .A2(new_n764), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n772), .B1(new_n542), .B2(new_n208), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n758), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n778), .A2(new_n780), .B1(new_n974), .B2(new_n799), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT52), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n329), .B1(new_n779), .B2(new_n784), .C1(new_n789), .C2(new_n421), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n793), .A2(new_n590), .B1(new_n787), .B2(new_n795), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1092), .B(new_n1093), .C1(G294), .C2(new_n853), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1091), .B(new_n1094), .C1(new_n601), .C2(new_n801), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n815), .A2(G150), .B1(new_n777), .B2(G159), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT117), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(KEYINPUT51), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n329), .B(new_n842), .C1(G143), .C2(new_n785), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n1099), .B1(new_n203), .B2(new_n795), .C1(new_n439), .C2(new_n793), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n782), .A2(new_n434), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1098), .B(new_n1102), .C1(new_n201), .C2(new_n801), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1097), .A2(KEYINPUT51), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1095), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1089), .B1(new_n1105), .B2(new_n771), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1079), .A2(new_n754), .B1(new_n1086), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1085), .A2(new_n1107), .ZN(G390));
  OAI21_X1  g0908(.A(new_n936), .B1(new_n746), .B2(KEYINPUT31), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n741), .A2(new_n723), .ZN(new_n1110));
  OAI211_X1 g0910(.A(G330), .B(new_n830), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n946), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n937), .A2(G330), .A3(new_n830), .A4(new_n906), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n838), .A2(new_n947), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n719), .A2(new_n690), .A3(new_n830), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n1117), .A2(new_n947), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1112), .A2(new_n1113), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n748), .A2(new_n448), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n641), .B(new_n1121), .C1(new_n722), .C2(new_n642), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(KEYINPUT119), .B1(new_n948), .B2(new_n944), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n942), .B1(new_n941), .B2(new_n898), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n831), .B1(new_n657), .B2(new_n676), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n906), .B1(new_n1127), .B2(new_n825), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT119), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1128), .A2(new_n1129), .A3(new_n943), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1125), .A2(new_n1126), .A3(new_n1130), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n943), .B(new_n921), .C1(new_n1118), .C2(new_n946), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n1131), .A2(new_n1113), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1113), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1124), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1113), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1131), .A2(new_n1113), .A3(new_n1132), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n1112), .A2(new_n1113), .A3(new_n1118), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1112), .A2(new_n1113), .B1(new_n947), .B2(new_n838), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1142), .A2(new_n1122), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1138), .A2(new_n1139), .A3(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1135), .A2(new_n1144), .A3(new_n710), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n867), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n815), .A2(G128), .B1(new_n777), .B2(G132), .ZN(new_n1147));
  XOR2_X1   g0947(.A(new_n1147), .B(KEYINPUT120), .Z(new_n1148));
  OAI21_X1  g0948(.A(KEYINPUT53), .B1(new_n795), .B2(new_n856), .ZN(new_n1149));
  INV_X1    g0949(.A(G125), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n248), .B1(new_n1150), .B2(new_n784), .C1(new_n789), .C2(new_n201), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G159), .B2(new_n792), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n795), .A2(KEYINPUT53), .A3(new_n856), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT54), .B(G143), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1153), .B1(new_n853), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n801), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(G137), .ZN(new_n1158));
  AND4_X1   g0958(.A1(new_n1149), .A2(new_n1152), .A3(new_n1156), .A4(new_n1158), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n778), .A2(new_n590), .B1(new_n542), .B2(new_n782), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n329), .B1(new_n794), .B2(new_n784), .C1(new_n795), .C2(new_n346), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n793), .A2(new_n439), .B1(new_n203), .B2(new_n789), .ZN(new_n1162));
  NOR3_X1   g0962(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(G107), .A2(new_n1157), .B1(new_n815), .B2(G283), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n1148), .A2(new_n1159), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n758), .B1(new_n291), .B2(new_n1146), .C1(new_n1165), .C2(new_n994), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(new_n1126), .B2(new_n768), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1167), .B1(new_n1168), .B2(new_n754), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1145), .A2(new_n1169), .ZN(G378));
  OAI21_X1  g0970(.A(new_n983), .B1(new_n799), .B2(new_n590), .ZN(new_n1171));
  XOR2_X1   g0971(.A(new_n1171), .B(KEYINPUT121), .Z(new_n1172));
  OAI22_X1  g0972(.A1(new_n778), .A2(new_n421), .B1(new_n436), .B2(new_n782), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n248), .A2(G41), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n787), .B2(new_n784), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n789), .A2(new_n202), .ZN(new_n1176));
  OR3_X1    g0976(.A1(new_n1175), .A2(new_n1060), .A3(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1173), .A2(new_n1177), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1172), .B(new_n1178), .C1(new_n542), .C2(new_n801), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n201), .B1(G33), .B2(G41), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n1180), .A2(KEYINPUT58), .B1(new_n1174), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(KEYINPUT122), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1180), .A2(KEYINPUT58), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n1150), .A2(new_n799), .B1(new_n801), .B2(new_n861), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n777), .A2(G128), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n792), .A2(G150), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n843), .A2(new_n1155), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1185), .B(new_n1189), .C1(G137), .C2(new_n853), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1191), .A2(KEYINPUT59), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(KEYINPUT59), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n976), .A2(G159), .ZN(new_n1194));
  AOI211_X1 g0994(.A(G33), .B(G41), .C1(new_n785), .C2(G124), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1183), .B(new_n1184), .C1(new_n1192), .C2(new_n1196), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1182), .A2(KEYINPUT122), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n771), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n710), .B(new_n754), .C1(new_n201), .C2(new_n867), .ZN(new_n1200));
  XOR2_X1   g1000(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1201));
  XNOR2_X1  g1001(.A(new_n315), .B(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n296), .A2(new_n885), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT123), .ZN(new_n1204));
  XOR2_X1   g1004(.A(new_n1202), .B(new_n1204), .Z(new_n1205));
  OAI211_X1 g1005(.A(new_n1199), .B(new_n1200), .C1(new_n1205), .C2(new_n769), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n898), .A2(new_n908), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(new_n925), .ZN(new_n1209));
  AND4_X1   g1009(.A1(KEYINPUT109), .A2(new_n908), .A3(new_n921), .A4(KEYINPUT40), .ZN(new_n1210));
  AOI21_X1  g1010(.A(KEYINPUT109), .B1(new_n929), .B2(new_n908), .ZN(new_n1211));
  OAI211_X1 g1011(.A(G330), .B(new_n1209), .C1(new_n1210), .C2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1205), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n924), .A2(new_n930), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1215), .A2(new_n1205), .A3(G330), .A4(new_n1209), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n951), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n951), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1214), .A2(new_n1219), .A3(new_n1216), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1207), .B1(new_n1221), .B2(new_n754), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n1214), .A2(new_n1219), .A3(new_n1216), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1219), .B1(new_n1214), .B2(new_n1216), .ZN(new_n1224));
  OAI21_X1  g1024(.A(KEYINPUT57), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1122), .B1(new_n1168), .B2(new_n1143), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n710), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1144), .A2(new_n1123), .ZN(new_n1228));
  AOI21_X1  g1028(.A(KEYINPUT57), .B1(new_n1221), .B2(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1222), .B1(new_n1227), .B2(new_n1229), .ZN(G375));
  NAND2_X1  g1030(.A1(new_n946), .A2(new_n768), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n758), .B1(G68), .B2(new_n1146), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n248), .B(new_n1059), .C1(G303), .C2(new_n785), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(G107), .A2(new_n853), .B1(new_n777), .B2(G283), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n843), .A2(G97), .B1(new_n976), .B2(G77), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n590), .A2(new_n801), .B1(new_n799), .B2(new_n794), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n329), .B(new_n1176), .C1(G128), .C2(new_n785), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n843), .A2(G159), .B1(new_n792), .B2(G50), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(G150), .A2(new_n853), .B1(new_n777), .B2(G137), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n861), .A2(new_n799), .B1(new_n801), .B2(new_n1154), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n1236), .A2(new_n1237), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1232), .B1(new_n1243), .B2(new_n771), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n1120), .A2(new_n754), .B1(new_n1231), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1124), .A2(new_n1041), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1116), .A2(new_n1122), .A3(new_n1119), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1245), .B1(new_n1246), .B2(new_n1247), .ZN(G381));
  OR4_X1    g1048(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1249), .A2(G387), .A3(G381), .ZN(new_n1250));
  INV_X1    g1050(.A(G378), .ZN(new_n1251));
  INV_X1    g1051(.A(G375), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1250), .A2(new_n1251), .A3(new_n1252), .ZN(G407));
  INV_X1    g1053(.A(G213), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1254), .A2(G343), .ZN(new_n1255));
  XOR2_X1   g1055(.A(new_n1255), .B(KEYINPUT124), .Z(new_n1256));
  NAND3_X1  g1056(.A1(new_n1252), .A2(new_n1251), .A3(new_n1256), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1257), .A2(KEYINPUT125), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1257), .A2(KEYINPUT125), .ZN(new_n1259));
  OAI211_X1 g1059(.A(G213), .B(G407), .C1(new_n1258), .C2(new_n1259), .ZN(G409));
  OAI211_X1 g1060(.A(G378), .B(new_n1222), .C1(new_n1227), .C2(new_n1229), .ZN(new_n1261));
  AND3_X1   g1061(.A1(new_n1221), .A2(new_n1228), .A3(new_n1041), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1206), .B1(new_n1263), .B2(new_n753), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1251), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1261), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1255), .ZN(new_n1267));
  INV_X1    g1067(.A(G384), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1116), .A2(new_n1122), .A3(KEYINPUT60), .A4(new_n1119), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n710), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1247), .ZN(new_n1271));
  OAI21_X1  g1071(.A(KEYINPUT60), .B1(new_n1142), .B2(new_n1122), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1270), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1245), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1268), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1247), .B1(new_n1124), .B2(KEYINPUT60), .ZN(new_n1276));
  OAI211_X1 g1076(.A(G384), .B(new_n1245), .C1(new_n1276), .C2(new_n1270), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1266), .A2(new_n1267), .A3(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT63), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1255), .A2(G2897), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1275), .A2(new_n1277), .A3(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(KEYINPUT126), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT126), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1275), .A2(new_n1287), .A3(new_n1277), .A4(new_n1284), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1278), .A2(G2897), .A3(new_n1256), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1283), .A2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1256), .B1(new_n1261), .B2(new_n1265), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1294), .A2(KEYINPUT63), .A3(new_n1279), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1085), .A2(new_n1107), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(G387), .A2(new_n1296), .ZN(new_n1297));
  XNOR2_X1  g1097(.A(G393), .B(new_n823), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n753), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1300), .A2(new_n1023), .A3(new_n1020), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1301), .A2(G390), .A3(new_n995), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1297), .A2(new_n1298), .A3(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1298), .B1(new_n1297), .B2(new_n1302), .ZN(new_n1304));
  NOR3_X1   g1104(.A1(new_n1303), .A2(new_n1304), .A3(KEYINPUT61), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1282), .A2(new_n1293), .A3(new_n1295), .A4(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT61), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1307), .B1(new_n1294), .B2(new_n1291), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT62), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1280), .A2(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1294), .A2(KEYINPUT62), .A3(new_n1279), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1308), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1306), .B1(new_n1312), .B2(new_n1313), .ZN(G405));
  INV_X1    g1114(.A(new_n1298), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(G387), .A2(new_n1296), .ZN(new_n1316));
  AOI21_X1  g1116(.A(G390), .B1(new_n1301), .B2(new_n995), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1315), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1297), .A2(new_n1302), .A3(new_n1298), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1318), .B(new_n1319), .C1(KEYINPUT127), .C2(new_n1279), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1279), .A2(KEYINPUT127), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1321), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1320), .A2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT127), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1261), .B1(new_n1324), .B2(new_n1278), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1325), .B1(new_n1251), .B2(G375), .ZN(new_n1326));
  XNOR2_X1  g1126(.A(new_n1323), .B(new_n1326), .ZN(G402));
endmodule


