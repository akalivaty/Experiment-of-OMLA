//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 1 1 1 1 0 0 0 0 1 1 1 1 1 0 0 0 1 1 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n614, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972;
  INV_X1    g000(.A(G125), .ZN(new_n187));
  INV_X1    g001(.A(G140), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  NAND2_X1  g003(.A1(G125), .A2(G140), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT16), .ZN(new_n192));
  OR3_X1    g006(.A1(new_n187), .A2(KEYINPUT16), .A3(G140), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n192), .A2(G146), .A3(new_n193), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G119), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(G128), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT68), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(new_n199), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT68), .A2(G119), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n200), .B1(new_n204), .B2(G128), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT23), .ZN(new_n206));
  OR3_X1    g020(.A1(new_n204), .A2(KEYINPUT23), .A3(G128), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(G110), .A3(new_n207), .ZN(new_n208));
  XOR2_X1   g022(.A(KEYINPUT24), .B(G110), .Z(new_n209));
  NAND2_X1  g023(.A1(new_n205), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n198), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n191), .A2(new_n195), .ZN(new_n212));
  AOI21_X1  g026(.A(G110), .B1(new_n206), .B2(new_n207), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n205), .A2(new_n209), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n197), .A2(KEYINPUT74), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT74), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n192), .A2(new_n217), .A3(G146), .A4(new_n193), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n211), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G953), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(G221), .A3(G234), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n222), .B(KEYINPUT22), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n223), .B(G137), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G902), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n211), .B(new_n224), .C1(new_n215), .C2(new_n219), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(KEYINPUT75), .A3(KEYINPUT25), .ZN(new_n230));
  INV_X1    g044(.A(G217), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n231), .B1(G234), .B2(new_n227), .ZN(new_n232));
  XOR2_X1   g046(.A(KEYINPUT75), .B(KEYINPUT25), .Z(new_n233));
  NAND4_X1  g047(.A1(new_n226), .A2(new_n227), .A3(new_n228), .A4(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n230), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  AND2_X1   g049(.A1(new_n226), .A2(new_n228), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n232), .A2(G902), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT69), .ZN(new_n242));
  AND2_X1   g056(.A1(KEYINPUT68), .A2(G119), .ZN(new_n243));
  NOR2_X1   g057(.A1(KEYINPUT68), .A2(G119), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n242), .B(G116), .C1(new_n243), .C2(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT2), .B(G113), .ZN(new_n246));
  INV_X1    g060(.A(G116), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n247), .B1(new_n202), .B2(new_n203), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT69), .B1(new_n199), .B2(G116), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n245), .B(new_n246), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(G116), .B1(new_n243), .B2(new_n244), .ZN(new_n252));
  INV_X1    g066(.A(new_n249), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n246), .B1(new_n254), .B2(new_n245), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n241), .B1(new_n251), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n245), .B1(new_n248), .B2(new_n249), .ZN(new_n257));
  INV_X1    g071(.A(new_n246), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(KEYINPUT70), .A3(new_n250), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT11), .ZN(new_n262));
  INV_X1    g076(.A(G134), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n262), .B1(new_n263), .B2(G137), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT65), .ZN(new_n265));
  INV_X1    g079(.A(G137), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n265), .B1(new_n266), .B2(G134), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(KEYINPUT11), .A3(G134), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n263), .A2(KEYINPUT65), .A3(G137), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n264), .A2(new_n267), .A3(new_n268), .A4(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n270), .B(G131), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n195), .A2(G143), .ZN(new_n272));
  INV_X1    g086(.A(G143), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G146), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT0), .ZN(new_n276));
  INV_X1    g090(.A(G128), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(new_n277), .A3(KEYINPUT64), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n278), .B1(new_n276), .B2(new_n277), .ZN(new_n279));
  AOI21_X1  g093(.A(KEYINPUT64), .B1(new_n276), .B2(new_n277), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n275), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n272), .B(new_n274), .C1(new_n276), .C2(new_n277), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI211_X1 g097(.A(KEYINPUT66), .B(KEYINPUT1), .C1(new_n273), .C2(G146), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G128), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT66), .B1(new_n272), .B2(KEYINPUT1), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n275), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT67), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n275), .A2(new_n277), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT1), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI211_X1 g106(.A(KEYINPUT67), .B(new_n275), .C1(new_n285), .C2(new_n286), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n289), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n270), .A2(G131), .ZN(new_n295));
  INV_X1    g109(.A(G131), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n266), .A2(G134), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n263), .A2(G137), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n296), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  AOI221_X4 g114(.A(KEYINPUT30), .B1(new_n271), .B2(new_n283), .C1(new_n294), .C2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT30), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n294), .A2(new_n300), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n271), .A2(new_n283), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n261), .B1(new_n301), .B2(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n307), .B(G101), .ZN(new_n308));
  OR2_X1    g122(.A1(KEYINPUT71), .A2(G237), .ZN(new_n309));
  NAND2_X1  g123(.A1(KEYINPUT71), .A2(G237), .ZN(new_n310));
  AOI21_X1  g124(.A(G953), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G210), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n308), .B(new_n312), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n303), .A2(new_n256), .A3(new_n260), .A4(new_n304), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n306), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT31), .ZN(new_n316));
  INV_X1    g130(.A(new_n313), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT72), .B(KEYINPUT28), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n303), .A2(new_n304), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n261), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n318), .B1(new_n320), .B2(new_n314), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT28), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n314), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n317), .B1(new_n321), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT31), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n306), .A2(new_n326), .A3(new_n313), .A4(new_n314), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n316), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT73), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G472), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n316), .A2(new_n325), .A3(KEYINPUT73), .A4(new_n327), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n330), .A2(new_n331), .A3(new_n227), .A4(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT32), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n320), .A2(new_n314), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n323), .B1(new_n337), .B2(new_n322), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n313), .A2(KEYINPUT29), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n227), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n313), .B1(new_n321), .B2(new_n324), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n306), .A2(new_n317), .A3(new_n314), .ZN(new_n342));
  AOI21_X1  g156(.A(KEYINPUT29), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(G472), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n344), .B1(new_n333), .B2(new_n334), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n240), .B1(new_n336), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n294), .A2(new_n187), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n283), .A2(G125), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n221), .A2(G224), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n349), .B(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G104), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT3), .B1(new_n352), .B2(G107), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT3), .ZN(new_n354));
  INV_X1    g168(.A(G107), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n355), .A3(G104), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n352), .A2(G107), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n353), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G101), .ZN(new_n359));
  INV_X1    g173(.A(G101), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n353), .A2(new_n356), .A3(new_n360), .A4(new_n357), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n359), .A2(KEYINPUT4), .A3(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT4), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n358), .A2(new_n363), .A3(G101), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n261), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT5), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n204), .A2(new_n368), .A3(G116), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n370), .B1(KEYINPUT5), .B2(new_n257), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n255), .B1(new_n371), .B2(G113), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT76), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(new_n355), .A3(G104), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT76), .B1(new_n355), .B2(G104), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n352), .A2(G107), .ZN(new_n376));
  OAI211_X1 g190(.A(G101), .B(new_n374), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n377), .A2(new_n361), .A3(KEYINPUT77), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT77), .B1(new_n377), .B2(new_n361), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n372), .A2(new_n380), .ZN(new_n381));
  XOR2_X1   g195(.A(G110), .B(G122), .Z(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n367), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n257), .A2(KEYINPUT5), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(G113), .A3(new_n369), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n386), .A2(new_n380), .A3(new_n259), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n365), .B1(new_n256), .B2(new_n260), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n382), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n384), .A2(new_n389), .A3(KEYINPUT6), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT82), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n383), .B1(new_n367), .B2(new_n381), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT6), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n393), .B(new_n382), .C1(new_n387), .C2(new_n388), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n395), .A2(KEYINPUT82), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n351), .B(new_n390), .C1(new_n394), .C2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT83), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n349), .A2(new_n350), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n377), .A2(new_n361), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(KEYINPUT85), .B1(new_n372), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT84), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n386), .A2(new_n259), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n404), .B1(new_n405), .B2(new_n401), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT85), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n405), .A2(new_n407), .A3(new_n401), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n372), .A2(KEYINPUT84), .A3(new_n402), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n403), .A2(new_n406), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  XOR2_X1   g224(.A(new_n382), .B(KEYINPUT8), .Z(new_n411));
  AOI21_X1  g225(.A(new_n400), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n349), .A2(KEYINPUT7), .A3(new_n350), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT86), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n349), .A2(KEYINPUT86), .A3(KEYINPUT7), .A4(new_n350), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OR2_X1    g231(.A1(new_n349), .A2(KEYINPUT7), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n412), .A2(new_n417), .A3(new_n384), .A4(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n392), .A2(new_n391), .A3(new_n393), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n395), .A2(KEYINPUT82), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n422), .A2(KEYINPUT83), .A3(new_n351), .A4(new_n390), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n399), .A2(new_n227), .A3(new_n419), .A4(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(G210), .B1(G237), .B2(G902), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT87), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n419), .A2(new_n227), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n429), .A2(new_n425), .A3(new_n399), .A4(new_n423), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n427), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(G475), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n309), .A2(new_n310), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(G214), .A3(new_n221), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT88), .ZN(new_n435));
  OAI21_X1  g249(.A(KEYINPUT89), .B1(new_n435), .B2(G143), .ZN(new_n436));
  OR2_X1    g250(.A1(KEYINPUT89), .A2(G143), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n436), .B1(new_n311), .B2(G214), .ZN(new_n440));
  NOR3_X1   g254(.A1(new_n439), .A2(new_n296), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT17), .ZN(new_n442));
  INV_X1    g256(.A(new_n198), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n296), .B1(new_n439), .B2(new_n440), .ZN(new_n444));
  INV_X1    g258(.A(new_n436), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n434), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n311), .A2(G214), .A3(new_n436), .A4(new_n437), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n447), .A3(G131), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n442), .B(new_n443), .C1(new_n449), .C2(KEYINPUT17), .ZN(new_n450));
  XOR2_X1   g264(.A(G113), .B(G122), .Z(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(KEYINPUT94), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(new_n352), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n446), .A2(new_n447), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT91), .ZN(new_n456));
  AOI22_X1  g270(.A1(new_n455), .A2(new_n456), .B1(KEYINPUT18), .B2(G131), .ZN(new_n457));
  NAND2_X1  g271(.A1(KEYINPUT18), .A2(G131), .ZN(new_n458));
  AOI211_X1 g272(.A(KEYINPUT91), .B(new_n458), .C1(new_n446), .C2(new_n447), .ZN(new_n459));
  INV_X1    g273(.A(new_n191), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G146), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n461), .A2(KEYINPUT90), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n212), .B1(new_n461), .B2(KEYINPUT90), .ZN(new_n463));
  OAI22_X1  g277(.A1(new_n457), .A2(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n450), .A2(new_n454), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n219), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT92), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n191), .A2(new_n467), .A3(KEYINPUT19), .ZN(new_n468));
  OR2_X1    g282(.A1(new_n467), .A2(KEYINPUT19), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(KEYINPUT19), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n469), .A2(new_n189), .A3(new_n190), .A4(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(G146), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(KEYINPUT93), .ZN(new_n473));
  OR2_X1    g287(.A1(new_n472), .A2(KEYINPUT93), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n449), .A2(new_n466), .A3(new_n473), .A4(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n454), .B1(new_n475), .B2(new_n464), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n432), .B(new_n227), .C1(new_n465), .C2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT20), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n454), .B1(new_n450), .B2(new_n464), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n227), .B1(new_n465), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(G475), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n475), .A2(new_n464), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n453), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n450), .A2(new_n454), .A3(new_n464), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n486), .A2(KEYINPUT20), .A3(new_n432), .A4(new_n227), .ZN(new_n487));
  INV_X1    g301(.A(G952), .ZN(new_n488));
  AOI211_X1 g302(.A(G953), .B(new_n488), .C1(G234), .C2(G237), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  AOI211_X1 g304(.A(new_n227), .B(new_n221), .C1(G234), .C2(G237), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  XOR2_X1   g306(.A(KEYINPUT21), .B(G898), .Z(new_n493));
  OAI21_X1  g307(.A(new_n490), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n479), .A2(new_n482), .A3(new_n487), .A4(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n247), .A2(G122), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n247), .A2(G122), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n496), .B1(KEYINPUT14), .B2(new_n497), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n498), .B(KEYINPUT98), .C1(KEYINPUT14), .C2(new_n497), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n499), .B(G107), .C1(KEYINPUT98), .C2(new_n498), .ZN(new_n500));
  INV_X1    g314(.A(new_n496), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n501), .A2(new_n497), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n355), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n273), .A2(G128), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n277), .A2(G143), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(KEYINPUT97), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n507), .A2(new_n263), .ZN(new_n508));
  OR2_X1    g322(.A1(new_n506), .A2(KEYINPUT97), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n506), .A2(KEYINPUT97), .ZN(new_n510));
  AOI21_X1  g324(.A(G134), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n500), .B(new_n503), .C1(new_n508), .C2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(KEYINPUT13), .B1(new_n273), .B2(G128), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT95), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n513), .B(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT13), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n515), .B(new_n505), .C1(new_n516), .C2(new_n504), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n517), .A2(KEYINPUT96), .A3(G134), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n502), .B(new_n355), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n507), .A2(new_n263), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n521), .A2(KEYINPUT96), .B1(new_n517), .B2(G134), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n512), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  XOR2_X1   g337(.A(KEYINPUT9), .B(G234), .Z(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NOR3_X1   g339(.A1(new_n525), .A2(new_n231), .A3(G953), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n512), .B(new_n526), .C1(new_n520), .C2(new_n522), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n227), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT15), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n532), .A3(G478), .ZN(new_n533));
  INV_X1    g347(.A(G478), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n530), .B(new_n227), .C1(KEYINPUT15), .C2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n495), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(G221), .B1(new_n525), .B2(G902), .ZN(new_n538));
  XOR2_X1   g352(.A(KEYINPUT79), .B(G469), .Z(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT10), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n272), .A2(KEYINPUT1), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G128), .ZN(new_n543));
  AOI22_X1  g357(.A1(new_n290), .A2(new_n291), .B1(new_n543), .B2(new_n275), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n541), .B1(new_n544), .B2(new_n401), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n283), .A2(new_n362), .A3(new_n364), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n270), .B(new_n296), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n294), .A2(new_n380), .A3(KEYINPUT10), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT80), .ZN(new_n551));
  XNOR2_X1  g365(.A(G110), .B(G140), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n221), .A2(G227), .ZN(new_n553));
  XOR2_X1   g367(.A(new_n552), .B(new_n553), .Z(new_n554));
  AND3_X1   g368(.A1(new_n550), .A2(new_n551), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n551), .B1(new_n550), .B2(new_n554), .ZN(new_n556));
  OR2_X1    g370(.A1(new_n544), .A2(new_n401), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n289), .A2(new_n292), .A3(new_n293), .A4(new_n401), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(KEYINPUT12), .B1(new_n559), .B2(new_n271), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT12), .ZN(new_n561));
  AOI211_X1 g375(.A(new_n561), .B(new_n548), .C1(new_n557), .C2(new_n558), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NOR3_X1   g377(.A1(new_n555), .A2(new_n556), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n548), .B1(new_n547), .B2(new_n549), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n554), .B1(new_n566), .B2(new_n550), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n227), .B(new_n540), .C1(new_n564), .C2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(G469), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n550), .A2(new_n554), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT78), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n550), .A2(KEYINPUT78), .A3(new_n554), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n572), .A2(new_n566), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n554), .ZN(new_n575));
  INV_X1    g389(.A(new_n550), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n575), .B1(new_n563), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(G902), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n568), .B1(new_n569), .B2(new_n578), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n537), .A2(new_n538), .A3(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(G214), .B1(G237), .B2(G902), .ZN(new_n581));
  XOR2_X1   g395(.A(new_n581), .B(KEYINPUT81), .Z(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n424), .A2(KEYINPUT87), .A3(new_n426), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n431), .A2(new_n580), .A3(new_n583), .A4(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n346), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(new_n360), .ZN(G3));
  INV_X1    g401(.A(KEYINPUT99), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n588), .B1(new_n424), .B2(new_n426), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n427), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n424), .A2(new_n588), .A3(new_n426), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n582), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n530), .A2(KEYINPUT33), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT33), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n528), .A2(new_n594), .A3(new_n529), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n593), .A2(G478), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n530), .A2(new_n534), .A3(new_n227), .ZN(new_n597));
  NAND2_X1  g411(.A1(G478), .A2(G902), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n479), .A2(new_n482), .A3(new_n487), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n592), .A2(new_n494), .A3(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n330), .A2(new_n227), .A3(new_n332), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(G472), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n333), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n579), .A2(new_n240), .A3(new_n538), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n602), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(KEYINPUT34), .B(G104), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G6));
  INV_X1    g424(.A(new_n495), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n592), .A2(new_n536), .A3(new_n611), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n612), .A2(new_n605), .A3(new_n607), .ZN(new_n613));
  XNOR2_X1  g427(.A(KEYINPUT35), .B(G107), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G9));
  AND3_X1   g429(.A1(new_n431), .A2(new_n583), .A3(new_n584), .ZN(new_n616));
  INV_X1    g430(.A(new_n605), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n616), .A2(new_n580), .A3(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n225), .A2(KEYINPUT36), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n220), .B(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n237), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n235), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT100), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G110), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT101), .B(KEYINPUT37), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G12));
  INV_X1    g441(.A(new_n536), .ZN(new_n628));
  INV_X1    g442(.A(G900), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n489), .B1(new_n491), .B2(new_n629), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n628), .A2(new_n600), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n592), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT102), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n592), .A2(KEYINPUT102), .A3(new_n631), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n330), .A2(new_n332), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n636), .A2(KEYINPUT32), .A3(new_n331), .A4(new_n227), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n637), .A2(new_n335), .A3(new_n344), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n579), .A2(new_n538), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n623), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n634), .A2(new_n635), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G128), .ZN(G30));
  AND2_X1   g458(.A1(new_n431), .A2(new_n584), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT38), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n630), .B(KEYINPUT39), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n639), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT40), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n582), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n646), .B(new_n650), .C1(new_n649), .C2(new_n648), .ZN(new_n651));
  INV_X1    g465(.A(new_n623), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n306), .A2(new_n314), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n313), .ZN(new_n654));
  AOI21_X1  g468(.A(G902), .B1(new_n337), .B2(new_n317), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n331), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n637), .A2(new_n335), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(KEYINPUT103), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT103), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n637), .A2(new_n660), .A3(new_n335), .A4(new_n657), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n662), .A2(new_n536), .A3(new_n600), .ZN(new_n663));
  OR3_X1    g477(.A1(new_n651), .A2(new_n652), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G143), .ZN(G45));
  INV_X1    g479(.A(new_n630), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n599), .A2(new_n600), .A3(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n592), .A2(new_n638), .A3(new_n640), .A4(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G146), .ZN(G48));
  INV_X1    g484(.A(new_n538), .ZN(new_n671));
  INV_X1    g485(.A(new_n568), .ZN(new_n672));
  OR3_X1    g486(.A1(new_n555), .A2(new_n556), .A3(new_n563), .ZN(new_n673));
  INV_X1    g487(.A(new_n567), .ZN(new_n674));
  AOI21_X1  g488(.A(G902), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  OR2_X1    g489(.A1(new_n675), .A2(KEYINPUT104), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n569), .B1(new_n675), .B2(KEYINPUT104), .ZN(new_n677));
  AOI211_X1 g491(.A(new_n671), .B(new_n672), .C1(new_n676), .C2(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n638), .A2(new_n240), .A3(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n602), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT41), .B(G113), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G15));
  INV_X1    g496(.A(new_n679), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n592), .A2(new_n536), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n683), .A2(new_n684), .A3(new_n685), .A4(new_n611), .ZN(new_n686));
  OAI21_X1  g500(.A(KEYINPUT105), .B1(new_n612), .B2(new_n679), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G116), .ZN(G18));
  NAND4_X1  g503(.A1(new_n592), .A2(new_n537), .A3(new_n652), .A4(new_n678), .ZN(new_n690));
  INV_X1    g504(.A(new_n638), .ZN(new_n691));
  OR3_X1    g505(.A1(new_n690), .A2(KEYINPUT106), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g506(.A(KEYINPUT106), .B1(new_n690), .B2(new_n691), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G119), .ZN(G21));
  NAND2_X1  g509(.A1(new_n590), .A2(new_n591), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n536), .A2(new_n600), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT110), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n696), .A2(new_n583), .A3(new_n494), .A4(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(G472), .A2(G902), .ZN(new_n700));
  OAI211_X1 g514(.A(KEYINPUT107), .B(new_n323), .C1(new_n337), .C2(new_n322), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n322), .B1(new_n320), .B2(new_n314), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n702), .B1(new_n703), .B2(new_n324), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n701), .A2(new_n704), .A3(new_n317), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n316), .A2(new_n327), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n700), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT108), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT108), .ZN(new_n709));
  OAI211_X1 g523(.A(new_n709), .B(new_n700), .C1(new_n705), .C2(new_n706), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g525(.A(KEYINPUT109), .B(G472), .Z(new_n712));
  NAND2_X1  g526(.A1(new_n603), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n678), .A2(new_n711), .A3(new_n240), .A4(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n699), .A2(new_n714), .ZN(new_n715));
  XOR2_X1   g529(.A(new_n715), .B(G122), .Z(G24));
  AND4_X1   g530(.A1(new_n668), .A2(new_n713), .A3(new_n710), .A4(new_n708), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n592), .A2(new_n717), .A3(new_n652), .A4(new_n678), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G125), .ZN(G27));
  AOI21_X1  g533(.A(new_n582), .B1(new_n431), .B2(new_n584), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n720), .A2(new_n638), .A3(new_n606), .A4(new_n668), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT42), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI211_X1 g537(.A(new_n582), .B(new_n667), .C1(new_n431), .C2(new_n584), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n335), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n333), .A2(KEYINPUT111), .A3(new_n334), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n726), .A2(new_n637), .A3(new_n344), .A4(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n724), .A2(new_n728), .A3(KEYINPUT42), .A4(new_n606), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n723), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(KEYINPUT112), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT112), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n723), .A2(new_n732), .A3(new_n729), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G131), .ZN(G33));
  NAND3_X1  g549(.A1(new_n720), .A2(new_n638), .A3(new_n606), .ZN(new_n736));
  INV_X1    g550(.A(new_n631), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n263), .ZN(G36));
  NAND2_X1  g553(.A1(new_n574), .A2(new_n577), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(KEYINPUT45), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(G469), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT113), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n741), .A2(KEYINPUT113), .A3(G469), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(G469), .A2(G902), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT114), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT46), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  AOI22_X1  g565(.A1(new_n744), .A2(new_n745), .B1(G469), .B2(G902), .ZN(new_n752));
  OAI21_X1  g566(.A(KEYINPUT114), .B1(new_n752), .B2(KEYINPUT46), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n672), .B1(new_n752), .B2(KEYINPUT46), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n751), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n538), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(new_n647), .ZN(new_n757));
  INV_X1    g571(.A(new_n720), .ZN(new_n758));
  INV_X1    g572(.A(new_n600), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n599), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT43), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n762), .A2(new_n605), .A3(new_n652), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT44), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n758), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n757), .B(new_n765), .C1(new_n764), .C2(new_n763), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G137), .ZN(G39));
  INV_X1    g581(.A(KEYINPUT47), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n756), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n755), .A2(KEYINPUT47), .A3(new_n538), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n638), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n239), .A3(new_n724), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G140), .ZN(G42));
  AOI21_X1  g587(.A(new_n672), .B1(new_n676), .B2(new_n677), .ZN(new_n774));
  XOR2_X1   g588(.A(new_n774), .B(KEYINPUT49), .Z(new_n775));
  NOR3_X1   g589(.A1(new_n646), .A2(new_n775), .A3(new_n239), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n662), .A2(new_n582), .A3(new_n671), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n776), .A2(new_n759), .A3(new_n599), .A4(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n738), .B1(new_n731), .B2(new_n733), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n718), .A2(new_n669), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n641), .B1(new_n632), .B2(new_n633), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n782), .B1(new_n635), .B2(new_n783), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n696), .A2(new_n583), .A3(new_n698), .ZN(new_n785));
  INV_X1    g599(.A(new_n622), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n639), .A2(new_n630), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n662), .A2(new_n785), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(KEYINPUT52), .B1(new_n784), .B2(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n718), .A2(new_n669), .ZN(new_n790));
  AND4_X1   g604(.A1(KEYINPUT52), .A2(new_n643), .A3(new_n788), .A4(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n781), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  OAI22_X1  g606(.A1(new_n602), .A2(new_n679), .B1(new_n699), .B2(new_n714), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n793), .B1(new_n686), .B2(new_n687), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n606), .A2(new_n604), .A3(new_n333), .A4(new_n494), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n628), .A2(new_n600), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(new_n616), .A3(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n798), .B1(new_n618), .B2(new_n623), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n431), .A2(new_n583), .A3(new_n584), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n599), .A2(new_n600), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT115), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n800), .A2(new_n795), .A3(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(KEYINPUT116), .B1(new_n803), .B2(new_n586), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n616), .A2(new_n638), .A3(new_n240), .A4(new_n580), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n601), .B(KEYINPUT115), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n796), .A2(new_n616), .A3(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n805), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n799), .B1(new_n804), .B2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n638), .A2(new_n628), .A3(new_n759), .A4(new_n666), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n640), .B(new_n720), .C1(new_n812), .C2(new_n717), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n794), .A2(new_n694), .A3(new_n810), .A4(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n780), .B1(new_n792), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n794), .A2(new_n694), .A3(new_n730), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT119), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n738), .ZN(new_n819));
  AND4_X1   g633(.A1(KEYINPUT53), .A2(new_n810), .A3(new_n819), .A4(new_n813), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n643), .A2(new_n788), .A3(new_n790), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT52), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n643), .A2(new_n788), .A3(new_n790), .A4(KEYINPUT52), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n794), .A2(new_n694), .A3(KEYINPUT119), .A4(new_n730), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n818), .A2(new_n820), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  XOR2_X1   g641(.A(KEYINPUT120), .B(KEYINPUT54), .Z(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n815), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT121), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n815), .A2(new_n827), .A3(KEYINPUT121), .A4(new_n829), .ZN(new_n833));
  AND4_X1   g647(.A1(new_n694), .A2(new_n794), .A3(new_n810), .A4(new_n813), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n834), .A2(new_n781), .A3(new_n825), .A4(new_n779), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT118), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT53), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n837), .B1(new_n792), .B2(new_n814), .ZN(new_n838));
  INV_X1    g652(.A(new_n733), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n732), .B1(new_n723), .B2(new_n729), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n819), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n841), .B1(new_n823), .B2(new_n824), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n842), .A2(new_n843), .A3(new_n834), .A4(new_n779), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n836), .A2(new_n838), .A3(new_n844), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n832), .A2(new_n833), .B1(new_n845), .B2(KEYINPUT54), .ZN(new_n846));
  INV_X1    g660(.A(new_n678), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n646), .A2(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n711), .A2(new_n713), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n240), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n762), .A2(new_n489), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n850), .A2(new_n583), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT50), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n848), .A2(KEYINPUT50), .A3(new_n852), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n758), .A2(new_n851), .A3(new_n847), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n858), .A2(new_n652), .A3(new_n849), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n240), .A2(new_n489), .ZN(new_n861));
  NOR4_X1   g675(.A1(new_n662), .A2(new_n847), .A3(new_n758), .A4(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n599), .A2(new_n600), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n774), .A2(new_n671), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n769), .A2(new_n770), .A3(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n850), .A2(new_n851), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n866), .A2(new_n720), .A3(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n860), .A2(KEYINPUT51), .A3(new_n864), .A4(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT51), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n866), .A2(new_n720), .A3(new_n867), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n857), .A2(new_n864), .A3(new_n859), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n488), .A2(G953), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n867), .A2(new_n592), .A3(new_n678), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n869), .A2(new_n873), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n728), .A2(new_n240), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n858), .A2(new_n877), .ZN(new_n878));
  XOR2_X1   g692(.A(new_n878), .B(KEYINPUT48), .Z(new_n879));
  NOR2_X1   g693(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n862), .A2(new_n601), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n846), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(G952), .A2(G953), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n778), .B1(new_n882), .B2(new_n883), .ZN(G75));
  AOI21_X1  g698(.A(new_n227), .B1(new_n815), .B2(new_n827), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(G210), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT56), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n422), .A2(new_n390), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(new_n351), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(KEYINPUT55), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n891), .B1(KEYINPUT122), .B2(new_n887), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n886), .A2(new_n887), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n892), .B1(new_n886), .B2(new_n887), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n221), .A2(G952), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(G51));
  NAND2_X1  g710(.A1(new_n815), .A2(new_n827), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n828), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n898), .A2(KEYINPUT123), .A3(new_n830), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n897), .A2(new_n900), .A3(new_n828), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n747), .B(KEYINPUT57), .Z(new_n902));
  NAND3_X1  g716(.A1(new_n899), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n673), .A2(new_n674), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n885), .A2(new_n744), .A3(new_n745), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n895), .B1(new_n905), .B2(new_n906), .ZN(G54));
  NAND3_X1  g721(.A1(new_n885), .A2(KEYINPUT58), .A3(G475), .ZN(new_n908));
  INV_X1    g722(.A(new_n486), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n908), .A2(new_n909), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n910), .A2(new_n911), .A3(new_n895), .ZN(G60));
  NAND2_X1  g726(.A1(new_n593), .A2(new_n595), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n598), .B(KEYINPUT59), .Z(new_n915));
  OAI21_X1  g729(.A(new_n914), .B1(new_n846), .B2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n895), .ZN(new_n917));
  INV_X1    g731(.A(new_n915), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n899), .A2(new_n901), .A3(new_n913), .A4(new_n918), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n916), .A2(new_n917), .A3(new_n919), .ZN(G63));
  NAND2_X1  g734(.A1(G217), .A2(G902), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT60), .Z(new_n922));
  NAND3_X1  g736(.A1(new_n897), .A2(new_n620), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n917), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n236), .B1(new_n897), .B2(new_n922), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT61), .ZN(G66));
  AOI21_X1  g741(.A(new_n221), .B1(new_n493), .B2(G224), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n928), .A2(KEYINPUT124), .ZN(new_n929));
  INV_X1    g743(.A(new_n928), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n794), .A2(new_n694), .A3(new_n810), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n930), .B1(new_n931), .B2(G953), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n929), .B1(new_n932), .B2(KEYINPUT124), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n888), .B1(G898), .B2(new_n221), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n933), .B(new_n934), .Z(G69));
  NOR2_X1   g749(.A1(new_n301), .A2(new_n305), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n468), .A2(new_n471), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n936), .B(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n772), .A2(new_n766), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n664), .A2(new_n784), .ZN(new_n940));
  XOR2_X1   g754(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n941));
  NOR2_X1   g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n940), .B1(KEYINPUT125), .B2(KEYINPUT62), .ZN(new_n944));
  INV_X1    g758(.A(new_n346), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n802), .B1(new_n628), .B2(new_n600), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n945), .A2(new_n946), .A3(new_n648), .A4(new_n720), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n943), .A2(new_n944), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n938), .B1(new_n948), .B2(G953), .ZN(new_n949));
  NAND2_X1  g763(.A1(G227), .A2(G900), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(G953), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n772), .A2(new_n766), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n757), .A2(new_n785), .A3(new_n877), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n781), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n952), .A2(new_n784), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n221), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n629), .A2(G953), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT126), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n949), .B(new_n951), .C1(new_n960), .C2(new_n938), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n957), .A2(new_n959), .ZN(new_n962));
  OAI211_X1 g776(.A(G953), .B(new_n950), .C1(new_n962), .C2(new_n938), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n961), .A2(new_n963), .ZN(G72));
  NAND4_X1  g778(.A1(new_n943), .A2(new_n931), .A3(new_n944), .A4(new_n947), .ZN(new_n965));
  NAND2_X1  g779(.A1(G472), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT63), .Z(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT127), .Z(new_n968));
  AOI21_X1  g782(.A(new_n654), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  AND4_X1   g783(.A1(new_n342), .A2(new_n845), .A3(new_n654), .A4(new_n967), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n952), .A2(new_n931), .A3(new_n784), .A4(new_n955), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n342), .B1(new_n971), .B2(new_n968), .ZN(new_n972));
  NOR4_X1   g786(.A1(new_n969), .A2(new_n970), .A3(new_n895), .A4(new_n972), .ZN(G57));
endmodule


