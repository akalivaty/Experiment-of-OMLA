

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592;

  OR2_X1 U327 ( .A1(n420), .A2(n419), .ZN(n421) );
  XNOR2_X1 U328 ( .A(n477), .B(n476), .ZN(n551) );
  XNOR2_X1 U329 ( .A(n475), .B(KEYINPUT48), .ZN(n476) );
  XNOR2_X1 U330 ( .A(n461), .B(n460), .ZN(n509) );
  AND2_X1 U331 ( .A1(G229GAT), .A2(G233GAT), .ZN(n295) );
  INV_X1 U332 ( .A(KEYINPUT91), .ZN(n370) );
  XNOR2_X1 U333 ( .A(n371), .B(n370), .ZN(n372) );
  NOR2_X1 U334 ( .A1(n414), .A2(n524), .ZN(n415) );
  XNOR2_X1 U335 ( .A(n373), .B(n372), .ZN(n376) );
  XNOR2_X1 U336 ( .A(n379), .B(n378), .ZN(n380) );
  NOR2_X1 U337 ( .A1(n417), .A2(n392), .ZN(n552) );
  XNOR2_X1 U338 ( .A(n430), .B(n295), .ZN(n431) );
  XNOR2_X1 U339 ( .A(n381), .B(n380), .ZN(n386) );
  XNOR2_X1 U340 ( .A(n432), .B(n431), .ZN(n436) );
  XNOR2_X1 U341 ( .A(n421), .B(KEYINPUT105), .ZN(n495) );
  XOR2_X1 U342 ( .A(n442), .B(n441), .Z(n576) );
  XNOR2_X1 U343 ( .A(n486), .B(KEYINPUT58), .ZN(n487) );
  XNOR2_X1 U344 ( .A(n462), .B(G29GAT), .ZN(n463) );
  XNOR2_X1 U345 ( .A(n488), .B(n487), .ZN(G1351GAT) );
  XNOR2_X1 U346 ( .A(n464), .B(n463), .ZN(G1328GAT) );
  INV_X1 U347 ( .A(KEYINPUT38), .ZN(n461) );
  XOR2_X1 U348 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n297) );
  NAND2_X1 U349 ( .A1(G231GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U350 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U351 ( .A(n298), .B(KEYINPUT12), .Z(n306) );
  XOR2_X1 U352 ( .A(G155GAT), .B(G78GAT), .Z(n300) );
  XNOR2_X1 U353 ( .A(G22GAT), .B(G211GAT), .ZN(n299) );
  XNOR2_X1 U354 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U355 ( .A(KEYINPUT85), .B(G64GAT), .Z(n302) );
  XNOR2_X1 U356 ( .A(KEYINPUT72), .B(G1GAT), .ZN(n301) );
  XNOR2_X1 U357 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U358 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U359 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U360 ( .A(G8GAT), .B(G183GAT), .Z(n361) );
  XOR2_X1 U361 ( .A(n307), .B(n361), .Z(n310) );
  XOR2_X1 U362 ( .A(G15GAT), .B(G127GAT), .Z(n334) );
  XNOR2_X1 U363 ( .A(G71GAT), .B(G57GAT), .ZN(n308) );
  XNOR2_X1 U364 ( .A(n308), .B(KEYINPUT13), .ZN(n452) );
  XNOR2_X1 U365 ( .A(n334), .B(n452), .ZN(n309) );
  XOR2_X1 U366 ( .A(n310), .B(n309), .Z(n586) );
  INV_X1 U367 ( .A(n586), .ZN(n572) );
  XOR2_X1 U368 ( .A(G92GAT), .B(G106GAT), .Z(n312) );
  XNOR2_X1 U369 ( .A(G134GAT), .B(G218GAT), .ZN(n311) );
  XNOR2_X1 U370 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U371 ( .A(KEYINPUT84), .B(KEYINPUT9), .Z(n314) );
  XNOR2_X1 U372 ( .A(KEYINPUT10), .B(KEYINPUT82), .ZN(n313) );
  XNOR2_X1 U373 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U374 ( .A(n316), .B(n315), .Z(n321) );
  XOR2_X1 U375 ( .A(KEYINPUT83), .B(KEYINPUT65), .Z(n318) );
  NAND2_X1 U376 ( .A1(G232GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U377 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U378 ( .A(KEYINPUT11), .B(n319), .ZN(n320) );
  XNOR2_X1 U379 ( .A(n321), .B(n320), .ZN(n326) );
  XOR2_X1 U380 ( .A(KEYINPUT71), .B(KEYINPUT7), .Z(n323) );
  XNOR2_X1 U381 ( .A(G43GAT), .B(G29GAT), .ZN(n322) );
  XNOR2_X1 U382 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U383 ( .A(KEYINPUT8), .B(n324), .ZN(n440) );
  INV_X1 U384 ( .A(n440), .ZN(n325) );
  XOR2_X1 U385 ( .A(n326), .B(n325), .Z(n330) );
  XNOR2_X1 U386 ( .A(G50GAT), .B(KEYINPUT81), .ZN(n327) );
  XNOR2_X1 U387 ( .A(n327), .B(G162GAT), .ZN(n377) );
  XOR2_X1 U388 ( .A(G99GAT), .B(G85GAT), .Z(n446) );
  XNOR2_X1 U389 ( .A(n377), .B(n446), .ZN(n328) );
  XOR2_X1 U390 ( .A(G36GAT), .B(G190GAT), .Z(n364) );
  XOR2_X1 U391 ( .A(n328), .B(n364), .Z(n329) );
  XOR2_X1 U392 ( .A(n330), .B(n329), .Z(n485) );
  INV_X1 U393 ( .A(n485), .ZN(n565) );
  XOR2_X1 U394 ( .A(KEYINPUT36), .B(n565), .Z(n589) );
  XOR2_X1 U395 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n389) );
  XOR2_X1 U396 ( .A(KEYINPUT90), .B(G183GAT), .Z(n332) );
  XNOR2_X1 U397 ( .A(G190GAT), .B(G71GAT), .ZN(n331) );
  XNOR2_X1 U398 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U399 ( .A(n333), .B(G99GAT), .Z(n336) );
  XNOR2_X1 U400 ( .A(G43GAT), .B(n334), .ZN(n335) );
  XNOR2_X1 U401 ( .A(n336), .B(n335), .ZN(n341) );
  XNOR2_X1 U402 ( .A(G134GAT), .B(G120GAT), .ZN(n337) );
  XNOR2_X1 U403 ( .A(n337), .B(KEYINPUT0), .ZN(n407) );
  XOR2_X1 U404 ( .A(G113GAT), .B(n407), .Z(n339) );
  NAND2_X1 U405 ( .A1(G227GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U406 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U407 ( .A(n341), .B(n340), .Z(n351) );
  XNOR2_X1 U408 ( .A(KEYINPUT88), .B(KEYINPUT89), .ZN(n342) );
  XNOR2_X1 U409 ( .A(n342), .B(KEYINPUT18), .ZN(n344) );
  INV_X1 U410 ( .A(KEYINPUT17), .ZN(n343) );
  XNOR2_X1 U411 ( .A(n344), .B(n343), .ZN(n346) );
  XNOR2_X1 U412 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n345) );
  XNOR2_X1 U413 ( .A(n346), .B(n345), .ZN(n358) );
  XOR2_X1 U414 ( .A(G176GAT), .B(KEYINPUT87), .Z(n348) );
  XNOR2_X1 U415 ( .A(KEYINPUT20), .B(KEYINPUT66), .ZN(n347) );
  XNOR2_X1 U416 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U417 ( .A(n358), .B(n349), .ZN(n350) );
  XNOR2_X1 U418 ( .A(n351), .B(n350), .ZN(n536) );
  XOR2_X1 U419 ( .A(KEYINPUT99), .B(KEYINPUT98), .Z(n353) );
  NAND2_X1 U420 ( .A1(G226GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U421 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U422 ( .A(n354), .B(G204GAT), .Z(n360) );
  XOR2_X1 U423 ( .A(KEYINPUT92), .B(G218GAT), .Z(n356) );
  XNOR2_X1 U424 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n355) );
  XNOR2_X1 U425 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U426 ( .A(G197GAT), .B(n357), .Z(n379) );
  XNOR2_X1 U427 ( .A(n358), .B(n379), .ZN(n359) );
  XOR2_X1 U428 ( .A(n360), .B(n359), .Z(n362) );
  XNOR2_X1 U429 ( .A(n362), .B(n361), .ZN(n366) );
  XNOR2_X1 U430 ( .A(G176GAT), .B(G92GAT), .ZN(n363) );
  XNOR2_X1 U431 ( .A(n363), .B(G64GAT), .ZN(n453) );
  XNOR2_X1 U432 ( .A(n453), .B(n364), .ZN(n365) );
  XNOR2_X1 U433 ( .A(n366), .B(n365), .ZN(n465) );
  NAND2_X1 U434 ( .A1(n536), .A2(n465), .ZN(n367) );
  XOR2_X1 U435 ( .A(KEYINPUT101), .B(n367), .Z(n387) );
  XOR2_X1 U436 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n369) );
  XNOR2_X1 U437 ( .A(KEYINPUT24), .B(KEYINPUT94), .ZN(n368) );
  XNOR2_X1 U438 ( .A(n369), .B(n368), .ZN(n373) );
  NAND2_X1 U439 ( .A1(G228GAT), .A2(G233GAT), .ZN(n371) );
  XOR2_X1 U440 ( .A(G155GAT), .B(KEYINPUT2), .Z(n375) );
  XNOR2_X1 U441 ( .A(KEYINPUT3), .B(KEYINPUT93), .ZN(n374) );
  XNOR2_X1 U442 ( .A(n375), .B(n374), .ZN(n403) );
  XOR2_X1 U443 ( .A(n376), .B(n403), .Z(n381) );
  XOR2_X1 U444 ( .A(G141GAT), .B(G22GAT), .Z(n425) );
  XNOR2_X1 U445 ( .A(n425), .B(n377), .ZN(n378) );
  XOR2_X1 U446 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n383) );
  XNOR2_X1 U447 ( .A(G78GAT), .B(G148GAT), .ZN(n382) );
  XNOR2_X1 U448 ( .A(n383), .B(n382), .ZN(n385) );
  XOR2_X1 U449 ( .A(G106GAT), .B(G204GAT), .Z(n384) );
  XNOR2_X1 U450 ( .A(n385), .B(n384), .ZN(n458) );
  XNOR2_X1 U451 ( .A(n386), .B(n458), .ZN(n416) );
  NAND2_X1 U452 ( .A1(n387), .A2(n416), .ZN(n388) );
  XNOR2_X1 U453 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U454 ( .A(KEYINPUT25), .B(n390), .ZN(n394) );
  XOR2_X1 U455 ( .A(n465), .B(KEYINPUT27), .Z(n417) );
  NOR2_X1 U456 ( .A1(n536), .A2(n416), .ZN(n391) );
  XNOR2_X1 U457 ( .A(KEYINPUT26), .B(n391), .ZN(n574) );
  INV_X1 U458 ( .A(n574), .ZN(n392) );
  XNOR2_X1 U459 ( .A(n552), .B(KEYINPUT100), .ZN(n393) );
  NOR2_X1 U460 ( .A1(n394), .A2(n393), .ZN(n414) );
  XOR2_X1 U461 ( .A(KEYINPUT97), .B(KEYINPUT6), .Z(n396) );
  XNOR2_X1 U462 ( .A(KEYINPUT5), .B(KEYINPUT95), .ZN(n395) );
  XNOR2_X1 U463 ( .A(n396), .B(n395), .ZN(n413) );
  XOR2_X1 U464 ( .A(KEYINPUT1), .B(G57GAT), .Z(n398) );
  XNOR2_X1 U465 ( .A(G141GAT), .B(G148GAT), .ZN(n397) );
  XNOR2_X1 U466 ( .A(n398), .B(n397), .ZN(n402) );
  XOR2_X1 U467 ( .A(G85GAT), .B(G162GAT), .Z(n400) );
  XNOR2_X1 U468 ( .A(G29GAT), .B(G127GAT), .ZN(n399) );
  XNOR2_X1 U469 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U470 ( .A(n402), .B(n401), .ZN(n411) );
  XOR2_X1 U471 ( .A(G113GAT), .B(G1GAT), .Z(n424) );
  XOR2_X1 U472 ( .A(n424), .B(n403), .Z(n405) );
  NAND2_X1 U473 ( .A1(G225GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U474 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U475 ( .A(n406), .B(KEYINPUT4), .Z(n409) );
  XNOR2_X1 U476 ( .A(n407), .B(KEYINPUT96), .ZN(n408) );
  XNOR2_X1 U477 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U478 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U479 ( .A(n413), .B(n412), .Z(n553) );
  INV_X1 U480 ( .A(n553), .ZN(n524) );
  XNOR2_X1 U481 ( .A(n415), .B(KEYINPUT104), .ZN(n420) );
  XOR2_X1 U482 ( .A(KEYINPUT28), .B(n416), .Z(n533) );
  NOR2_X1 U483 ( .A1(n417), .A2(n533), .ZN(n418) );
  NAND2_X1 U484 ( .A1(n418), .A2(n524), .ZN(n538) );
  NOR2_X1 U485 ( .A1(n538), .A2(n536), .ZN(n419) );
  NOR2_X1 U486 ( .A1(n589), .A2(n495), .ZN(n422) );
  NAND2_X1 U487 ( .A1(n572), .A2(n422), .ZN(n423) );
  XNOR2_X1 U488 ( .A(KEYINPUT37), .B(n423), .ZN(n523) );
  XOR2_X1 U489 ( .A(G36GAT), .B(G50GAT), .Z(n427) );
  XNOR2_X1 U490 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U491 ( .A(n427), .B(n426), .ZN(n432) );
  XOR2_X1 U492 ( .A(KEYINPUT69), .B(G8GAT), .Z(n429) );
  XNOR2_X1 U493 ( .A(KEYINPUT29), .B(KEYINPUT72), .ZN(n428) );
  XNOR2_X1 U494 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U495 ( .A(KEYINPUT73), .B(G197GAT), .Z(n434) );
  XNOR2_X1 U496 ( .A(G169GAT), .B(G15GAT), .ZN(n433) );
  XOR2_X1 U497 ( .A(n434), .B(n433), .Z(n435) );
  XNOR2_X1 U498 ( .A(n436), .B(n435), .ZN(n442) );
  XOR2_X1 U499 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n438) );
  XNOR2_X1 U500 ( .A(KEYINPUT67), .B(KEYINPUT70), .ZN(n437) );
  XNOR2_X1 U501 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U502 ( .A(n440), .B(n439), .Z(n441) );
  INV_X1 U503 ( .A(n576), .ZN(n569) );
  XOR2_X1 U504 ( .A(KEYINPUT79), .B(KEYINPUT75), .Z(n444) );
  XNOR2_X1 U505 ( .A(KEYINPUT78), .B(KEYINPUT31), .ZN(n443) );
  XNOR2_X1 U506 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U507 ( .A(n445), .B(KEYINPUT33), .Z(n448) );
  XNOR2_X1 U508 ( .A(G120GAT), .B(n446), .ZN(n447) );
  XNOR2_X1 U509 ( .A(n448), .B(n447), .ZN(n457) );
  XOR2_X1 U510 ( .A(KEYINPUT74), .B(KEYINPUT32), .Z(n450) );
  NAND2_X1 U511 ( .A1(G230GAT), .A2(G233GAT), .ZN(n449) );
  XNOR2_X1 U512 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U513 ( .A(n451), .B(KEYINPUT80), .Z(n455) );
  XNOR2_X1 U514 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U515 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U516 ( .A(n457), .B(n456), .ZN(n459) );
  XNOR2_X1 U517 ( .A(n459), .B(n458), .ZN(n581) );
  NOR2_X1 U518 ( .A1(n569), .A2(n581), .ZN(n496) );
  NAND2_X1 U519 ( .A1(n523), .A2(n496), .ZN(n460) );
  NAND2_X1 U520 ( .A1(n509), .A2(n524), .ZN(n464) );
  XOR2_X1 U521 ( .A(KEYINPUT39), .B(KEYINPUT108), .Z(n462) );
  XOR2_X1 U522 ( .A(KEYINPUT54), .B(KEYINPUT123), .Z(n479) );
  BUF_X1 U523 ( .A(n465), .Z(n527) );
  XNOR2_X1 U524 ( .A(KEYINPUT41), .B(n581), .ZN(n560) );
  NOR2_X1 U525 ( .A1(n569), .A2(n560), .ZN(n466) );
  XNOR2_X1 U526 ( .A(n466), .B(KEYINPUT46), .ZN(n467) );
  NOR2_X1 U527 ( .A1(n565), .A2(n467), .ZN(n468) );
  NAND2_X1 U528 ( .A1(n468), .A2(n572), .ZN(n469) );
  XNOR2_X1 U529 ( .A(n469), .B(KEYINPUT47), .ZN(n474) );
  NOR2_X1 U530 ( .A1(n589), .A2(n572), .ZN(n470) );
  XNOR2_X1 U531 ( .A(KEYINPUT45), .B(n470), .ZN(n471) );
  NAND2_X1 U532 ( .A1(n471), .A2(n569), .ZN(n472) );
  NOR2_X1 U533 ( .A1(n581), .A2(n472), .ZN(n473) );
  NOR2_X1 U534 ( .A1(n474), .A2(n473), .ZN(n477) );
  INV_X1 U535 ( .A(KEYINPUT116), .ZN(n475) );
  NAND2_X1 U536 ( .A1(n527), .A2(n551), .ZN(n478) );
  XNOR2_X1 U537 ( .A(n479), .B(n478), .ZN(n480) );
  NOR2_X1 U538 ( .A1(n524), .A2(n480), .ZN(n481) );
  XNOR2_X1 U539 ( .A(n481), .B(KEYINPUT64), .ZN(n575) );
  NAND2_X1 U540 ( .A1(n416), .A2(n575), .ZN(n483) );
  INV_X1 U541 ( .A(KEYINPUT55), .ZN(n482) );
  XOR2_X1 U542 ( .A(n483), .B(n482), .Z(n484) );
  NAND2_X1 U543 ( .A1(n484), .A2(n536), .ZN(n571) );
  NOR2_X1 U544 ( .A1(n485), .A2(n571), .ZN(n488) );
  INV_X1 U545 ( .A(G190GAT), .ZN(n486) );
  XOR2_X1 U546 ( .A(n560), .B(KEYINPUT109), .Z(n542) );
  NOR2_X1 U547 ( .A1(n542), .A2(n571), .ZN(n491) );
  XNOR2_X1 U548 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n489) );
  XNOR2_X1 U549 ( .A(n489), .B(G176GAT), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n491), .B(n490), .ZN(G1349GAT) );
  XOR2_X1 U551 ( .A(KEYINPUT107), .B(KEYINPUT34), .Z(n499) );
  NOR2_X1 U552 ( .A1(n565), .A2(n572), .ZN(n492) );
  XOR2_X1 U553 ( .A(KEYINPUT16), .B(n492), .Z(n493) );
  XNOR2_X1 U554 ( .A(n493), .B(KEYINPUT86), .ZN(n494) );
  NOR2_X1 U555 ( .A1(n495), .A2(n494), .ZN(n511) );
  NAND2_X1 U556 ( .A1(n511), .A2(n496), .ZN(n497) );
  XOR2_X1 U557 ( .A(KEYINPUT106), .B(n497), .Z(n504) );
  NAND2_X1 U558 ( .A1(n504), .A2(n524), .ZN(n498) );
  XNOR2_X1 U559 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U560 ( .A(G1GAT), .B(n500), .ZN(G1324GAT) );
  NAND2_X1 U561 ( .A1(n504), .A2(n527), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n501), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U563 ( .A(G15GAT), .B(KEYINPUT35), .Z(n503) );
  NAND2_X1 U564 ( .A1(n536), .A2(n504), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n503), .B(n502), .ZN(G1326GAT) );
  NAND2_X1 U566 ( .A1(n504), .A2(n533), .ZN(n505) );
  XNOR2_X1 U567 ( .A(n505), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U568 ( .A1(n509), .A2(n527), .ZN(n506) );
  XNOR2_X1 U569 ( .A(n506), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U570 ( .A1(n509), .A2(n536), .ZN(n507) );
  XNOR2_X1 U571 ( .A(n507), .B(KEYINPUT40), .ZN(n508) );
  XNOR2_X1 U572 ( .A(G43GAT), .B(n508), .ZN(G1330GAT) );
  NAND2_X1 U573 ( .A1(n509), .A2(n533), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n510), .B(G50GAT), .ZN(G1331GAT) );
  NOR2_X1 U575 ( .A1(n542), .A2(n576), .ZN(n522) );
  AND2_X1 U576 ( .A1(n511), .A2(n522), .ZN(n519) );
  NAND2_X1 U577 ( .A1(n519), .A2(n524), .ZN(n512) );
  XNOR2_X1 U578 ( .A(KEYINPUT42), .B(n512), .ZN(n513) );
  XNOR2_X1 U579 ( .A(G57GAT), .B(n513), .ZN(G1332GAT) );
  NAND2_X1 U580 ( .A1(n519), .A2(n527), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n514), .B(KEYINPUT110), .ZN(n515) );
  XNOR2_X1 U582 ( .A(G64GAT), .B(n515), .ZN(G1333GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n517) );
  NAND2_X1 U584 ( .A1(n519), .A2(n536), .ZN(n516) );
  XNOR2_X1 U585 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U586 ( .A(G71GAT), .B(n518), .ZN(G1334GAT) );
  XOR2_X1 U587 ( .A(G78GAT), .B(KEYINPUT43), .Z(n521) );
  NAND2_X1 U588 ( .A1(n519), .A2(n533), .ZN(n520) );
  XNOR2_X1 U589 ( .A(n521), .B(n520), .ZN(G1335GAT) );
  XOR2_X1 U590 ( .A(G85GAT), .B(KEYINPUT113), .Z(n526) );
  AND2_X1 U591 ( .A1(n523), .A2(n522), .ZN(n532) );
  NAND2_X1 U592 ( .A1(n532), .A2(n524), .ZN(n525) );
  XNOR2_X1 U593 ( .A(n526), .B(n525), .ZN(G1336GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n529) );
  NAND2_X1 U595 ( .A1(n532), .A2(n527), .ZN(n528) );
  XNOR2_X1 U596 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U597 ( .A(G92GAT), .B(n530), .ZN(G1337GAT) );
  NAND2_X1 U598 ( .A1(n532), .A2(n536), .ZN(n531) );
  XNOR2_X1 U599 ( .A(n531), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U600 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n534), .B(KEYINPUT44), .ZN(n535) );
  XNOR2_X1 U602 ( .A(G106GAT), .B(n535), .ZN(G1339GAT) );
  XOR2_X1 U603 ( .A(G113GAT), .B(KEYINPUT117), .Z(n540) );
  NAND2_X1 U604 ( .A1(n536), .A2(n551), .ZN(n537) );
  NOR2_X1 U605 ( .A1(n538), .A2(n537), .ZN(n548) );
  NAND2_X1 U606 ( .A1(n548), .A2(n576), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(G1340GAT) );
  INV_X1 U608 ( .A(n548), .ZN(n541) );
  NOR2_X1 U609 ( .A1(n542), .A2(n541), .ZN(n544) );
  XNOR2_X1 U610 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(G1341GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n546) );
  NAND2_X1 U613 ( .A1(n548), .A2(n586), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U615 ( .A(G127GAT), .B(n547), .Z(G1342GAT) );
  XOR2_X1 U616 ( .A(G134GAT), .B(KEYINPUT51), .Z(n550) );
  NAND2_X1 U617 ( .A1(n548), .A2(n565), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  NAND2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n554) );
  NOR2_X1 U620 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U621 ( .A(KEYINPUT119), .B(n555), .ZN(n559) );
  INV_X1 U622 ( .A(n559), .ZN(n566) );
  NAND2_X1 U623 ( .A1(n566), .A2(n576), .ZN(n556) );
  XNOR2_X1 U624 ( .A(G141GAT), .B(n556), .ZN(G1344GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT120), .B(KEYINPUT52), .Z(n558) );
  XNOR2_X1 U626 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n557) );
  XNOR2_X1 U627 ( .A(n558), .B(n557), .ZN(n562) );
  NOR2_X1 U628 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U629 ( .A(n562), .B(n561), .Z(G1345GAT) );
  XOR2_X1 U630 ( .A(G155GAT), .B(KEYINPUT121), .Z(n564) );
  NAND2_X1 U631 ( .A1(n566), .A2(n586), .ZN(n563) );
  XNOR2_X1 U632 ( .A(n564), .B(n563), .ZN(G1346GAT) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(KEYINPUT122), .ZN(n568) );
  XNOR2_X1 U635 ( .A(G162GAT), .B(n568), .ZN(G1347GAT) );
  NOR2_X1 U636 ( .A1(n569), .A2(n571), .ZN(n570) );
  XOR2_X1 U637 ( .A(G169GAT), .B(n570), .Z(G1348GAT) );
  NOR2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U639 ( .A(G183GAT), .B(n573), .Z(G1350GAT) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n588) );
  INV_X1 U641 ( .A(n588), .ZN(n585) );
  NAND2_X1 U642 ( .A1(n576), .A2(n585), .ZN(n580) );
  XOR2_X1 U643 ( .A(KEYINPUT124), .B(KEYINPUT59), .Z(n578) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n577) );
  XNOR2_X1 U645 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n583) );
  NAND2_X1 U648 ( .A1(n585), .A2(n581), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(n584) );
  XOR2_X1 U650 ( .A(G204GAT), .B(n584), .Z(G1353GAT) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n587), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n591) );
  XNOR2_X1 U654 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n591), .B(n590), .ZN(n592) );
  XOR2_X1 U656 ( .A(G218GAT), .B(n592), .Z(G1355GAT) );
endmodule

