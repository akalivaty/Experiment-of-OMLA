//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 0 0 1 0 1 1 0 1 1 0 1 0 0 0 1 0 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n753, new_n754, new_n755, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028;
  INV_X1    g000(.A(KEYINPUT29), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT65), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT11), .ZN(new_n189));
  INV_X1    g003(.A(G137), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n189), .B1(G134), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G134), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT64), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G134), .ZN(new_n195));
  AOI21_X1  g009(.A(G137), .B1(new_n193), .B2(new_n195), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n191), .B1(new_n196), .B2(new_n189), .ZN(new_n197));
  INV_X1    g011(.A(G131), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n193), .A2(new_n195), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(new_n190), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n188), .B1(new_n197), .B2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT64), .B(G134), .ZN(new_n202));
  AOI21_X1  g016(.A(G131), .B1(new_n202), .B2(G137), .ZN(new_n203));
  NOR3_X1   g017(.A1(new_n202), .A2(KEYINPUT11), .A3(G137), .ZN(new_n204));
  OAI211_X1 g018(.A(KEYINPUT65), .B(new_n203), .C1(new_n204), .C2(new_n191), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n201), .A2(new_n205), .ZN(new_n206));
  OAI22_X1  g020(.A1(new_n204), .A2(new_n191), .B1(new_n190), .B2(new_n199), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G131), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT0), .A2(G128), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  XOR2_X1   g031(.A(KEYINPUT0), .B(G128), .Z(new_n218));
  OAI21_X1  g032(.A(new_n217), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n209), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n211), .A2(new_n213), .A3(G128), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n223), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(new_n212), .A3(G146), .ZN(new_n226));
  AOI21_X1  g040(.A(G128), .B1(new_n211), .B2(new_n213), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n224), .A2(new_n226), .A3(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n190), .A2(G134), .ZN(new_n230));
  OAI21_X1  g044(.A(G131), .B1(new_n196), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT66), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI211_X1 g047(.A(KEYINPUT66), .B(G131), .C1(new_n196), .C2(new_n230), .ZN(new_n234));
  AOI22_X1  g048(.A1(new_n201), .A2(new_n205), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n229), .B1(new_n235), .B2(KEYINPUT67), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n233), .A2(new_n234), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n206), .A2(KEYINPUT67), .A3(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n220), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT74), .ZN(new_n240));
  XNOR2_X1  g054(.A(G116), .B(G119), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT2), .B(G113), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n243), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n241), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n244), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n242), .A2(KEYINPUT70), .A3(new_n243), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n239), .A2(new_n240), .A3(new_n251), .ZN(new_n252));
  NOR3_X1   g066(.A1(new_n197), .A2(new_n188), .A3(new_n200), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n194), .A2(G134), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n192), .A2(KEYINPUT64), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n189), .B(new_n190), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n191), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(KEYINPUT65), .B1(new_n258), .B2(new_n203), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n237), .B1(new_n253), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n235), .A2(KEYINPUT67), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(new_n229), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n250), .B1(new_n264), .B2(new_n220), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n235), .A2(new_n229), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n220), .A2(new_n266), .A3(new_n250), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT74), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n252), .B(KEYINPUT28), .C1(new_n265), .C2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n267), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n270), .A2(KEYINPUT28), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G237), .ZN(new_n273));
  INV_X1    g087(.A(G953), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n273), .A2(new_n274), .A3(G210), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n275), .B(KEYINPUT27), .ZN(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT26), .B(G101), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n276), .B(new_n277), .ZN(new_n278));
  XOR2_X1   g092(.A(new_n278), .B(KEYINPUT73), .Z(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n269), .A2(new_n272), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT69), .ZN(new_n282));
  OR2_X1    g096(.A1(new_n215), .A2(new_n218), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n206), .A2(new_n208), .B1(new_n283), .B2(new_n217), .ZN(new_n284));
  INV_X1    g098(.A(new_n229), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n285), .B1(new_n260), .B2(new_n261), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n284), .B1(new_n286), .B2(new_n263), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n282), .B1(new_n287), .B2(KEYINPUT30), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT30), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n239), .A2(KEYINPUT69), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n220), .A2(KEYINPUT30), .A3(new_n266), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n251), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n270), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n187), .B(new_n281), .C1(new_n295), .C2(new_n278), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n220), .A2(new_n266), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n297), .B(new_n251), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n271), .B1(new_n298), .B2(KEYINPUT28), .ZN(new_n299));
  INV_X1    g113(.A(new_n278), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n300), .A2(new_n187), .ZN(new_n301));
  AOI21_X1  g115(.A(G902), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n296), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G472), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n269), .A2(new_n272), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n279), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n293), .B1(new_n288), .B2(new_n290), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT71), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n267), .A2(new_n308), .A3(new_n278), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n308), .B1(new_n267), .B2(new_n278), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(KEYINPUT31), .B1(new_n307), .B2(new_n311), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n287), .A2(new_n282), .A3(KEYINPUT30), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT69), .B1(new_n239), .B2(new_n289), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n294), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  OR2_X1    g129(.A1(new_n309), .A2(new_n310), .ZN(new_n316));
  XOR2_X1   g130(.A(KEYINPUT72), .B(KEYINPUT31), .Z(new_n317));
  NAND3_X1  g131(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n306), .A2(new_n312), .A3(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT32), .ZN(new_n320));
  NOR2_X1   g134(.A1(G472), .A2(G902), .ZN(new_n321));
  AND3_X1   g135(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n320), .B1(new_n319), .B2(new_n321), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n304), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT75), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n326), .B(new_n304), .C1(new_n322), .C2(new_n323), .ZN(new_n327));
  INV_X1    g141(.A(G217), .ZN(new_n328));
  INV_X1    g142(.A(G902), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n328), .B1(G234), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT80), .ZN(new_n331));
  XNOR2_X1  g145(.A(G125), .B(G140), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n210), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT79), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT79), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n332), .A2(new_n335), .A3(new_n210), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n332), .A2(KEYINPUT16), .ZN(new_n338));
  INV_X1    g152(.A(G125), .ZN(new_n339));
  OR3_X1    g153(.A1(new_n339), .A2(KEYINPUT16), .A3(G140), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(G146), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT78), .ZN(new_n343));
  INV_X1    g157(.A(G128), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G119), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n344), .A2(G119), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT23), .ZN(new_n347));
  OAI211_X1 g161(.A(KEYINPUT77), .B(new_n345), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G119), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G128), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n349), .A2(G128), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT77), .ZN(new_n352));
  OAI211_X1 g166(.A(KEYINPUT23), .B(new_n350), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G110), .ZN(new_n354));
  AND3_X1   g168(.A1(new_n348), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(KEYINPUT24), .B(G110), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT76), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n358), .B1(new_n346), .B2(new_n351), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n350), .A2(new_n345), .A3(KEYINPUT76), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n357), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n343), .B1(new_n355), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n360), .ZN(new_n363));
  AOI21_X1  g177(.A(KEYINPUT76), .B1(new_n350), .B2(new_n345), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n356), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n348), .A2(new_n353), .A3(new_n354), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(KEYINPUT78), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n342), .B1(new_n362), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n348), .A2(new_n353), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G110), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n359), .A2(new_n360), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n370), .B1(new_n371), .B2(new_n356), .ZN(new_n372));
  INV_X1    g186(.A(new_n341), .ZN(new_n373));
  AOI21_X1  g187(.A(G146), .B1(new_n338), .B2(new_n340), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n331), .B1(new_n368), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n342), .ZN(new_n378));
  NOR3_X1   g192(.A1(new_n355), .A2(new_n361), .A3(new_n343), .ZN(new_n379));
  AOI21_X1  g193(.A(KEYINPUT78), .B1(new_n365), .B2(new_n366), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OAI221_X1 g195(.A(new_n370), .B1(new_n371), .B2(new_n356), .C1(new_n373), .C2(new_n374), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(KEYINPUT80), .A3(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(KEYINPUT22), .B(G137), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n274), .A2(G221), .A3(G234), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n384), .B(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n377), .A2(new_n383), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n381), .A2(new_n382), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(new_n331), .A3(new_n386), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(KEYINPUT25), .B1(new_n391), .B2(new_n329), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT25), .ZN(new_n393));
  AOI211_X1 g207(.A(new_n393), .B(G902), .C1(new_n388), .C2(new_n390), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n330), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT81), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI211_X1 g211(.A(KEYINPUT81), .B(new_n330), .C1(new_n392), .C2(new_n394), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n330), .A2(G902), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n391), .A2(new_n399), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n397), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n325), .A2(new_n327), .A3(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(KEYINPUT9), .B(G234), .ZN(new_n403));
  OAI21_X1  g217(.A(G221), .B1(new_n403), .B2(G902), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n404), .B(KEYINPUT82), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(G214), .B1(G237), .B2(G902), .ZN(new_n407));
  INV_X1    g221(.A(G104), .ZN(new_n408));
  OAI21_X1  g222(.A(KEYINPUT3), .B1(new_n408), .B2(G107), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT3), .ZN(new_n410));
  INV_X1    g224(.A(G107), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n411), .A3(G104), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n408), .A2(G107), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n409), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT4), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(new_n415), .A3(G101), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n414), .A2(G101), .ZN(new_n417));
  INV_X1    g231(.A(G101), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n409), .A2(new_n412), .A3(new_n418), .A4(new_n413), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT4), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n416), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  OR2_X1    g235(.A1(new_n250), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n408), .A2(G107), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n411), .A2(G104), .ZN(new_n424));
  OAI21_X1  g238(.A(G101), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n419), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT5), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(new_n349), .A3(G116), .ZN(new_n429));
  OAI211_X1 g243(.A(G113), .B(new_n429), .C1(new_n242), .C2(new_n428), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n427), .A2(new_n246), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n422), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(G110), .B(G122), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n422), .A2(new_n433), .A3(new_n431), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(KEYINPUT6), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n229), .A2(new_n339), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n219), .A2(G125), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n274), .A2(G224), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n440), .B(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT6), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n432), .A2(new_n443), .A3(new_n434), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n437), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(G210), .B1(G237), .B2(G902), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT89), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT7), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n440), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n441), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n451), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n427), .B1(new_n246), .B2(new_n430), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT88), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n433), .B(KEYINPUT8), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT88), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n431), .A2(new_n457), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n455), .B(new_n456), .C1(new_n458), .C2(new_n454), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n440), .A2(new_n449), .A3(KEYINPUT7), .A4(new_n441), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n453), .A2(new_n459), .A3(new_n436), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n329), .ZN(new_n462));
  NOR3_X1   g276(.A1(new_n446), .A2(new_n448), .A3(new_n462), .ZN(new_n463));
  XOR2_X1   g277(.A(new_n447), .B(KEYINPUT90), .Z(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n461), .A2(new_n329), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n465), .B1(new_n466), .B2(new_n445), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n407), .B1(new_n463), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(KEYINPUT92), .B1(new_n344), .B2(G143), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT92), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(new_n212), .A3(G128), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n344), .A2(G143), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n202), .A3(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n202), .B1(new_n472), .B2(new_n473), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(G122), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G116), .ZN(new_n479));
  INV_X1    g293(.A(G116), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(G122), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n411), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n479), .A2(new_n481), .A3(G107), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n479), .A2(KEYINPUT14), .A3(G107), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n479), .A2(new_n481), .A3(KEYINPUT14), .A4(G107), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(KEYINPUT93), .B1(new_n477), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n472), .A2(new_n473), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n199), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n474), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT93), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n492), .A2(new_n493), .A3(new_n486), .A4(new_n487), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT13), .ZN(new_n496));
  AOI22_X1  g310(.A1(new_n472), .A2(new_n496), .B1(new_n344), .B2(G143), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n497), .B1(new_n496), .B2(new_n472), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G134), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n499), .A2(new_n474), .A3(new_n483), .A4(new_n484), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  NOR3_X1   g315(.A1(new_n403), .A2(new_n328), .A3(G953), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n495), .A2(new_n500), .A3(new_n502), .ZN(new_n505));
  AOI21_X1  g319(.A(G902), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G478), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n507), .A2(KEYINPUT15), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n506), .A2(new_n509), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n273), .A2(new_n274), .A3(G214), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(G143), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT91), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT18), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n516), .B1(new_n517), .B2(new_n198), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n515), .A2(KEYINPUT91), .A3(KEYINPUT18), .A4(G131), .ZN(new_n519));
  OR2_X1    g333(.A1(new_n332), .A2(new_n210), .ZN(new_n520));
  AOI22_X1  g334(.A1(new_n518), .A2(new_n519), .B1(new_n337), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n515), .A2(new_n198), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT17), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n515), .B(new_n198), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n375), .B(new_n524), .C1(new_n525), .C2(KEYINPUT17), .ZN(new_n526));
  XNOR2_X1  g340(.A(G113), .B(G122), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(new_n408), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n522), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n528), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n332), .B(KEYINPUT19), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n373), .B1(new_n210), .B2(new_n531), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n532), .A2(new_n525), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n530), .B1(new_n533), .B2(new_n521), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n529), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(G475), .A2(G902), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(KEYINPUT20), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT20), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n535), .A2(new_n539), .A3(new_n536), .ZN(new_n540));
  INV_X1    g354(.A(new_n529), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n528), .B1(new_n522), .B2(new_n526), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n329), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI22_X1  g357(.A1(new_n538), .A2(new_n540), .B1(G475), .B2(new_n543), .ZN(new_n544));
  AND2_X1   g358(.A1(new_n274), .A2(G952), .ZN(new_n545));
  NAND2_X1  g359(.A1(G234), .A2(G237), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  XOR2_X1   g361(.A(new_n547), .B(KEYINPUT94), .Z(new_n548));
  XNOR2_X1  g362(.A(KEYINPUT21), .B(G898), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n546), .A2(G902), .A3(G953), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n548), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  XOR2_X1   g366(.A(new_n552), .B(KEYINPUT95), .Z(new_n553));
  NAND3_X1  g367(.A1(new_n513), .A2(new_n544), .A3(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n468), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(G110), .B(G140), .ZN(new_n556));
  INV_X1    g370(.A(G227), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n557), .A2(G953), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n556), .B(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n212), .A2(KEYINPUT1), .A3(G146), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n228), .B(new_n561), .C1(new_n225), .C2(new_n221), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n427), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n426), .A2(new_n224), .A3(new_n226), .A4(new_n228), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n209), .A2(KEYINPUT12), .A3(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT83), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT12), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n563), .A2(new_n564), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n201), .A2(new_n205), .B1(new_n207), .B2(G131), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n209), .A2(KEYINPUT83), .A3(KEYINPUT12), .A4(new_n565), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n568), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n219), .B(new_n416), .C1(new_n417), .C2(new_n420), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT10), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n563), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n229), .A2(KEYINPUT10), .A3(new_n427), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n571), .A2(new_n575), .A3(new_n577), .A4(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n560), .B1(new_n574), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(KEYINPUT84), .A3(new_n560), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n577), .A2(new_n575), .A3(new_n578), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n209), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT84), .B1(new_n579), .B2(new_n560), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(KEYINPUT85), .B1(new_n580), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n585), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n588), .A2(new_n583), .A3(new_n581), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT85), .ZN(new_n590));
  INV_X1    g404(.A(new_n579), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n572), .A2(new_n573), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n591), .B1(new_n592), .B2(new_n568), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n589), .B(new_n590), .C1(new_n593), .C2(new_n560), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n587), .A2(new_n594), .A3(new_n329), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT86), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n595), .A2(new_n596), .A3(G469), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n572), .A2(new_n573), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n206), .A2(new_n208), .B1(new_n563), .B2(new_n564), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT83), .B1(new_n599), .B2(KEYINPUT12), .ZN(new_n600));
  OAI21_X1  g414(.A(KEYINPUT87), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT87), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n568), .A2(new_n602), .A3(new_n572), .A4(new_n573), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n601), .A2(new_n579), .A3(new_n560), .A4(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n560), .B1(new_n583), .B2(new_n579), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(G469), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n607), .A2(new_n608), .A3(new_n329), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n597), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n596), .B1(new_n595), .B2(G469), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n406), .B(new_n555), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT96), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n595), .A2(G469), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(KEYINPUT86), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n616), .A2(new_n597), .A3(new_n609), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n617), .A2(KEYINPUT96), .A3(new_n406), .A4(new_n555), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n402), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(new_n418), .ZN(G3));
  INV_X1    g435(.A(G472), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n319), .B2(new_n329), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT97), .ZN(new_n624));
  OR2_X1    g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI22_X1  g439(.A1(new_n623), .A2(new_n624), .B1(new_n321), .B2(new_n319), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n617), .A2(new_n401), .A3(new_n406), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n507), .A2(new_n329), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n630), .B1(new_n506), .B2(new_n507), .ZN(new_n631));
  INV_X1    g445(.A(new_n505), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n502), .B1(new_n495), .B2(new_n500), .ZN(new_n633));
  OAI21_X1  g447(.A(KEYINPUT33), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT33), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n504), .A2(new_n635), .A3(new_n505), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n634), .A2(new_n636), .A3(G478), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n631), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(KEYINPUT98), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT98), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n631), .A2(new_n637), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n538), .A2(new_n540), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n543), .A2(G475), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n407), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n448), .B1(new_n446), .B2(new_n462), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n466), .A2(new_n447), .A3(new_n445), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n553), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n646), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n629), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT99), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT34), .B(G104), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G6));
  INV_X1    g471(.A(KEYINPUT101), .ZN(new_n658));
  XOR2_X1   g472(.A(new_n553), .B(KEYINPUT100), .Z(new_n659));
  OAI211_X1 g473(.A(new_n544), .B(new_n659), .C1(new_n512), .C2(new_n511), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n658), .B1(new_n651), .B2(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n645), .A2(new_n513), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n662), .A2(new_n650), .A3(KEYINPUT101), .A4(new_n659), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n629), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT35), .B(G107), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G9));
  NOR2_X1   g481(.A1(new_n387), .A2(KEYINPUT36), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n389), .B(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n399), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n397), .A2(new_n398), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT102), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n397), .A2(KEYINPUT102), .A3(new_n398), .A4(new_n670), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n675), .A2(new_n625), .A3(new_n626), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(KEYINPUT103), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n614), .A2(new_n618), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n675), .A2(new_n625), .A3(new_n626), .A4(new_n679), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n677), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT37), .B(G110), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT104), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n681), .B(new_n683), .ZN(G12));
  OAI21_X1  g498(.A(new_n406), .B1(new_n610), .B2(new_n611), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n673), .A2(new_n674), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n548), .B1(G900), .B2(new_n551), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n662), .A2(new_n687), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n685), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n689), .A2(new_n325), .A3(new_n327), .A4(new_n650), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G128), .ZN(G30));
  INV_X1    g505(.A(new_n685), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n687), .B(KEYINPUT39), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(KEYINPUT40), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT40), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n692), .A2(new_n696), .A3(new_n693), .ZN(new_n697));
  OR2_X1    g511(.A1(new_n322), .A2(new_n323), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n307), .A2(new_n311), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n699), .B1(new_n279), .B2(new_n298), .ZN(new_n700));
  OAI21_X1  g514(.A(G472), .B1(new_n700), .B2(G902), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n464), .B1(new_n446), .B2(new_n462), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n649), .ZN(new_n704));
  XOR2_X1   g518(.A(new_n704), .B(KEYINPUT38), .Z(new_n705));
  NOR2_X1   g519(.A1(new_n513), .A2(new_n544), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n407), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n705), .A2(new_n671), .A3(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n695), .A2(new_n697), .A3(new_n702), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G143), .ZN(G45));
  INV_X1    g524(.A(new_n641), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n640), .B1(new_n631), .B2(new_n637), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n645), .B(new_n687), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT105), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n642), .A2(KEYINPUT105), .A3(new_n645), .A4(new_n687), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n685), .A2(new_n686), .A3(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n718), .A2(new_n325), .A3(new_n327), .A4(new_n650), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G146), .ZN(G48));
  NAND2_X1  g534(.A1(new_n579), .A2(new_n560), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n721), .B1(new_n574), .B2(KEYINPUT87), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n605), .B1(new_n722), .B2(new_n603), .ZN(new_n723));
  OAI21_X1  g537(.A(G469), .B1(new_n723), .B2(G902), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n724), .A2(new_n609), .A3(new_n406), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT106), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n724), .A2(new_n609), .A3(KEYINPUT106), .A4(new_n406), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n729), .A2(new_n653), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n730), .A2(new_n325), .A3(new_n327), .A4(new_n401), .ZN(new_n731));
  XNOR2_X1  g545(.A(KEYINPUT41), .B(G113), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(KEYINPUT107), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n731), .B(new_n733), .ZN(G15));
  AND2_X1   g548(.A1(new_n729), .A2(new_n664), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n735), .A2(new_n325), .A3(new_n327), .A4(new_n401), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G116), .ZN(G18));
  INV_X1    g551(.A(new_n554), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n673), .A2(new_n738), .A3(new_n674), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n727), .A2(new_n650), .A3(new_n728), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n325), .A2(new_n741), .A3(new_n327), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G119), .ZN(G21));
  NAND2_X1  g557(.A1(new_n319), .A2(new_n329), .ZN(new_n744));
  XOR2_X1   g558(.A(KEYINPUT108), .B(G472), .Z(new_n745));
  OAI211_X1 g559(.A(new_n312), .B(new_n318), .C1(new_n280), .C2(new_n299), .ZN(new_n746));
  AOI22_X1  g560(.A1(new_n744), .A2(new_n745), .B1(new_n321), .B2(new_n746), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n747), .A2(new_n401), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n650), .A2(new_n706), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n748), .A2(new_n659), .A3(new_n729), .A4(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G122), .ZN(G24));
  AND2_X1   g566(.A1(new_n747), .A2(new_n671), .ZN(new_n753));
  INV_X1    g567(.A(new_n717), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n753), .A2(new_n650), .A3(new_n754), .A4(new_n729), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G125), .ZN(G27));
  NOR2_X1   g570(.A1(new_n405), .A2(new_n647), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n703), .A2(new_n649), .A3(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n608), .A2(new_n329), .ZN(new_n759));
  AOI21_X1  g573(.A(G902), .B1(new_n604), .B2(new_n606), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n759), .B1(new_n760), .B2(new_n608), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n593), .A2(KEYINPUT109), .A3(new_n560), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT109), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n580), .A2(new_n763), .ZN(new_n764));
  OAI211_X1 g578(.A(G469), .B(new_n589), .C1(new_n762), .C2(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n758), .B1(new_n761), .B2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n717), .A2(new_n767), .A3(KEYINPUT42), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n325), .A2(new_n768), .A3(new_n327), .A4(new_n401), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n715), .A2(new_n716), .A3(new_n766), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(new_n324), .A3(new_n401), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT42), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT110), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n769), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n773), .B1(new_n769), .B2(new_n772), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G131), .ZN(G33));
  NOR2_X1   g591(.A1(new_n767), .A2(new_n688), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n325), .A2(new_n327), .A3(new_n401), .A4(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G134), .ZN(G36));
  OAI211_X1 g594(.A(KEYINPUT45), .B(new_n589), .C1(new_n762), .C2(new_n764), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n587), .A2(new_n594), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n781), .B(G469), .C1(KEYINPUT45), .C2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n759), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(KEYINPUT46), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT111), .B1(new_n785), .B2(new_n609), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT46), .ZN(new_n788));
  INV_X1    g602(.A(new_n783), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n788), .B1(new_n789), .B2(new_n759), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n785), .A2(KEYINPUT111), .A3(new_n609), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n787), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(new_n406), .A3(new_n693), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT112), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n642), .A2(new_n544), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n796), .A2(KEYINPUT43), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(KEYINPUT43), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n797), .A2(new_n671), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n627), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT44), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n799), .A2(new_n627), .A3(KEYINPUT44), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n703), .A2(new_n407), .A3(new_n649), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n802), .A2(new_n803), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT113), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n802), .A2(KEYINPUT113), .A3(new_n803), .A4(new_n805), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n795), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G137), .ZN(G39));
  NAND2_X1  g626(.A1(new_n792), .A2(new_n406), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT47), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n791), .A2(new_n790), .ZN(new_n816));
  OAI211_X1 g630(.A(KEYINPUT47), .B(new_n406), .C1(new_n816), .C2(new_n786), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  OR3_X1    g632(.A1(new_n717), .A2(new_n401), .A3(new_n804), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n819), .B1(new_n325), .B2(new_n327), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n818), .A2(KEYINPUT114), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT47), .B1(new_n792), .B2(new_n406), .ZN(new_n822));
  INV_X1    g636(.A(new_n817), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n820), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n821), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(G140), .ZN(G42));
  INV_X1    g642(.A(new_n796), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n724), .A2(new_n609), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n705), .B(new_n829), .C1(KEYINPUT49), .C2(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n831), .B1(KEYINPUT49), .B2(new_n830), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n401), .A2(new_n757), .ZN(new_n833));
  XOR2_X1   g647(.A(new_n833), .B(KEYINPUT115), .Z(new_n834));
  INV_X1    g648(.A(new_n702), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n832), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT53), .ZN(new_n837));
  INV_X1    g651(.A(new_n628), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n704), .A2(new_n407), .A3(new_n659), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n839), .A2(new_n840), .A3(new_n645), .A4(new_n642), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n704), .A2(new_n407), .A3(new_n659), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT117), .B1(new_n646), .B2(new_n842), .ZN(new_n843));
  OR2_X1    g657(.A1(new_n468), .A2(new_n660), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n841), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n838), .A2(new_n625), .A3(new_n626), .A4(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n846), .B1(new_n402), .B2(new_n619), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n513), .A2(new_n544), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n687), .A2(new_n406), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n804), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n673), .A2(new_n674), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n610), .A2(new_n611), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n325), .A2(new_n853), .A3(new_n327), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n753), .A2(new_n770), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n779), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n681), .A2(new_n847), .A3(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n736), .A2(new_n731), .A3(new_n742), .A4(new_n751), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT116), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n751), .A2(new_n742), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n861), .A2(KEYINPUT116), .A3(new_n731), .A4(new_n736), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n857), .A2(new_n776), .A3(new_n860), .A4(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n761), .A2(new_n765), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n749), .A2(new_n671), .A3(new_n849), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n702), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n719), .A2(new_n690), .A3(new_n755), .A4(new_n866), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT52), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n837), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT54), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT52), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n867), .B(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n769), .A2(new_n772), .A3(KEYINPUT53), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n858), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n872), .A2(new_n857), .A3(new_n874), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n869), .A2(new_n870), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n548), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n797), .A2(new_n877), .A3(new_n798), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(new_n748), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n879), .A2(new_n804), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n830), .A2(new_n406), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n880), .B1(new_n818), .B2(new_n881), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n729), .A2(new_n805), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n835), .A2(new_n401), .A3(new_n877), .A4(new_n883), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n884), .A2(new_n645), .A3(new_n642), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n883), .A2(new_n878), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n753), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT120), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n886), .A2(KEYINPUT120), .A3(new_n753), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n885), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n705), .A2(new_n647), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n878), .A2(new_n748), .A3(new_n729), .A4(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT50), .ZN(new_n894));
  OAI21_X1  g708(.A(KEYINPUT119), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n893), .A2(new_n894), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n895), .B(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n882), .A2(new_n891), .A3(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT51), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n882), .A2(new_n891), .A3(KEYINPUT51), .A4(new_n897), .ZN(new_n901));
  OAI221_X1 g715(.A(new_n545), .B1(new_n740), .B2(new_n879), .C1(new_n884), .C2(new_n646), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n324), .A2(new_n401), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n886), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT48), .ZN(new_n905));
  OR2_X1    g719(.A1(new_n904), .A2(KEYINPUT48), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n902), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n900), .A2(new_n901), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n869), .A2(KEYINPUT118), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT118), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n910), .B(new_n837), .C1(new_n863), .C2(new_n868), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n863), .A2(new_n868), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n909), .B(new_n911), .C1(new_n837), .C2(new_n912), .ZN(new_n913));
  AOI211_X1 g727(.A(new_n876), .B(new_n908), .C1(new_n913), .C2(KEYINPUT54), .ZN(new_n914));
  NOR2_X1   g728(.A1(G952), .A2(G953), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n836), .B1(new_n914), .B2(new_n915), .ZN(G75));
  NOR2_X1   g730(.A1(new_n274), .A2(G952), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n329), .B1(new_n869), .B2(new_n875), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n920), .A2(new_n465), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n437), .A2(new_n444), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n922), .A2(new_n442), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n923), .A2(new_n446), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT55), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT56), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n918), .B1(new_n921), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n919), .A2(G210), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n925), .B1(new_n929), .B2(new_n926), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n928), .A2(new_n930), .ZN(G51));
  XNOR2_X1  g745(.A(new_n759), .B(KEYINPUT121), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT57), .Z(new_n933));
  AOI21_X1  g747(.A(new_n870), .B1(new_n869), .B2(new_n875), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n933), .B1(new_n876), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n607), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n919), .A2(new_n789), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n917), .B1(new_n936), .B2(new_n937), .ZN(G54));
  AND2_X1   g752(.A1(KEYINPUT58), .A2(G475), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n919), .A2(new_n535), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n535), .B1(new_n919), .B2(new_n939), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n940), .A2(new_n941), .A3(new_n917), .ZN(G60));
  NAND2_X1  g756(.A1(new_n634), .A2(new_n636), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n630), .B(KEYINPUT59), .Z(new_n944));
  OAI211_X1 g758(.A(new_n943), .B(new_n944), .C1(new_n876), .C2(new_n934), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n918), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n863), .A2(new_n868), .A3(new_n837), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n947), .B1(KEYINPUT118), .B2(new_n869), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n870), .B1(new_n948), .B2(new_n911), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n944), .B1(new_n949), .B2(new_n876), .ZN(new_n950));
  INV_X1    g764(.A(new_n943), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n946), .B1(new_n950), .B2(new_n951), .ZN(G63));
  NAND2_X1  g766(.A1(new_n869), .A2(new_n875), .ZN(new_n953));
  NAND2_X1  g767(.A1(G217), .A2(G902), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT60), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n391), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n917), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT61), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n955), .B1(new_n869), .B2(new_n875), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n669), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n959), .A2(KEYINPUT122), .A3(new_n960), .A4(new_n962), .ZN(new_n963));
  OR2_X1    g777(.A1(new_n960), .A2(KEYINPUT122), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n960), .A2(KEYINPUT122), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n918), .B1(new_n961), .B2(new_n391), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n953), .A2(new_n669), .A3(new_n956), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n964), .B(new_n965), .C1(new_n966), .C2(new_n967), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n963), .A2(new_n968), .ZN(G66));
  AOI21_X1  g783(.A(new_n274), .B1(new_n550), .B2(G224), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n681), .A2(new_n847), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n860), .A2(new_n862), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n970), .B1(new_n972), .B2(new_n274), .ZN(new_n973));
  INV_X1    g787(.A(G898), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n922), .B1(new_n974), .B2(G953), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n973), .B(new_n975), .ZN(G69));
  INV_X1    g790(.A(G900), .ZN(new_n977));
  OAI21_X1  g791(.A(G953), .B1(new_n557), .B2(new_n977), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT125), .Z(new_n979));
  NAND2_X1  g793(.A1(new_n827), .A2(new_n811), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n903), .A2(new_n750), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n795), .A2(new_n981), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n690), .A2(new_n755), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n983), .A2(new_n719), .A3(new_n779), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n982), .A2(new_n776), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(KEYINPUT126), .B1(new_n980), .B2(new_n985), .ZN(new_n986));
  AOI22_X1  g800(.A1(new_n821), .A2(new_n826), .B1(new_n795), .B2(new_n810), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT126), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n984), .A2(new_n776), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n987), .A2(new_n988), .A3(new_n982), .A4(new_n989), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n986), .A2(new_n990), .A3(new_n274), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n291), .A2(new_n292), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(new_n531), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n993), .B1(G900), .B2(G953), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n993), .B(KEYINPUT123), .Z(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n983), .A2(new_n709), .A3(new_n719), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT62), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n983), .A2(KEYINPUT62), .A3(new_n709), .A4(new_n719), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n646), .B1(new_n513), .B2(new_n645), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n1003), .A2(KEYINPUT124), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(KEYINPUT124), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n805), .ZN(new_n1006));
  OR4_X1    g820(.A1(new_n402), .A2(new_n694), .A3(new_n1004), .A4(new_n1006), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n827), .A2(new_n1002), .A3(new_n811), .A4(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n997), .B1(new_n1008), .B2(new_n274), .ZN(new_n1009));
  INV_X1    g823(.A(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n979), .B1(new_n995), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(new_n979), .ZN(new_n1012));
  AOI211_X1 g826(.A(new_n1012), .B(new_n1009), .C1(new_n991), .C2(new_n994), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n1011), .A2(new_n1013), .ZN(G72));
  XOR2_X1   g828(.A(KEYINPUT127), .B(KEYINPUT63), .Z(new_n1015));
  NOR2_X1   g829(.A1(new_n622), .A2(new_n329), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1015), .B(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(new_n295), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n699), .B1(new_n1018), .B2(new_n300), .ZN(new_n1019));
  AOI211_X1 g833(.A(new_n1017), .B(new_n1019), .C1(new_n948), .C2(new_n911), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n1018), .A2(new_n278), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n986), .A2(new_n990), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1018), .A2(new_n278), .ZN(new_n1023));
  OR2_X1    g837(.A1(new_n1008), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n972), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(new_n1023), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1017), .B1(new_n1026), .B2(new_n1021), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1027), .A2(new_n918), .ZN(new_n1028));
  NOR3_X1   g842(.A1(new_n1020), .A2(new_n1025), .A3(new_n1028), .ZN(G57));
endmodule


