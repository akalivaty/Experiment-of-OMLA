//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 0 1 1 1 0 1 1 0 0 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 0 0 1 1 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983;
  INV_X1    g000(.A(G104), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT3), .B1(new_n187), .B2(G107), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G104), .ZN(new_n191));
  INV_X1    g005(.A(G101), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n187), .A2(G107), .ZN(new_n193));
  NAND4_X1  g007(.A1(new_n188), .A2(new_n191), .A3(new_n192), .A4(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n187), .A2(G107), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n190), .A2(G104), .ZN(new_n196));
  OAI21_X1  g010(.A(G101), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT5), .ZN(new_n200));
  INV_X1    g014(.A(G119), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(G116), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT72), .ZN(new_n203));
  INV_X1    g017(.A(G116), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(G119), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n201), .A2(KEYINPUT72), .A3(G116), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(G119), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  OAI211_X1 g022(.A(G113), .B(new_n202), .C1(new_n208), .C2(new_n200), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT2), .B(G113), .ZN(new_n210));
  OR2_X1    g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n199), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n188), .A2(new_n191), .A3(new_n193), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G101), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT84), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AND2_X1   g030(.A1(new_n194), .A2(KEYINPUT4), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n213), .A2(KEYINPUT84), .A3(G101), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT4), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n213), .A2(new_n221), .A3(G101), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n208), .A2(KEYINPUT71), .A3(new_n210), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n210), .B1(new_n208), .B2(KEYINPUT71), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n212), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(G110), .B(G122), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n227), .B(new_n212), .C1(new_n220), .C2(new_n225), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(KEYINPUT6), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT65), .ZN(new_n232));
  INV_X1    g046(.A(G143), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n232), .B1(new_n233), .B2(G146), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(G146), .ZN(new_n235));
  INV_X1    g049(.A(G146), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(KEYINPUT65), .A3(G143), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n234), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  AND2_X1   g052(.A1(KEYINPUT0), .A2(G128), .ZN(new_n239));
  NOR2_X1   g053(.A1(KEYINPUT0), .A2(G128), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT66), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n243), .B1(new_n233), .B2(G146), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n236), .A2(KEYINPUT66), .A3(G143), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n244), .A2(new_n245), .A3(new_n235), .A4(new_n239), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n242), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G125), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n244), .A2(new_n245), .A3(new_n235), .ZN(new_n249));
  OR2_X1    g063(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n250));
  NAND2_X1  g064(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n250), .A2(G128), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n249), .A2(new_n253), .ZN(new_n254));
  AOI22_X1  g068(.A1(new_n250), .A2(new_n251), .B1(G143), .B2(new_n236), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT70), .B(G128), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n238), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G125), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n254), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n248), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G953), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G224), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n262), .B(KEYINPUT86), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n260), .B(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT6), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n226), .A2(new_n265), .A3(new_n228), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n231), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  XOR2_X1   g081(.A(new_n227), .B(KEYINPUT8), .Z(new_n268));
  NAND2_X1  g082(.A1(new_n209), .A2(new_n211), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n198), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n268), .B1(new_n270), .B2(new_n212), .ZN(new_n271));
  AND4_X1   g085(.A1(KEYINPUT7), .A2(new_n248), .A3(new_n259), .A4(new_n262), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n248), .A2(new_n259), .B1(KEYINPUT7), .B2(new_n262), .ZN(new_n273));
  NOR3_X1   g087(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(G902), .B1(new_n274), .B2(new_n230), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n267), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(G210), .B1(G237), .B2(G902), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n277), .B(KEYINPUT87), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  AND3_X1   g093(.A1(new_n267), .A2(new_n275), .A3(new_n277), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G237), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n283), .A2(new_n261), .A3(G214), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n284), .B(G143), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT18), .ZN(new_n286));
  INV_X1    g100(.A(G131), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n284), .B(new_n233), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(KEYINPUT18), .A3(G131), .ZN(new_n290));
  XNOR2_X1  g104(.A(G125), .B(G140), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n291), .B(new_n236), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n288), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(KEYINPUT16), .ZN(new_n294));
  OR3_X1    g108(.A1(new_n258), .A2(KEYINPUT16), .A3(G140), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n294), .A2(G146), .A3(new_n295), .ZN(new_n296));
  XOR2_X1   g110(.A(new_n291), .B(KEYINPUT19), .Z(new_n297));
  OAI21_X1  g111(.A(new_n296), .B1(new_n297), .B2(G146), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n289), .A2(G131), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n285), .A2(new_n287), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n293), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  XOR2_X1   g116(.A(G113), .B(G122), .Z(new_n303));
  XOR2_X1   g117(.A(KEYINPUT88), .B(G104), .Z(new_n304));
  XOR2_X1   g118(.A(new_n303), .B(new_n304), .Z(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT17), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n299), .A2(new_n300), .A3(new_n308), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n294), .A2(G146), .A3(new_n295), .ZN(new_n310));
  AOI21_X1  g124(.A(G146), .B1(new_n294), .B2(new_n295), .ZN(new_n311));
  OAI21_X1  g125(.A(KEYINPUT89), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n294), .A2(new_n295), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n236), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT89), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n314), .A2(new_n315), .A3(new_n296), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n289), .A2(KEYINPUT17), .A3(G131), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n309), .A2(new_n312), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(new_n293), .A3(new_n305), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n307), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT20), .ZN(new_n321));
  NOR2_X1   g135(.A1(G475), .A2(G902), .ZN(new_n322));
  AND3_X1   g136(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n321), .B1(new_n320), .B2(new_n322), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n318), .A2(new_n293), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n306), .ZN(new_n326));
  AOI21_X1  g140(.A(G902), .B1(new_n326), .B2(new_n319), .ZN(new_n327));
  XOR2_X1   g141(.A(KEYINPUT90), .B(G475), .Z(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  OAI22_X1  g143(.A1(new_n323), .A2(new_n324), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G134), .ZN(new_n331));
  INV_X1    g145(.A(G128), .ZN(new_n332));
  OAI21_X1  g146(.A(KEYINPUT91), .B1(new_n332), .B2(G143), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT91), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(new_n233), .A3(G128), .ZN(new_n335));
  AOI21_X1  g149(.A(KEYINPUT13), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n336), .A2(KEYINPUT92), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n256), .A2(G143), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n333), .A2(new_n335), .A3(KEYINPUT13), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n336), .A2(KEYINPUT92), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n331), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(G116), .B(G122), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(new_n190), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n333), .A2(new_n335), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n338), .A2(new_n331), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  OR2_X1    g162(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT93), .ZN(new_n350));
  OR2_X1    g164(.A1(new_n204), .A2(G122), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n190), .B1(new_n351), .B2(KEYINPUT14), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n352), .B(new_n344), .ZN(new_n353));
  INV_X1    g167(.A(new_n347), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n331), .B1(new_n338), .B2(new_n346), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT9), .B(G234), .ZN(new_n357));
  INV_X1    g171(.A(G217), .ZN(new_n358));
  NOR3_X1   g172(.A1(new_n357), .A2(new_n358), .A3(G953), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n349), .A2(new_n350), .A3(new_n356), .A4(new_n359), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n356), .B(new_n359), .C1(new_n343), .C2(new_n348), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT93), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n356), .B1(new_n343), .B2(new_n348), .ZN(new_n363));
  INV_X1    g177(.A(new_n359), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n360), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G902), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G478), .ZN(new_n369));
  NOR2_X1   g183(.A1(KEYINPUT94), .A2(KEYINPUT15), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(KEYINPUT94), .A2(KEYINPUT15), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n369), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n373), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n375), .B1(new_n366), .B2(new_n367), .ZN(new_n376));
  NAND2_X1  g190(.A1(G234), .A2(G237), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n377), .A2(G952), .A3(new_n261), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(G902), .A3(G953), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(KEYINPUT21), .B(G898), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n379), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NOR4_X1   g197(.A1(new_n330), .A2(new_n374), .A3(new_n376), .A4(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(G214), .B1(G237), .B2(G902), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n282), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G469), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n331), .A2(G137), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT11), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(KEYINPUT67), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT67), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(KEYINPUT11), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G137), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n394), .A2(G134), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n388), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT68), .ZN(new_n398));
  NAND2_X1  g212(.A1(KEYINPUT11), .A2(G134), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n398), .B1(new_n399), .B2(G137), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n394), .A2(KEYINPUT68), .A3(KEYINPUT11), .A4(G134), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(G131), .B1(new_n397), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n400), .A2(new_n401), .ZN(new_n404));
  AOI22_X1  g218(.A1(new_n390), .A2(new_n392), .B1(new_n331), .B2(G137), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n404), .B(new_n287), .C1(new_n405), .C2(new_n388), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n236), .A2(G143), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n332), .B1(new_n408), .B2(KEYINPUT1), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n249), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n244), .A2(new_n245), .A3(new_n235), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(new_n252), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n199), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n254), .A2(new_n257), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n415), .A2(new_n199), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n407), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(KEYINPUT12), .ZN(new_n418));
  AOI21_X1  g232(.A(KEYINPUT65), .B1(new_n236), .B2(G143), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n236), .A2(G143), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AND2_X1   g235(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n422));
  NOR2_X1   g236(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n408), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n332), .A2(KEYINPUT70), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT70), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(G128), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n421), .A2(new_n237), .B1(new_n424), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(KEYINPUT74), .B1(new_n429), .B2(new_n412), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT74), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n254), .A2(new_n257), .A3(new_n431), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n430), .A2(new_n432), .A3(KEYINPUT10), .A4(new_n199), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT10), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n413), .A2(new_n434), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n222), .A2(new_n246), .A3(new_n242), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n219), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n407), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n433), .A2(new_n435), .A3(new_n437), .A4(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(G110), .B(G140), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n261), .A2(G227), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n440), .B(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT12), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n444), .B(new_n407), .C1(new_n414), .C2(new_n416), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n418), .A2(new_n439), .A3(new_n443), .A4(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n433), .A2(new_n437), .A3(new_n435), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n407), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n443), .B1(new_n448), .B2(new_n439), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n446), .B1(new_n449), .B2(KEYINPUT85), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT85), .ZN(new_n451));
  AOI211_X1 g265(.A(new_n451), .B(new_n443), .C1(new_n448), .C2(new_n439), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n387), .B(new_n367), .C1(new_n450), .C2(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n387), .A2(new_n367), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  AND2_X1   g269(.A1(new_n448), .A2(new_n439), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n443), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n418), .A2(new_n439), .A3(new_n445), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n442), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n453), .B(new_n455), .C1(new_n387), .C2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G221), .ZN(new_n462));
  INV_X1    g276(.A(new_n357), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n462), .B1(new_n463), .B2(new_n367), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n386), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(G472), .A2(G902), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT32), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n223), .A2(new_n224), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n242), .A2(new_n246), .ZN(new_n473));
  INV_X1    g287(.A(new_n406), .ZN(new_n474));
  INV_X1    g288(.A(new_n388), .ZN(new_n475));
  XNOR2_X1  g289(.A(KEYINPUT67), .B(KEYINPUT11), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n475), .B1(new_n476), .B2(new_n395), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n287), .B1(new_n477), .B2(new_n404), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n473), .B1(new_n474), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(G131), .B1(new_n388), .B2(new_n395), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n415), .A2(new_n406), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  XOR2_X1   g296(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n483));
  AOI21_X1  g297(.A(new_n472), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n479), .A2(KEYINPUT73), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n406), .A2(new_n480), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(new_n430), .A3(new_n432), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT73), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n488), .B(new_n473), .C1(new_n474), .C2(new_n478), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n485), .A2(KEYINPUT30), .A3(new_n487), .A4(new_n489), .ZN(new_n490));
  AND2_X1   g304(.A1(new_n484), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n485), .A2(new_n487), .A3(new_n472), .A4(new_n489), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n283), .A2(new_n261), .A3(G210), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n493), .B(KEYINPUT27), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT26), .B(G101), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n494), .B(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(KEYINPUT31), .B1(new_n491), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(KEYINPUT75), .ZN(new_n499));
  INV_X1    g313(.A(new_n496), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT28), .ZN(new_n501));
  INV_X1    g315(.A(new_n472), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n482), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n501), .B1(new_n492), .B2(new_n503), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n487), .A2(new_n472), .ZN(new_n505));
  AOI21_X1  g319(.A(KEYINPUT28), .B1(new_n505), .B2(new_n479), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n500), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n489), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n488), .B1(new_n407), .B2(new_n473), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n500), .B1(new_n510), .B2(new_n505), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n484), .A2(new_n490), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT31), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n511), .A2(new_n512), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT75), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT31), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n499), .A2(new_n507), .A3(new_n514), .A4(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n518), .A2(KEYINPUT76), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT76), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n516), .B1(new_n515), .B2(KEYINPUT31), .ZN(new_n521));
  AOI211_X1 g335(.A(KEYINPUT75), .B(new_n513), .C1(new_n511), .C2(new_n512), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AND2_X1   g337(.A1(new_n507), .A2(new_n514), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n520), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n471), .B1(new_n519), .B2(new_n525), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n510), .A2(new_n487), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n492), .B1(new_n527), .B2(new_n472), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT28), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n506), .B(KEYINPUT78), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT29), .A4(new_n496), .ZN(new_n531));
  OR3_X1    g345(.A1(new_n504), .A2(new_n506), .A3(new_n500), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT29), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n512), .A2(new_n492), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n500), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n532), .A2(KEYINPUT77), .A3(new_n533), .A4(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT77), .ZN(new_n537));
  AOI22_X1  g351(.A1(new_n490), .A2(new_n484), .B1(new_n510), .B2(new_n505), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n533), .B1(new_n538), .B2(new_n496), .ZN(new_n539));
  NOR3_X1   g353(.A1(new_n504), .A2(new_n506), .A3(new_n500), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n531), .A2(new_n536), .A3(new_n367), .A4(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G472), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n518), .A2(KEYINPUT76), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n523), .A2(new_n520), .A3(new_n524), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n469), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n526), .B(new_n543), .C1(new_n546), .C2(KEYINPUT32), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT83), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n358), .B1(G234), .B2(new_n367), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n549), .A2(G902), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT22), .B(G137), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n261), .A2(G221), .A3(G234), .ZN(new_n552));
  XOR2_X1   g366(.A(new_n551), .B(new_n552), .Z(new_n553));
  NAND3_X1  g367(.A1(new_n256), .A2(KEYINPUT23), .A3(G119), .ZN(new_n554));
  AOI21_X1  g368(.A(KEYINPUT23), .B1(new_n332), .B2(G119), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n555), .B1(new_n201), .B2(G128), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(KEYINPUT79), .B1(new_n557), .B2(G110), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n201), .A2(G128), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n559), .B1(new_n428), .B2(new_n201), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT24), .B(G110), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT79), .ZN(new_n563));
  INV_X1    g377(.A(G110), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n554), .A2(new_n556), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n558), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n310), .B1(new_n236), .B2(new_n291), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n557), .A2(G110), .ZN(new_n569));
  OAI221_X1 g383(.A(new_n569), .B1(new_n560), .B2(new_n561), .C1(new_n311), .C2(new_n310), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n568), .A2(KEYINPUT80), .A3(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT80), .B1(new_n568), .B2(new_n570), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n553), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n553), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n575), .A2(new_n578), .A3(KEYINPUT82), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT82), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n580), .B1(new_n574), .B2(new_n577), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n574), .A2(new_n367), .A3(new_n577), .ZN(new_n583));
  NAND2_X1  g397(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n586));
  OR3_X1    g400(.A1(new_n583), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n549), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n588), .B1(new_n583), .B2(new_n585), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n550), .A2(new_n582), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n547), .A2(new_n548), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n548), .B1(new_n547), .B2(new_n590), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n467), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(G101), .ZN(G3));
  AND3_X1   g409(.A1(new_n590), .A2(new_n465), .A3(new_n461), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n468), .B1(new_n519), .B2(new_n525), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n367), .B1(new_n519), .B2(new_n525), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(G472), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n596), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n277), .B1(new_n267), .B2(new_n275), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n385), .B1(new_n280), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT95), .ZN(new_n603));
  INV_X1    g417(.A(new_n383), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT95), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n605), .B(new_n385), .C1(new_n280), .C2(new_n601), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n603), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT96), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT33), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n609), .B1(new_n363), .B2(new_n364), .ZN(new_n610));
  AOI22_X1  g424(.A1(new_n366), .A2(new_n609), .B1(new_n361), .B2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n369), .A2(G902), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(G478), .B1(new_n366), .B2(new_n367), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n608), .B1(new_n616), .B2(new_n330), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n614), .B1(new_n611), .B2(new_n612), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n320), .A2(new_n322), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT20), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n326), .A2(new_n319), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n367), .ZN(new_n623));
  AOI22_X1  g437(.A1(new_n620), .A2(new_n621), .B1(new_n623), .B2(new_n328), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n618), .A2(new_n624), .A3(KEYINPUT96), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n617), .A2(new_n625), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n600), .A2(new_n607), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT34), .B(G104), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G6));
  OAI21_X1  g443(.A(new_n624), .B1(new_n374), .B2(new_n376), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n600), .A2(new_n607), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(KEYINPUT35), .B(G107), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G9));
  NAND2_X1  g447(.A1(new_n587), .A2(new_n589), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n568), .A2(new_n570), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n576), .A2(KEYINPUT36), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n550), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n466), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n640), .A2(new_n597), .A3(new_n386), .A4(new_n599), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT37), .B(G110), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G12));
  NAND2_X1  g457(.A1(new_n603), .A2(new_n606), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n597), .A2(new_n470), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n544), .A2(new_n545), .ZN(new_n646));
  AOI22_X1  g460(.A1(new_n646), .A2(new_n471), .B1(G472), .B2(new_n542), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n644), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n648), .A2(new_n640), .ZN(new_n649));
  OR2_X1    g463(.A1(new_n380), .A2(G900), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n378), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n630), .A2(new_n652), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(new_n332), .ZN(G30));
  NAND2_X1  g469(.A1(new_n534), .A2(new_n496), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n656), .B(new_n367), .C1(new_n528), .C2(new_n496), .ZN(new_n657));
  AOI22_X1  g471(.A1(new_n646), .A2(new_n471), .B1(G472), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n645), .A2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n651), .B(KEYINPUT39), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n466), .A2(new_n661), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n662), .A2(KEYINPUT40), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n281), .B(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n639), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n330), .B1(new_n374), .B2(new_n376), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n665), .A2(new_n385), .A3(new_n666), .A4(new_n668), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n660), .A2(new_n663), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n670), .B1(KEYINPUT40), .B2(new_n662), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G143), .ZN(G45));
  INV_X1    g486(.A(new_n612), .ZN(new_n673));
  AOI221_X4 g487(.A(new_n673), .B1(new_n610), .B2(new_n361), .C1(new_n366), .C2(new_n609), .ZN(new_n674));
  OAI211_X1 g488(.A(new_n330), .B(new_n651), .C1(new_n674), .C2(new_n614), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT98), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n616), .A2(KEYINPUT98), .A3(new_n330), .A4(new_n651), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n649), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(new_n236), .ZN(G48));
  NOR2_X1   g496(.A1(new_n626), .A2(new_n607), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n367), .B1(new_n450), .B2(new_n452), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(G469), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n465), .A3(new_n453), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT99), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n547), .A2(new_n683), .A3(new_n688), .A4(new_n590), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT41), .B(G113), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G15));
  NOR2_X1   g505(.A1(new_n607), .A2(new_n630), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n547), .A2(new_n688), .A3(new_n590), .A4(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(KEYINPUT100), .ZN(new_n694));
  INV_X1    g508(.A(new_n590), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n695), .B1(new_n645), .B2(new_n647), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT100), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n696), .A2(new_n697), .A3(new_n692), .A4(new_n688), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT101), .B(G116), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G18));
  NOR2_X1   g515(.A1(new_n644), .A2(new_n686), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n639), .A2(new_n384), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n547), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G119), .ZN(G21));
  NAND2_X1  g519(.A1(new_n529), .A2(new_n530), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n500), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n498), .A2(new_n514), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n469), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n709), .B1(new_n598), .B2(G472), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n644), .A2(new_n383), .A3(new_n667), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n710), .A2(new_n688), .A3(new_n590), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G122), .ZN(G24));
  INV_X1    g527(.A(new_n709), .ZN(new_n714));
  AOI21_X1  g528(.A(G902), .B1(new_n544), .B2(new_n545), .ZN(new_n715));
  INV_X1    g529(.A(G472), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n639), .B(new_n714), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT102), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n679), .A2(new_n644), .A3(new_n686), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n680), .A2(new_n702), .ZN(new_n722));
  OAI21_X1  g536(.A(KEYINPUT102), .B1(new_n722), .B2(new_n717), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G125), .ZN(G27));
  AOI21_X1  g539(.A(KEYINPUT32), .B1(new_n646), .B2(new_n468), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(KEYINPUT105), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT105), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n728), .B1(new_n546), .B2(KEYINPUT32), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n727), .A2(new_n647), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n457), .A2(KEYINPUT103), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT103), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n456), .A2(new_n732), .A3(new_n443), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n731), .A2(new_n459), .A3(new_n733), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n453), .B(new_n455), .C1(new_n734), .C2(new_n387), .ZN(new_n735));
  INV_X1    g549(.A(new_n385), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n464), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n735), .A2(new_n281), .A3(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT42), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n679), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n730), .A2(new_n590), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n679), .A2(new_n738), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT104), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n547), .A2(new_n742), .A3(new_n743), .A4(new_n590), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n739), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n743), .B1(new_n696), .B2(new_n742), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n741), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(KEYINPUT106), .B(G131), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(G33));
  INV_X1    g563(.A(new_n738), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n696), .A2(new_n653), .A3(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G134), .ZN(G36));
  NOR2_X1   g566(.A1(new_n618), .A2(new_n330), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(KEYINPUT43), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n599), .A2(new_n597), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n755), .A2(KEYINPUT108), .A3(new_n639), .ZN(new_n756));
  AOI21_X1  g570(.A(KEYINPUT108), .B1(new_n755), .B2(new_n639), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n754), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n759));
  OR2_X1    g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n453), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT45), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n387), .B1(new_n460), .B2(new_n762), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n731), .A2(KEYINPUT45), .A3(new_n459), .A4(new_n733), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT107), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n765), .B1(new_n763), .B2(new_n764), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n455), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT46), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n761), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI211_X1 g584(.A(KEYINPUT46), .B(new_n455), .C1(new_n766), .C2(new_n767), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n772), .A2(new_n465), .A3(new_n661), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n281), .A2(new_n385), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n758), .A2(new_n759), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n760), .A2(new_n773), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(KEYINPUT109), .B(G137), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n777), .B(new_n778), .ZN(G39));
  NOR4_X1   g593(.A1(new_n547), .A2(new_n590), .A3(new_n679), .A4(new_n774), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n772), .A2(KEYINPUT47), .A3(new_n465), .ZN(new_n781));
  AOI21_X1  g595(.A(KEYINPUT47), .B1(new_n772), .B2(new_n465), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G140), .ZN(G42));
  OAI211_X1 g598(.A(new_n630), .B(KEYINPUT113), .C1(new_n624), .C2(new_n618), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT113), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n616), .A2(new_n786), .A3(new_n330), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n282), .A2(new_n385), .A3(new_n604), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n790), .A2(new_n597), .A3(new_n599), .A4(new_n596), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n641), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n526), .A2(new_n543), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n590), .B1(new_n793), .B2(new_n726), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(KEYINPUT83), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n591), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n792), .B1(new_n796), .B2(new_n467), .ZN(new_n797));
  NOR4_X1   g611(.A1(new_n330), .A2(new_n374), .A3(new_n376), .A4(new_n652), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n547), .A2(new_n775), .A3(new_n798), .ZN(new_n799));
  AOI22_X1  g613(.A1(new_n799), .A2(new_n640), .B1(new_n718), .B2(new_n742), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n797), .A2(new_n747), .A3(new_n751), .A4(new_n800), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n648), .B(new_n640), .C1(new_n653), .C2(new_n680), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT114), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n465), .B1(new_n652), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n804), .B1(new_n803), .B2(new_n652), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n666), .A2(new_n735), .A3(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n644), .A2(new_n667), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n806), .A2(new_n659), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n724), .A2(new_n802), .A3(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n724), .A2(new_n802), .A3(KEYINPUT52), .A4(new_n808), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n801), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n689), .A2(new_n712), .A3(new_n704), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT112), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n699), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n815), .B1(new_n699), .B2(new_n814), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT53), .B1(new_n813), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n811), .A2(new_n812), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n747), .A2(new_n751), .ZN(new_n821));
  INV_X1    g635(.A(new_n792), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n594), .A2(new_n800), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  AND4_X1   g638(.A1(KEYINPUT53), .A2(new_n818), .A3(new_n820), .A4(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(KEYINPUT54), .B1(new_n819), .B2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n824), .A2(new_n820), .ZN(new_n828));
  OR2_X1    g642(.A1(new_n816), .A2(new_n817), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n699), .A2(new_n814), .A3(KEYINPUT53), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n824), .A2(new_n820), .A3(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n830), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n774), .A2(new_n686), .ZN(new_n835));
  AND4_X1   g649(.A1(new_n590), .A2(new_n660), .A3(new_n379), .A4(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n616), .A2(new_n330), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n754), .A2(new_n379), .A3(new_n835), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n718), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT115), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n839), .A2(new_n718), .A3(KEYINPUT115), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n838), .A2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n782), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n772), .A2(KEYINPUT47), .A3(new_n465), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n685), .A2(new_n453), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(new_n464), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  AND4_X1   g664(.A1(new_n590), .A2(new_n710), .A3(new_n379), .A4(new_n754), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(new_n775), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n665), .A2(new_n385), .A3(new_n686), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT50), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n856), .B(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n845), .A2(new_n854), .A3(KEYINPUT51), .A4(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(G952), .ZN(new_n860));
  AOI211_X1 g674(.A(new_n860), .B(G953), .C1(new_n851), .C2(new_n702), .ZN(new_n861));
  INV_X1    g675(.A(new_n626), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n836), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n730), .A2(new_n590), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n839), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n866), .A2(KEYINPUT48), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(KEYINPUT48), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n864), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n859), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT51), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n856), .A2(new_n857), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT50), .B1(new_n851), .B2(new_n855), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n844), .B(new_n838), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n781), .A2(new_n782), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n852), .B1(new_n875), .B2(new_n849), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n871), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT116), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI211_X1 g693(.A(KEYINPUT116), .B(new_n871), .C1(new_n874), .C2(new_n876), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n870), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n826), .A2(new_n834), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT117), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT117), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n826), .A2(new_n881), .A3(new_n884), .A4(new_n834), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n860), .A2(new_n261), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n883), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT49), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n848), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n590), .A2(new_n737), .A3(new_n753), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT110), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n892), .B1(new_n891), .B2(new_n890), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT111), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n665), .B1(new_n848), .B2(new_n888), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n894), .A2(new_n660), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n887), .A2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT118), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n887), .A2(KEYINPUT118), .A3(new_n896), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(G75));
  NOR2_X1   g715(.A1(new_n261), .A2(G952), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n830), .A2(new_n833), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n904), .A2(new_n367), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT56), .B1(new_n905), .B2(G210), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n231), .A2(new_n266), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(new_n264), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT55), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n903), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n905), .A2(new_n278), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT119), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT56), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n909), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n910), .B1(new_n912), .B2(new_n914), .ZN(G51));
  XNOR2_X1  g729(.A(new_n904), .B(new_n831), .ZN(new_n916));
  XNOR2_X1  g730(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(new_n454), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n919), .B1(new_n452), .B2(new_n450), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n766), .A2(new_n767), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n905), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n902), .B1(new_n920), .B2(new_n922), .ZN(G54));
  AND3_X1   g737(.A1(new_n905), .A2(KEYINPUT58), .A3(G475), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n903), .B1(new_n924), .B2(new_n320), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n925), .B1(new_n320), .B2(new_n924), .ZN(G60));
  NAND2_X1  g740(.A1(new_n826), .A2(new_n834), .ZN(new_n927));
  XNOR2_X1  g741(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n928));
  NAND2_X1  g742(.A1(G478), .A2(G902), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n928), .B(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n611), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n611), .A2(new_n930), .ZN(new_n932));
  AOI211_X1 g746(.A(new_n902), .B(new_n931), .C1(new_n916), .C2(new_n932), .ZN(G63));
  XNOR2_X1  g747(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n934));
  NAND2_X1  g748(.A1(G217), .A2(G902), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n934), .B(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n904), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n637), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n938), .B(new_n903), .C1(new_n582), .C2(new_n937), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT61), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(G66));
  INV_X1    g755(.A(G224), .ZN(new_n942));
  OAI21_X1  g756(.A(G953), .B1(new_n382), .B2(new_n942), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n818), .A2(new_n797), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n943), .B1(new_n944), .B2(G953), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n907), .B1(G898), .B2(new_n261), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT124), .Z(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT123), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n945), .B(new_n948), .ZN(G69));
  NAND2_X1  g763(.A1(new_n482), .A2(new_n483), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n490), .A2(new_n950), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(new_n297), .Z(new_n952));
  AOI21_X1  g766(.A(new_n952), .B1(G900), .B2(G953), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n773), .A2(new_n807), .A3(new_n865), .ZN(new_n954));
  AND4_X1   g768(.A1(new_n747), .A2(new_n783), .A3(new_n954), .A4(new_n751), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n724), .A2(new_n802), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n777), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n956), .B1(new_n777), .B2(new_n957), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n955), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n953), .B1(new_n960), .B2(G953), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n261), .B1(G227), .B2(G900), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(KEYINPUT127), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n662), .A2(new_n788), .A3(new_n774), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n796), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n777), .A2(new_n783), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n957), .A2(new_n671), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT62), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n969), .A2(G953), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n952), .B(KEYINPUT125), .Z(new_n971));
  OAI211_X1 g785(.A(new_n961), .B(new_n963), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n962), .A2(KEYINPUT127), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n972), .B(new_n973), .Z(G72));
  OAI211_X1 g788(.A(new_n944), .B(new_n955), .C1(new_n958), .C2(new_n959), .ZN(new_n975));
  NAND2_X1  g789(.A1(G472), .A2(G902), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT63), .Z(new_n977));
  AOI211_X1 g791(.A(new_n496), .B(new_n534), .C1(new_n975), .C2(new_n977), .ZN(new_n978));
  OR2_X1    g792(.A1(new_n819), .A2(new_n825), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n535), .A2(new_n515), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n979), .A2(new_n977), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n969), .A2(new_n944), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n656), .B1(new_n982), .B2(new_n977), .ZN(new_n983));
  NOR4_X1   g797(.A1(new_n978), .A2(new_n981), .A3(new_n902), .A4(new_n983), .ZN(G57));
endmodule


