//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 0 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1244, new_n1245, new_n1246, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND3_X1  g0013(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n214));
  INV_X1    g0014(.A(new_n201), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n210), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n213), .B1(new_n214), .B2(new_n216), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G58), .B(G77), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(KEYINPUT17), .ZN(new_n244));
  INV_X1    g0044(.A(KEYINPUT70), .ZN(new_n245));
  NAND2_X1  g0045(.A1(G58), .A2(G68), .ZN(new_n246));
  AOI21_X1  g0046(.A(new_n208), .B1(new_n215), .B2(new_n246), .ZN(new_n247));
  NOR2_X1   g0047(.A1(G20), .A2(G33), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G159), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n245), .B1(new_n247), .B2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(new_n246), .ZN(new_n253));
  OAI21_X1  g0053(.A(G20), .B1(new_n253), .B2(new_n201), .ZN(new_n254));
  OAI211_X1 g0054(.A(new_n254), .B(KEYINPUT70), .C1(new_n250), .C2(new_n249), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT7), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT3), .B(G33), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n257), .B1(new_n258), .B2(G20), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT3), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n218), .B1(new_n259), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT16), .ZN(new_n267));
  OR3_X1    g0067(.A1(new_n256), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n261), .A2(KEYINPUT71), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT71), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(new_n260), .A3(KEYINPUT3), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n269), .A2(new_n263), .A3(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n257), .A2(G20), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n218), .B1(new_n274), .B2(new_n259), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n267), .B1(new_n275), .B2(new_n256), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G1), .A2(G13), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n268), .A2(new_n276), .A3(new_n279), .ZN(new_n280));
  XOR2_X1   g0080(.A(KEYINPUT8), .B(G58), .Z(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n282), .B1(new_n207), .B2(G20), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(new_n279), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n283), .A2(new_n286), .B1(new_n285), .B2(new_n282), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n280), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G200), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT73), .ZN(new_n291));
  INV_X1    g0091(.A(G223), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(G1698), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n293), .A2(new_n261), .A3(new_n263), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT72), .ZN(new_n295));
  NAND2_X1  g0095(.A1(G33), .A2(G87), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n261), .A2(new_n263), .A3(G226), .A4(G1698), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT72), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n293), .A2(new_n261), .A3(new_n263), .A4(new_n298), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n295), .A2(new_n296), .A3(new_n297), .A4(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G33), .A2(G41), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n301), .A2(G1), .A3(G13), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G41), .ZN(new_n305));
  INV_X1    g0105(.A(G45), .ZN(new_n306));
  AOI21_X1  g0106(.A(G1), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n307), .A2(new_n302), .A3(G274), .ZN(new_n308));
  INV_X1    g0108(.A(G232), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n302), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n308), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n291), .B1(new_n304), .B2(new_n313), .ZN(new_n314));
  AOI211_X1 g0114(.A(KEYINPUT73), .B(new_n312), .C1(new_n300), .C2(new_n303), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n290), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT75), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n298), .B1(new_n258), .B2(new_n293), .ZN(new_n318));
  AND4_X1   g0118(.A1(new_n298), .A2(new_n293), .A3(new_n261), .A4(new_n263), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n297), .A2(new_n296), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n302), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NOR3_X1   g0122(.A1(new_n322), .A2(G190), .A3(new_n312), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  AND3_X1   g0124(.A1(new_n316), .A2(new_n317), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n317), .B1(new_n316), .B2(new_n324), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n289), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT76), .ZN(new_n328));
  OAI21_X1  g0128(.A(KEYINPUT73), .B1(new_n322), .B2(new_n312), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n304), .A2(new_n291), .A3(new_n313), .ZN(new_n330));
  AOI21_X1  g0130(.A(G200), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(KEYINPUT75), .B1(new_n331), .B2(new_n323), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n316), .A2(new_n317), .A3(new_n324), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT76), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n334), .A2(new_n335), .A3(new_n289), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n244), .B1(new_n328), .B2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n288), .B1(new_n332), .B2(new_n333), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n338), .A2(KEYINPUT17), .ZN(new_n339));
  OAI21_X1  g0139(.A(KEYINPUT77), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n335), .B1(new_n334), .B2(new_n289), .ZN(new_n341));
  AOI211_X1 g0141(.A(KEYINPUT76), .B(new_n288), .C1(new_n332), .C2(new_n333), .ZN(new_n342));
  OAI21_X1  g0142(.A(KEYINPUT17), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT77), .ZN(new_n344));
  INV_X1    g0144(.A(new_n339), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G169), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(new_n314), .B2(new_n315), .ZN(new_n348));
  INV_X1    g0148(.A(G179), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n304), .A2(new_n349), .A3(new_n313), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n288), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT18), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT18), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n351), .A2(new_n354), .A3(new_n288), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT74), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT74), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n353), .A2(new_n358), .A3(new_n355), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n340), .A2(new_n346), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n279), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n260), .A2(G20), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n281), .A2(new_n364), .B1(G150), .B2(new_n248), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n203), .A2(G20), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n363), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT65), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n202), .B1(new_n207), .B2(G20), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n286), .A2(new_n369), .B1(new_n202), .B2(new_n285), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n367), .A2(KEYINPUT65), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g0173(.A(new_n373), .B(KEYINPUT9), .ZN(new_n374));
  INV_X1    g0174(.A(new_n308), .ZN(new_n375));
  INV_X1    g0175(.A(new_n311), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n375), .B1(G226), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(G222), .A2(G1698), .ZN(new_n378));
  INV_X1    g0178(.A(G1698), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n379), .A2(G223), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n258), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n381), .B(new_n303), .C1(G77), .C2(new_n258), .ZN(new_n382));
  AND2_X1   g0182(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G190), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n290), .B2(new_n383), .ZN(new_n385));
  OAI22_X1  g0185(.A1(new_n374), .A2(new_n385), .B1(KEYINPUT67), .B2(KEYINPUT10), .ZN(new_n386));
  NAND2_X1  g0186(.A1(KEYINPUT67), .A2(KEYINPUT10), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n386), .B(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n373), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n383), .A2(new_n349), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n389), .B(new_n390), .C1(G169), .C2(new_n383), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n375), .B1(G238), .B2(new_n376), .ZN(new_n393));
  NAND2_X1  g0193(.A1(G33), .A2(G97), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n309), .A2(G1698), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(G226), .B2(G1698), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n394), .B1(new_n396), .B2(new_n264), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n303), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n393), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT13), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n399), .A2(KEYINPUT13), .ZN(new_n402));
  OR2_X1    g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT14), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n403), .A2(new_n404), .A3(G169), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n401), .A2(new_n402), .ZN(new_n406));
  OAI21_X1  g0206(.A(KEYINPUT14), .B1(new_n406), .B2(new_n347), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(G179), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n405), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n248), .A2(G50), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n410), .B(KEYINPUT68), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n364), .A2(G77), .B1(G20), .B2(new_n218), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n363), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OR2_X1    g0213(.A1(new_n413), .A2(KEYINPUT11), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(KEYINPUT11), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT69), .B1(new_n284), .B2(G68), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n416), .B(KEYINPUT12), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n218), .B1(new_n207), .B2(G20), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n417), .B1(new_n286), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n414), .A2(new_n415), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n409), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n403), .A2(G200), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n420), .B1(new_n406), .B2(G190), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n281), .A2(new_n248), .B1(G20), .B2(G77), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT66), .ZN(new_n427));
  INV_X1    g0227(.A(new_n364), .ZN(new_n428));
  XNOR2_X1  g0228(.A(KEYINPUT15), .B(G87), .ZN(new_n429));
  OAI22_X1  g0229(.A1(new_n426), .A2(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n426), .A2(new_n427), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n279), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(G77), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n433), .B1(new_n207), .B2(G20), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n286), .A2(new_n434), .B1(new_n433), .B2(new_n285), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n258), .A2(new_n379), .ZN(new_n437));
  INV_X1    g0237(.A(G107), .ZN(new_n438));
  OAI22_X1  g0238(.A1(new_n437), .A2(new_n309), .B1(new_n438), .B2(new_n258), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n258), .A2(G1698), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n440), .A2(new_n219), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n303), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(G244), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n442), .B(new_n308), .C1(new_n443), .C2(new_n311), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n436), .B1(new_n347), .B2(new_n444), .ZN(new_n445));
  OR2_X1    g0245(.A1(new_n444), .A2(G179), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n444), .A2(G200), .ZN(new_n448));
  INV_X1    g0248(.A(G190), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n436), .B(new_n448), .C1(new_n449), .C2(new_n444), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n425), .A2(new_n447), .A3(new_n450), .ZN(new_n451));
  NOR3_X1   g0251(.A1(new_n392), .A2(new_n422), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n362), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT23), .B1(new_n208), .B2(G107), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT86), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT86), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n456), .B(KEYINPUT23), .C1(new_n208), .C2(G107), .ZN(new_n457));
  OR3_X1    g0257(.A1(new_n208), .A2(KEYINPUT23), .A3(G107), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n208), .A2(G33), .A3(G116), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n455), .A2(new_n457), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  XNOR2_X1  g0260(.A(new_n460), .B(KEYINPUT87), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n258), .A2(new_n208), .A3(G87), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT22), .ZN(new_n463));
  XNOR2_X1  g0263(.A(new_n462), .B(new_n463), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n461), .A2(KEYINPUT24), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT24), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT87), .ZN(new_n467));
  XNOR2_X1  g0267(.A(new_n460), .B(new_n467), .ZN(new_n468));
  XNOR2_X1  g0268(.A(new_n462), .B(KEYINPUT22), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n279), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n207), .A2(G33), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n284), .A2(new_n472), .A3(new_n278), .A4(new_n277), .ZN(new_n473));
  XNOR2_X1  g0273(.A(new_n473), .B(KEYINPUT82), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G107), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n284), .A2(G107), .ZN(new_n476));
  XNOR2_X1  g0276(.A(new_n476), .B(KEYINPUT25), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n471), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n258), .A2(G257), .A3(G1698), .ZN(new_n481));
  NAND2_X1  g0281(.A1(G33), .A2(G294), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n481), .B(new_n482), .C1(new_n437), .C2(new_n221), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n483), .A2(KEYINPUT88), .A3(new_n303), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n306), .A2(G1), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n485), .B(KEYINPUT83), .C1(KEYINPUT5), .C2(new_n305), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n207), .B(G45), .C1(new_n305), .C2(KEYINPUT5), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT83), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n305), .A2(KEYINPUT5), .ZN(new_n490));
  AND3_X1   g0290(.A1(new_n486), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(G274), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n303), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n487), .A2(new_n488), .B1(KEYINPUT5), .B2(new_n305), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n303), .B1(new_n495), .B2(new_n486), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G264), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n484), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(KEYINPUT88), .B1(new_n483), .B2(new_n303), .ZN(new_n499));
  NOR3_X1   g0299(.A1(new_n498), .A2(G190), .A3(new_n499), .ZN(new_n500));
  OR2_X1    g0300(.A1(new_n500), .A2(KEYINPUT89), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n483), .A2(new_n303), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n502), .A2(new_n497), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n494), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n500), .A2(KEYINPUT89), .B1(new_n290), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n480), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(G169), .B1(new_n498), .B2(new_n499), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n503), .A2(G179), .A3(new_n494), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n471), .A2(new_n479), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n302), .B1(G250), .B2(new_n485), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n511), .B1(new_n492), .B2(new_n485), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G116), .ZN(new_n513));
  OAI221_X1 g0313(.A(new_n513), .B1(new_n440), .B2(new_n443), .C1(new_n219), .C2(new_n437), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n512), .B1(new_n514), .B2(new_n303), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n515), .A2(G169), .ZN(new_n516));
  AOI211_X1 g0316(.A(G179), .B(new_n512), .C1(new_n514), .C2(new_n303), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT84), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT82), .ZN(new_n520));
  XNOR2_X1  g0320(.A(new_n473), .B(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n519), .B1(new_n521), .B2(new_n429), .ZN(new_n522));
  INV_X1    g0322(.A(new_n429), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n474), .A2(KEYINPUT84), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT85), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT19), .ZN(new_n527));
  XNOR2_X1  g0327(.A(KEYINPUT79), .B(G97), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n527), .B1(new_n528), .B2(new_n428), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n208), .B1(new_n394), .B2(new_n527), .ZN(new_n530));
  INV_X1    g0330(.A(G97), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(KEYINPUT79), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT79), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(G97), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n220), .A2(new_n438), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n530), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n258), .A2(new_n208), .A3(G68), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n529), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n539), .A2(new_n279), .B1(new_n285), .B2(new_n429), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n525), .A2(new_n526), .A3(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n526), .B1(new_n525), .B2(new_n540), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n518), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(KEYINPUT7), .B1(new_n264), .B2(new_n208), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n545), .B1(new_n272), .B2(new_n273), .ZN(new_n546));
  OAI21_X1  g0346(.A(KEYINPUT81), .B1(new_n546), .B2(new_n438), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n248), .A2(G77), .ZN(new_n548));
  XOR2_X1   g0348(.A(new_n548), .B(KEYINPUT78), .Z(new_n549));
  NAND4_X1  g0349(.A1(new_n535), .A2(KEYINPUT80), .A3(KEYINPUT6), .A4(new_n438), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT80), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n438), .A2(KEYINPUT6), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n551), .B1(new_n528), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n531), .A2(new_n438), .ZN(new_n554));
  NOR2_X1   g0354(.A1(G97), .A2(G107), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n550), .B(new_n553), .C1(KEYINPUT6), .C2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n549), .B1(new_n557), .B2(G20), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n274), .A2(new_n259), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT81), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n559), .A2(new_n560), .A3(G107), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n547), .A2(new_n558), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n279), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n521), .A2(G97), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n284), .A2(new_n531), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  AOI22_X1  g0367(.A1(G257), .A2(new_n496), .B1(new_n491), .B2(new_n493), .ZN(new_n568));
  NAND2_X1  g0368(.A1(G33), .A2(G283), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n258), .A2(G250), .A3(G1698), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n258), .A2(G244), .A3(new_n379), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT4), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n569), .B(new_n570), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n571), .A2(new_n572), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n303), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(G169), .B1(new_n568), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n568), .A2(new_n575), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n576), .B1(new_n578), .B2(new_n349), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n567), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n562), .A2(new_n279), .B1(new_n564), .B2(new_n565), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n577), .A2(G200), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n578), .A2(G190), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n515), .A2(new_n290), .ZN(new_n585));
  AOI211_X1 g0385(.A(new_n449), .B(new_n512), .C1(new_n514), .C2(new_n303), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n540), .B1(new_n220), .B2(new_n521), .ZN(new_n587));
  NOR3_X1   g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n544), .A2(new_n580), .A3(new_n584), .A4(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT20), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n569), .A2(new_n208), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n593), .B1(new_n535), .B2(new_n260), .ZN(new_n594));
  INV_X1    g0394(.A(G116), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n277), .A2(new_n278), .B1(G20), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n592), .B1(new_n594), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n528), .A2(G33), .ZN(new_n599));
  OAI211_X1 g0399(.A(KEYINPUT20), .B(new_n596), .C1(new_n599), .C2(new_n593), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  MUX2_X1   g0401(.A(new_n284), .B(new_n473), .S(G116), .Z(new_n602));
  AOI21_X1  g0402(.A(new_n347), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n258), .A2(G264), .A3(G1698), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n258), .A2(G257), .A3(new_n379), .ZN(new_n605));
  INV_X1    g0405(.A(G303), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n604), .B(new_n605), .C1(new_n606), .C2(new_n258), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n303), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n496), .A2(G270), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n608), .A2(new_n609), .A3(new_n494), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n603), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT21), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n603), .A2(KEYINPUT21), .A3(new_n610), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n601), .A2(new_n602), .ZN(new_n615));
  AOI22_X1  g0415(.A1(G270), .A2(new_n496), .B1(new_n491), .B2(new_n493), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n615), .A2(G179), .A3(new_n608), .A4(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n613), .A2(new_n614), .A3(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(G190), .A3(new_n608), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n615), .B1(new_n610), .B2(G200), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n510), .A2(new_n591), .A3(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n453), .A2(new_n622), .ZN(G372));
  INV_X1    g0423(.A(new_n453), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT26), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT91), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n577), .A2(new_n347), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n627), .B1(G179), .B2(new_n577), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n626), .B1(new_n628), .B2(new_n581), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n567), .A2(new_n579), .A3(KEYINPUT91), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n544), .A2(new_n589), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n625), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n543), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n541), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n588), .B1(new_n635), .B2(new_n518), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n628), .A2(new_n581), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n636), .A2(KEYINPUT92), .A3(KEYINPUT26), .A4(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n544), .A2(new_n637), .A3(KEYINPUT26), .A4(new_n589), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT92), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n633), .A2(new_n638), .A3(new_n641), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n509), .A2(KEYINPUT90), .A3(new_n618), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT90), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n507), .A2(new_n508), .ZN(new_n645));
  OAI21_X1  g0445(.A(KEYINPUT24), .B1(new_n461), .B2(new_n464), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n468), .A2(new_n466), .A3(new_n469), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n363), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n645), .B1(new_n648), .B2(new_n478), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n614), .A2(new_n617), .ZN(new_n650));
  AOI21_X1  g0450(.A(KEYINPUT21), .B1(new_n603), .B2(new_n610), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n644), .B1(new_n649), .B2(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n643), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n590), .A2(new_n506), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n642), .A2(new_n656), .A3(new_n544), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n624), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n356), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n340), .A2(new_n346), .ZN(new_n660));
  INV_X1    g0460(.A(new_n447), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n422), .B1(new_n661), .B2(new_n425), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n659), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n388), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n658), .A2(new_n391), .A3(new_n664), .ZN(G369));
  NAND3_X1  g0465(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n667));
  XOR2_X1   g0467(.A(new_n667), .B(KEYINPUT93), .Z(new_n668));
  OAI21_X1  g0468(.A(G213), .B1(new_n666), .B2(KEYINPUT27), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(G343), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n480), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n510), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT95), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n649), .B2(new_n671), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n509), .A2(KEYINPUT95), .A3(new_n672), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n672), .A2(new_n615), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n621), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n652), .B2(new_n681), .ZN(new_n683));
  XNOR2_X1  g0483(.A(KEYINPUT94), .B(G330), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n652), .A2(new_n672), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n671), .B(KEYINPUT96), .ZN(new_n689));
  AOI22_X1  g0489(.A1(new_n679), .A2(new_n688), .B1(new_n509), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n687), .A2(new_n690), .ZN(G399));
  INV_X1    g0491(.A(new_n211), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G41), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(G1), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n528), .A2(new_n220), .A3(new_n438), .A4(new_n595), .ZN(new_n696));
  OAI22_X1  g0496(.A1(new_n695), .A2(new_n696), .B1(new_n216), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  INV_X1    g0498(.A(new_n689), .ZN(new_n699));
  INV_X1    g0499(.A(new_n544), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n700), .B1(new_n654), .B2(new_n655), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n699), .B1(new_n701), .B2(new_n642), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n702), .A2(KEYINPUT29), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n509), .A2(KEYINPUT98), .A3(new_n618), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT98), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n705), .B1(new_n649), .B2(new_n652), .ZN(new_n706));
  NOR4_X1   g0506(.A1(new_n590), .A2(new_n704), .A3(new_n706), .A4(new_n506), .ZN(new_n707));
  OAI21_X1  g0507(.A(KEYINPUT26), .B1(new_n631), .B2(new_n632), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n636), .A2(new_n637), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n708), .B(new_n544), .C1(KEYINPUT26), .C2(new_n709), .ZN(new_n710));
  OAI211_X1 g0510(.A(KEYINPUT29), .B(new_n671), .C1(new_n707), .C2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n515), .A2(G179), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n712), .A2(new_n504), .A3(new_n577), .A4(new_n610), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n610), .A2(new_n349), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n715), .A2(new_n578), .A3(new_n515), .A4(new_n503), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(KEYINPUT30), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n503), .A2(new_n515), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT30), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n718), .A2(new_n719), .A3(new_n578), .A4(new_n715), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n714), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT31), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n721), .A2(new_n722), .A3(new_n689), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT97), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n722), .B1(new_n721), .B2(new_n671), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n725), .A2(new_n724), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n726), .B(new_n727), .C1(new_n622), .C2(new_n699), .ZN(new_n728));
  AOI22_X1  g0528(.A1(new_n703), .A2(new_n711), .B1(new_n684), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n698), .B1(new_n729), .B2(G1), .ZN(G364));
  INV_X1    g0530(.A(new_n685), .ZN(new_n731));
  INV_X1    g0531(.A(G13), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(G20), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n207), .B1(new_n733), .B2(G45), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n693), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n731), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(new_n684), .B2(new_n683), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n278), .B1(G20), .B2(new_n347), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n208), .A2(G179), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n741), .A2(G190), .A3(G200), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(new_n220), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G190), .A2(G200), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G159), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(KEYINPUT32), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n208), .A2(new_n349), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G200), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G190), .ZN(new_n751));
  AOI211_X1 g0551(.A(new_n743), .B(new_n748), .C1(G68), .C2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n749), .A2(new_n744), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n258), .B1(new_n753), .B2(new_n433), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n749), .A2(G190), .A3(new_n290), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n754), .B1(G58), .B2(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n741), .A2(new_n449), .A3(G200), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n747), .A2(KEYINPUT32), .B1(G107), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n750), .A2(new_n449), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n349), .A2(new_n290), .A3(G190), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  AOI22_X1  g0563(.A1(new_n761), .A2(G50), .B1(G97), .B2(new_n763), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n752), .A2(new_n757), .A3(new_n760), .A4(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(G322), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n755), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(G311), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n264), .B1(new_n753), .B2(new_n768), .ZN(new_n769));
  AOI211_X1 g0569(.A(new_n767), .B(new_n769), .C1(G329), .C2(new_n746), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n761), .A2(G326), .ZN(new_n771));
  XNOR2_X1  g0571(.A(KEYINPUT33), .B(G317), .ZN(new_n772));
  INV_X1    g0572(.A(new_n742), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n751), .A2(new_n772), .B1(new_n773), .B2(G303), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n759), .A2(G283), .B1(new_n763), .B2(G294), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n770), .A2(new_n771), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n740), .B1(new_n765), .B2(new_n776), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n736), .B(KEYINPUT99), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n692), .A2(new_n264), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G355), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(G116), .B2(new_n211), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n692), .A2(new_n258), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n216), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n783), .B1(new_n306), .B2(new_n784), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n239), .A2(new_n306), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n781), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G13), .A2(G33), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G20), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n739), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n778), .B1(new_n787), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n777), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n790), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n794), .B1(new_n683), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n738), .A2(new_n796), .ZN(G396));
  NAND2_X1  g0597(.A1(new_n661), .A2(new_n671), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n450), .B1(new_n436), .B2(new_n671), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(new_n447), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n702), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n728), .A2(new_n684), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n736), .B1(new_n802), .B2(new_n803), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n740), .A2(new_n789), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n778), .B1(G77), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n761), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n809), .A2(new_n606), .B1(new_n758), .B2(new_n220), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(G107), .B2(new_n773), .ZN(new_n811));
  INV_X1    g0611(.A(G294), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n755), .A2(new_n812), .B1(new_n745), .B2(new_n768), .ZN(new_n813));
  INV_X1    g0613(.A(new_n753), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n258), .B(new_n813), .C1(G116), .C2(new_n814), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n751), .A2(G283), .B1(G97), .B2(new_n763), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n811), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(G132), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n258), .B1(new_n745), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(G50), .B2(new_n773), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n758), .A2(new_n218), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(G58), .B2(new_n763), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n756), .A2(G143), .B1(new_n814), .B2(G159), .ZN(new_n823));
  INV_X1    g0623(.A(new_n751), .ZN(new_n824));
  INV_X1    g0624(.A(G150), .ZN(new_n825));
  INV_X1    g0625(.A(G137), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n823), .B1(new_n824), .B2(new_n825), .C1(new_n826), .C2(new_n809), .ZN(new_n827));
  XNOR2_X1  g0627(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n820), .B(new_n822), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n827), .A2(new_n828), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n817), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n808), .B1(new_n831), .B2(new_n739), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n801), .B2(new_n789), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(KEYINPUT101), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n806), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(G384));
  NAND2_X1  g0636(.A1(new_n246), .A2(G77), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n216), .A2(new_n837), .B1(G50), .B2(new_n218), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n838), .A2(G1), .A3(new_n732), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n839), .B(KEYINPUT102), .Z(new_n840));
  AOI211_X1 g0640(.A(new_n595), .B(new_n214), .C1(new_n557), .C2(KEYINPUT35), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(KEYINPUT35), .B2(new_n557), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT36), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n840), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(new_n843), .B2(new_n842), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n624), .A2(new_n703), .A3(new_n711), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n846), .A2(new_n391), .A3(new_n664), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT108), .ZN(new_n848));
  INV_X1    g0648(.A(new_n798), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(new_n702), .B2(new_n801), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT103), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n421), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n409), .A2(KEYINPUT103), .A3(new_n420), .ZN(new_n853));
  INV_X1    g0653(.A(new_n425), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n420), .A2(new_n672), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n852), .A2(new_n853), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n855), .B1(new_n854), .B2(new_n409), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT104), .B1(new_n850), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n657), .A2(new_n689), .A3(new_n801), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n798), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT104), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n863), .A2(new_n864), .A3(new_n859), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n267), .B1(new_n256), .B2(new_n266), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n268), .A2(new_n279), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n287), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n868), .A2(new_n670), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n361), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n341), .A2(new_n342), .ZN(new_n871));
  XOR2_X1   g0671(.A(new_n670), .B(KEYINPUT105), .Z(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n288), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n352), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g0674(.A(KEYINPUT106), .B(KEYINPUT37), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n868), .B1(new_n351), .B2(new_n670), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n328), .A2(new_n336), .A3(new_n878), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n871), .A2(new_n877), .B1(new_n879), .B2(KEYINPUT37), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT38), .B1(new_n870), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT38), .ZN(new_n883));
  AOI211_X1 g0683(.A(new_n883), .B(new_n880), .C1(new_n361), .C2(new_n869), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n861), .B(new_n865), .C1(new_n882), .C2(new_n884), .ZN(new_n885));
  OR2_X1    g0685(.A1(new_n659), .A2(new_n872), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n870), .A2(KEYINPUT38), .A3(new_n881), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n343), .A2(new_n345), .A3(new_n659), .ZN(new_n889));
  INV_X1    g0689(.A(new_n873), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n871), .A2(new_n877), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n876), .B1(new_n874), .B2(new_n338), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT107), .B1(new_n895), .B2(new_n883), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n889), .A2(new_n890), .B1(new_n892), .B2(new_n893), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT107), .ZN(new_n898));
  NOR3_X1   g0698(.A1(new_n897), .A2(new_n898), .A3(KEYINPUT38), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n888), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT39), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n852), .A2(new_n853), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n671), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n870), .A2(new_n881), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n883), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n907), .A2(KEYINPUT39), .A3(new_n888), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n902), .A2(new_n905), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n887), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n848), .B(new_n910), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n859), .A2(new_n801), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n622), .A2(new_n699), .ZN(new_n913));
  OR3_X1    g0713(.A1(new_n721), .A2(new_n722), .A3(new_n671), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n725), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n912), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n882), .B2(new_n884), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT40), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n912), .A2(new_n917), .A3(KEYINPUT40), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n920), .A2(new_n921), .B1(new_n900), .B2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n453), .B2(new_n916), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n924), .A2(new_n624), .A3(new_n917), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n926), .A2(new_n684), .A3(new_n927), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n911), .A2(new_n928), .B1(new_n207), .B2(new_n733), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n911), .A2(new_n928), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n845), .B1(new_n929), .B2(new_n930), .ZN(G367));
  OAI211_X1 g0731(.A(new_n580), .B(new_n584), .C1(new_n581), .C2(new_n689), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT109), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n509), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n699), .B1(new_n934), .B2(new_n580), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n580), .A2(new_n689), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n938), .A2(KEYINPUT42), .A3(new_n679), .A4(new_n688), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT42), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n679), .A2(new_n688), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n940), .B1(new_n941), .B2(new_n937), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n935), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n672), .A2(new_n587), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n636), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n544), .B2(new_n944), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n946), .A2(KEYINPUT43), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n943), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT110), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n943), .A2(KEYINPUT110), .A3(new_n947), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n946), .A2(KEYINPUT43), .ZN(new_n953));
  OR3_X1    g0753(.A1(new_n943), .A2(new_n947), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n952), .A2(KEYINPUT111), .A3(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(KEYINPUT111), .B1(new_n952), .B2(new_n954), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n956), .A2(new_n957), .B1(new_n687), .B2(new_n937), .ZN(new_n958));
  INV_X1    g0758(.A(new_n957), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n687), .A2(new_n937), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n959), .A2(new_n960), .A3(new_n955), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n693), .B(KEYINPUT41), .Z(new_n962));
  INV_X1    g0762(.A(new_n690), .ZN(new_n963));
  OAI21_X1  g0763(.A(KEYINPUT112), .B1(new_n963), .B2(new_n937), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT112), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n690), .A2(new_n938), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT45), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n964), .A2(KEYINPUT45), .A3(new_n966), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n963), .A2(KEYINPUT44), .A3(new_n937), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT44), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n690), .B2(new_n938), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n969), .A2(new_n970), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n686), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n679), .A2(new_n688), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n941), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(new_n731), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n729), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT113), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n980), .A2(KEYINPUT113), .A3(new_n729), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n969), .A2(new_n970), .A3(new_n687), .A4(new_n974), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n976), .A2(new_n983), .A3(new_n984), .A4(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n962), .B1(new_n986), .B2(new_n729), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n958), .B(new_n961), .C1(new_n987), .C2(new_n735), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n791), .B1(new_n211), .B2(new_n429), .C1(new_n783), .C2(new_n235), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n778), .A2(new_n989), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n761), .A2(G311), .B1(G107), .B2(new_n763), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n991), .B1(new_n812), .B2(new_n824), .C1(new_n528), .C2(new_n758), .ZN(new_n992));
  AOI22_X1  g0792(.A1(G283), .A2(new_n814), .B1(new_n746), .B2(G317), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n258), .B1(new_n756), .B2(G303), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n773), .A2(KEYINPUT46), .A3(G116), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT46), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n742), .B2(new_n595), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n993), .A2(new_n994), .A3(new_n995), .A4(new_n997), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n753), .A2(new_n202), .B1(new_n745), .B2(new_n826), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(G150), .B2(new_n756), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n751), .A2(G159), .B1(new_n761), .B2(G143), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n773), .A2(G58), .B1(new_n763), .B2(G68), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n258), .B1(new_n758), .B2(new_n433), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT114), .Z(new_n1005));
  OAI22_X1  g0805(.A1(new_n992), .A2(new_n998), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT47), .Z(new_n1007));
  OAI221_X1 g0807(.A(new_n990), .B1(new_n740), .B2(new_n1007), .C1(new_n946), .C2(new_n795), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n988), .A2(new_n1008), .ZN(G387));
  NAND2_X1  g0809(.A1(new_n680), .A2(new_n790), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n281), .A2(new_n202), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT50), .Z(new_n1012));
  AOI211_X1 g0812(.A(G45), .B(new_n696), .C1(G68), .C2(G77), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n783), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n306), .B2(new_n232), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n779), .A2(new_n696), .B1(new_n438), .B2(new_n692), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1015), .A2(KEYINPUT115), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n791), .ZN(new_n1018));
  AOI21_X1  g0818(.A(KEYINPUT115), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n778), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n755), .A2(new_n202), .B1(new_n745), .B2(new_n825), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n264), .B(new_n1021), .C1(G68), .C2(new_n814), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n773), .A2(G77), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n751), .A2(new_n281), .B1(new_n759), .B2(G97), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n761), .A2(G159), .B1(new_n523), .B2(new_n763), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n756), .A2(G317), .B1(new_n814), .B2(G303), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(new_n824), .B2(new_n768), .C1(new_n766), .C2(new_n809), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT48), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(G283), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n763), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1030), .B1(new_n1031), .B2(new_n1032), .C1(new_n812), .C2(new_n742), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(KEYINPUT49), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n758), .A2(new_n595), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n258), .B(new_n1037), .C1(G326), .C2(new_n746), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1035), .A2(KEYINPUT49), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1026), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1020), .B1(new_n1041), .B2(new_n739), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n980), .A2(new_n735), .B1(new_n1010), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n983), .A2(new_n984), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n693), .B1(new_n980), .B2(new_n729), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1043), .B1(new_n1045), .B2(new_n1046), .ZN(G393));
  NAND2_X1  g0847(.A1(new_n976), .A2(new_n985), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n1044), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1049), .A2(new_n693), .A3(new_n986), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n976), .A2(new_n735), .A3(new_n985), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n791), .B1(new_n211), .B2(new_n528), .C1(new_n783), .C2(new_n242), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n778), .A2(new_n1052), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n824), .A2(new_n606), .B1(new_n595), .B2(new_n1032), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n264), .B1(new_n745), .B2(new_n766), .C1(new_n812), .C2(new_n753), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n438), .A2(new_n758), .B1(new_n742), .B2(new_n1031), .ZN(new_n1056));
  OR3_X1    g0856(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G317), .A2(new_n761), .B1(new_n756), .B2(G311), .ZN(new_n1058));
  XOR2_X1   g0858(.A(KEYINPUT116), .B(KEYINPUT52), .Z(new_n1059));
  XNOR2_X1  g0859(.A(new_n1058), .B(new_n1059), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G150), .A2(new_n761), .B1(new_n756), .B2(G159), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT51), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n751), .A2(G50), .B1(new_n759), .B2(G87), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n814), .A2(new_n281), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n264), .B1(new_n746), .B2(G143), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n773), .A2(G68), .B1(new_n763), .B2(G77), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n1057), .A2(new_n1060), .B1(new_n1062), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1053), .B1(new_n1068), .B2(new_n739), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n938), .B2(new_n795), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n1051), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1050), .A2(new_n1071), .ZN(G390));
  OAI21_X1  g0872(.A(new_n904), .B1(new_n850), .B2(new_n860), .ZN(new_n1073));
  NOR3_X1   g0873(.A1(new_n882), .A2(new_n884), .A3(new_n901), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n898), .B1(new_n897), .B2(KEYINPUT38), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n328), .A2(new_n336), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n339), .B1(new_n1076), .B2(KEYINPUT17), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n873), .B1(new_n1077), .B2(new_n659), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n892), .A2(new_n893), .ZN(new_n1079));
  OAI211_X1 g0879(.A(KEYINPUT107), .B(new_n883), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1075), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(KEYINPUT39), .B1(new_n1081), .B2(new_n888), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1073), .B1(new_n1074), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n880), .B1(new_n361), .B2(new_n869), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n1075), .A2(new_n1080), .B1(new_n1084), .B2(KEYINPUT38), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1085), .A2(new_n905), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n671), .B(new_n800), .C1(new_n707), .C2(new_n710), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n798), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT117), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n860), .A2(KEYINPUT118), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT118), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n859), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1089), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1086), .A2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n728), .A2(new_n684), .A3(new_n801), .A4(new_n859), .ZN(new_n1096));
  AND3_X1   g0896(.A1(new_n1083), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n912), .A2(new_n917), .A3(G330), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n1083), .B2(new_n1095), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n908), .B1(KEYINPUT39), .B2(new_n1085), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n788), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n778), .B1(new_n281), .B2(new_n807), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n742), .A2(new_n825), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT53), .ZN(new_n1105));
  INV_X1    g0905(.A(G125), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n755), .A2(new_n818), .B1(new_n745), .B2(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(KEYINPUT54), .B(G143), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n258), .B1(new_n753), .B2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n751), .A2(G137), .B1(G159), .B2(new_n763), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n761), .A2(G128), .B1(new_n759), .B2(G50), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1105), .A2(new_n1110), .A3(new_n1111), .A4(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n743), .A2(new_n258), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT120), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n753), .A2(new_n528), .B1(new_n745), .B2(new_n812), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(G116), .B2(new_n756), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n751), .A2(G107), .B1(new_n761), .B2(G283), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n821), .B1(G77), .B2(new_n763), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1113), .B1(new_n1115), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1103), .B1(new_n1121), .B2(new_n739), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n1100), .A2(new_n735), .B1(new_n1102), .B2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1083), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1101), .A2(new_n1073), .B1(new_n1086), .B2(new_n1094), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1124), .B1(new_n1125), .B2(new_n1098), .ZN(new_n1126));
  OAI211_X1 g0926(.A(G330), .B(new_n801), .C1(new_n913), .C2(new_n915), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1090), .A2(new_n1092), .A3(new_n1127), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n1128), .A2(new_n1096), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT117), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1088), .B(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n728), .A2(new_n684), .A3(new_n801), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n860), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n1098), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1129), .A2(new_n1131), .B1(new_n1134), .B2(new_n863), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n362), .A2(new_n452), .A3(new_n917), .A4(G330), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n846), .A2(new_n1137), .A3(new_n391), .A4(new_n664), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n694), .B1(new_n1126), .B2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1124), .B(new_n1142), .C1(new_n1125), .C2(new_n1098), .ZN(new_n1143));
  AOI21_X1  g0943(.A(KEYINPUT119), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1140), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1145));
  AND4_X1   g0945(.A1(KEYINPUT119), .A2(new_n1145), .A3(new_n693), .A4(new_n1143), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1123), .B1(new_n1144), .B2(new_n1146), .ZN(G378));
  NAND2_X1  g0947(.A1(new_n924), .A2(G330), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n389), .A2(new_n670), .ZN(new_n1149));
  XOR2_X1   g0949(.A(new_n1149), .B(KEYINPUT121), .Z(new_n1150));
  XNOR2_X1  g0950(.A(new_n392), .B(new_n1150), .ZN(new_n1151));
  XOR2_X1   g0951(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1152));
  XNOR2_X1  g0952(.A(new_n1151), .B(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1148), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n924), .A2(new_n1153), .A3(G330), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT123), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(new_n910), .B2(KEYINPUT122), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT122), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1160), .B(KEYINPUT123), .C1(new_n887), .C2(new_n909), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1157), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n924), .A2(G330), .A3(new_n1153), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1153), .B1(new_n924), .B2(G330), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n885), .A2(new_n886), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1074), .A2(new_n1082), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1166), .B1(new_n1167), .B2(new_n905), .ZN(new_n1168));
  OAI21_X1  g0968(.A(KEYINPUT123), .B1(new_n1168), .B2(new_n1160), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n910), .A2(KEYINPUT122), .A3(new_n1158), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1165), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1143), .A2(new_n1139), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1162), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT57), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NOR3_X1   g0975(.A1(new_n1163), .A2(new_n1164), .A3(new_n1168), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n910), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1174), .B1(new_n1143), .B2(new_n1139), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n694), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1175), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1162), .A2(new_n1171), .A3(new_n735), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n736), .B1(G50), .B2(new_n807), .ZN(new_n1183));
  INV_X1    g0983(.A(G58), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n809), .A2(new_n595), .B1(new_n758), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G97), .B2(new_n751), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n264), .A2(new_n305), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(G283), .B2(new_n746), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n756), .A2(G107), .B1(new_n814), .B2(new_n523), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n773), .A2(G77), .B1(new_n763), .B2(G68), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1186), .A2(new_n1188), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT58), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1187), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n1106), .A2(new_n809), .B1(new_n824), .B2(new_n818), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n756), .A2(G128), .B1(new_n814), .B2(G137), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n742), .B2(new_n1108), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1196), .B(new_n1198), .C1(G150), .C2(new_n763), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n759), .A2(G159), .ZN(new_n1202));
  AOI211_X1 g1002(.A(G33), .B(G41), .C1(new_n746), .C2(G124), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1195), .B1(new_n1192), .B2(new_n1191), .C1(new_n1204), .C2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1183), .B1(new_n1206), .B2(new_n739), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n1153), .B2(new_n789), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1182), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1181), .A2(new_n1210), .ZN(G375));
  NOR2_X1   g1011(.A1(new_n1093), .A2(new_n789), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n761), .A2(G294), .B1(new_n814), .B2(G107), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n595), .B2(new_n824), .ZN(new_n1214));
  XOR2_X1   g1014(.A(new_n1214), .B(KEYINPUT124), .Z(new_n1215));
  OAI22_X1  g1015(.A1(new_n1032), .A2(new_n429), .B1(new_n758), .B2(new_n433), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n264), .B1(new_n745), .B2(new_n606), .C1(new_n755), .C2(new_n1031), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1216), .B(new_n1217), .C1(G97), .C2(new_n773), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n773), .A2(G159), .B1(new_n746), .B2(G128), .ZN(new_n1219));
  XOR2_X1   g1019(.A(new_n1219), .B(KEYINPUT125), .Z(new_n1220));
  OAI22_X1  g1020(.A1(new_n818), .A2(new_n809), .B1(new_n824), .B2(new_n1108), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n258), .B1(new_n753), .B2(new_n825), .C1(new_n826), .C2(new_n755), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n1032), .A2(new_n202), .B1(new_n758), .B2(new_n1184), .ZN(new_n1223));
  NOR3_X1   g1023(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1215), .A2(new_n1218), .B1(new_n1220), .B2(new_n1224), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n778), .B1(G68), .B2(new_n807), .C1(new_n1225), .C2(new_n740), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1212), .A2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n1136), .B2(new_n735), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1142), .A2(new_n962), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1228), .B1(new_n1229), .B2(new_n1231), .ZN(G381));
  OR2_X1    g1032(.A1(G393), .A2(G396), .ZN(new_n1233));
  OR4_X1    g1033(.A1(G384), .A2(new_n1233), .A3(G390), .A4(G381), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1234), .A2(G387), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1209), .B1(new_n1175), .B2(new_n1180), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1145), .A2(new_n693), .A3(new_n1143), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1123), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT126), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1123), .A2(new_n1237), .A3(KEYINPUT126), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1235), .A2(new_n1236), .A3(new_n1242), .ZN(G407));
  INV_X1    g1043(.A(G213), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1244), .A2(G343), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1236), .A2(new_n1242), .A3(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(G407), .A2(G213), .A3(new_n1246), .ZN(G409));
  XOR2_X1   g1047(.A(G393), .B(G396), .Z(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n988), .A2(new_n1008), .A3(G390), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(G390), .B1(new_n988), .B2(new_n1008), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1249), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(G390), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(G387), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1255), .A2(new_n1248), .A3(new_n1250), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1253), .A2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1231), .B1(KEYINPUT60), .B2(new_n1140), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1135), .A2(new_n1138), .A3(KEYINPUT60), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n693), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1228), .B1(new_n1258), .B2(new_n1260), .ZN(new_n1261));
  AND2_X1   g1061(.A1(new_n1261), .A2(new_n835), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1261), .A2(new_n835), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1245), .A2(G2897), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1264), .B(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1176), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1177), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1268), .A2(new_n1269), .A3(new_n735), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1208), .B(new_n1270), .C1(new_n1173), .C2(new_n962), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n1236), .A2(G378), .B1(new_n1242), .B2(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1267), .B1(new_n1272), .B2(new_n1245), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1181), .A2(G378), .A3(new_n1210), .ZN(new_n1274));
  AOI21_X1  g1074(.A(KEYINPUT126), .B1(new_n1123), .B2(new_n1237), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1241), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1271), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1274), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT62), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1245), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1278), .A2(new_n1279), .A3(new_n1280), .A4(new_n1264), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT61), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1273), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1245), .B1(new_n1274), .B2(new_n1277), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1279), .B1(new_n1284), .B2(new_n1264), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1257), .B1(new_n1283), .B2(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1253), .A2(new_n1282), .A3(new_n1256), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT127), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(new_n1287), .B(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1284), .A2(new_n1264), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT63), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1284), .A2(KEYINPUT63), .A3(new_n1264), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1289), .A2(new_n1292), .A3(new_n1273), .A4(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1286), .A2(new_n1294), .ZN(G405));
  NAND2_X1  g1095(.A1(G375), .A2(new_n1242), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1274), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1264), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1296), .B(new_n1274), .C1(new_n1262), .C2(new_n1263), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  XNOR2_X1  g1100(.A(new_n1300), .B(new_n1257), .ZN(G402));
endmodule


