//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 1 0 0 0 0 0 0 0 1 0 0 0 1 1 0 1 1 1 0 1 0 1 0 1 1 1 0 0 0 0 1 1 0 1 1 1 0 1 0 1 1 1 1 1 1 0 0 1 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n574, new_n575, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n641, new_n642, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1226,
    new_n1227, new_n1228, new_n1229;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT66), .Z(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G125), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT67), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n465), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n463), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n475), .B1(new_n472), .B2(new_n473), .ZN(new_n476));
  OAI21_X1  g051(.A(G2105), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n464), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n478), .A2(new_n467), .ZN(new_n479));
  INV_X1    g054(.A(G2105), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT69), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n465), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n479), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n466), .A2(G2105), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT70), .ZN(new_n486));
  AOI22_X1  g061(.A1(new_n484), .A2(G137), .B1(G101), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n477), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G160));
  NAND2_X1  g064(.A1(new_n484), .A2(G136), .ZN(new_n490));
  XOR2_X1   g065(.A(new_n490), .B(KEYINPUT71), .Z(new_n491));
  OR2_X1    g066(.A1(G100), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G112), .C2(new_n480), .ZN(new_n493));
  XOR2_X1   g068(.A(new_n493), .B(KEYINPUT72), .Z(new_n494));
  NAND3_X1  g069(.A1(new_n479), .A2(G2105), .A3(new_n482), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n494), .B1(G124), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n491), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g073(.A(new_n498), .B(KEYINPUT73), .ZN(G162));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G114), .ZN(new_n502));
  AND3_X1   g077(.A1(new_n502), .A2(KEYINPUT74), .A3(G2105), .ZN(new_n503));
  AOI21_X1  g078(.A(KEYINPUT74), .B1(new_n502), .B2(G2105), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n501), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G126), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n495), .B2(new_n506), .ZN(new_n507));
  AND2_X1   g082(.A1(new_n480), .A2(G138), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n479), .A2(new_n482), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT4), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n469), .A2(new_n471), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT4), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n511), .A2(new_n512), .A3(new_n508), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n507), .B1(new_n510), .B2(new_n513), .ZN(G164));
  AND2_X1   g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  AND2_X1   g093(.A1(new_n518), .A2(G62), .ZN(new_n519));
  NAND2_X1  g094(.A1(G75), .A2(G543), .ZN(new_n520));
  XOR2_X1   g095(.A(new_n520), .B(KEYINPUT78), .Z(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  OAI21_X1  g097(.A(G651), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G50), .ZN(new_n524));
  AND2_X1   g099(.A1(KEYINPUT75), .A2(KEYINPUT6), .ZN(new_n525));
  NOR2_X1   g100(.A1(KEYINPUT75), .A2(KEYINPUT6), .ZN(new_n526));
  OAI21_X1  g101(.A(G651), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(KEYINPUT76), .ZN(new_n528));
  INV_X1    g103(.A(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(KEYINPUT6), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT76), .ZN(new_n531));
  OAI211_X1 g106(.A(new_n531), .B(G651), .C1(new_n525), .C2(new_n526), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n528), .A2(G543), .A3(new_n530), .A4(new_n532), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n528), .A2(new_n518), .A3(new_n530), .A4(new_n532), .ZN(new_n534));
  INV_X1    g109(.A(G88), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n524), .A2(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n536), .A2(KEYINPUT77), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n536), .A2(KEYINPUT77), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n523), .B1(new_n537), .B2(new_n538), .ZN(G303));
  INV_X1    g114(.A(G303), .ZN(G166));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT79), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT7), .ZN(new_n543));
  AND2_X1   g118(.A1(G63), .A2(G651), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n543), .B1(new_n518), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n532), .A2(new_n530), .ZN(new_n546));
  OR2_X1    g121(.A1(KEYINPUT75), .A2(KEYINPUT6), .ZN(new_n547));
  NAND2_X1  g122(.A1(KEYINPUT75), .A2(KEYINPUT6), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n531), .B1(new_n549), .B2(G651), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n551), .A2(G89), .A3(new_n518), .ZN(new_n552));
  INV_X1    g127(.A(new_n533), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G51), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n545), .A2(new_n552), .A3(new_n554), .ZN(G286));
  INV_X1    g130(.A(G286), .ZN(G168));
  INV_X1    g131(.A(G52), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n558));
  OAI22_X1  g133(.A1(new_n533), .A2(new_n557), .B1(new_n558), .B2(new_n529), .ZN(new_n559));
  INV_X1    g134(.A(G90), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n534), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n559), .A2(new_n561), .ZN(G171));
  NAND2_X1  g137(.A1(G68), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G56), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n517), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G651), .ZN(new_n566));
  INV_X1    g141(.A(G43), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n533), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(G81), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n534), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G860), .ZN(G153));
  NAND4_X1  g147(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g148(.A1(G1), .A2(G3), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT8), .ZN(new_n575));
  NAND4_X1  g150(.A1(G319), .A2(G483), .A3(G661), .A4(new_n575), .ZN(G188));
  INV_X1    g151(.A(KEYINPUT80), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n551), .A2(new_n577), .A3(G53), .A4(G543), .ZN(new_n578));
  INV_X1    g153(.A(G53), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT80), .B1(new_n533), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n580), .A3(KEYINPUT9), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n518), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n582), .A2(new_n529), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT81), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n534), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n530), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n529), .B1(new_n547), .B2(new_n548), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n586), .B1(new_n587), .B2(new_n531), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n588), .A2(KEYINPUT81), .A3(new_n518), .A4(new_n528), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n585), .A2(G91), .A3(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT9), .ZN(new_n591));
  OAI211_X1 g166(.A(KEYINPUT80), .B(new_n591), .C1(new_n533), .C2(new_n579), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n581), .A2(new_n583), .A3(new_n590), .A4(new_n592), .ZN(G299));
  INV_X1    g168(.A(G171), .ZN(G301));
  NAND2_X1  g169(.A1(new_n585), .A2(new_n589), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(G87), .ZN(new_n597));
  INV_X1    g172(.A(G74), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n529), .B1(new_n517), .B2(new_n598), .ZN(new_n599));
  AND2_X1   g174(.A1(G49), .A2(G543), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n551), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT82), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n551), .A2(KEYINPUT82), .A3(new_n600), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n599), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n597), .A2(new_n605), .ZN(G288));
  NAND2_X1  g181(.A1(new_n553), .A2(G48), .ZN(new_n607));
  INV_X1    g182(.A(G61), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n517), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT83), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(G73), .A2(G543), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(new_n609), .B2(new_n610), .ZN(new_n614));
  OAI21_X1  g189(.A(G651), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n607), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(new_n596), .B2(G86), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(G305));
  INV_X1    g193(.A(G47), .ZN(new_n619));
  INV_X1    g194(.A(G85), .ZN(new_n620));
  OAI22_X1  g195(.A1(new_n619), .A2(new_n533), .B1(new_n534), .B2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT84), .ZN(new_n622));
  AND2_X1   g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  AOI22_X1  g199(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n625));
  OAI22_X1  g200(.A1(new_n623), .A2(new_n624), .B1(new_n529), .B2(new_n625), .ZN(G290));
  NAND2_X1  g201(.A1(G301), .A2(G868), .ZN(new_n627));
  NAND2_X1  g202(.A1(G79), .A2(G543), .ZN(new_n628));
  INV_X1    g203(.A(G66), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n517), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(G651), .ZN(new_n631));
  INV_X1    g206(.A(G54), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(new_n533), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n585), .A2(G92), .A3(new_n589), .ZN(new_n634));
  INV_X1    g209(.A(KEYINPUT10), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g211(.A1(new_n585), .A2(new_n589), .A3(KEYINPUT10), .A4(G92), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n633), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n627), .B1(new_n638), .B2(G868), .ZN(G284));
  OAI21_X1  g214(.A(new_n627), .B1(new_n638), .B2(G868), .ZN(G321));
  NAND2_X1  g215(.A1(G286), .A2(G868), .ZN(new_n641));
  AND4_X1   g216(.A1(new_n581), .A2(new_n583), .A3(new_n590), .A4(new_n592), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n641), .B1(new_n642), .B2(G868), .ZN(G297));
  OAI21_X1  g218(.A(new_n641), .B1(new_n642), .B2(G868), .ZN(G280));
  INV_X1    g219(.A(G559), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n638), .B1(new_n645), .B2(G860), .ZN(G148));
  NAND2_X1  g221(.A1(new_n636), .A2(new_n637), .ZN(new_n647));
  INV_X1    g222(.A(new_n633), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(KEYINPUT85), .B1(new_n649), .B2(G559), .ZN(new_n650));
  INV_X1    g225(.A(KEYINPUT85), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n638), .A2(new_n651), .A3(new_n645), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(G868), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n654), .A2(KEYINPUT86), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(KEYINPUT86), .ZN(new_n656));
  OAI211_X1 g231(.A(new_n655), .B(new_n656), .C1(G868), .C2(new_n571), .ZN(G323));
  XNOR2_X1  g232(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g233(.A1(new_n511), .A2(new_n486), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT12), .Z(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT13), .Z(new_n661));
  INV_X1    g236(.A(G2100), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  OR2_X1    g239(.A1(G99), .A2(G2105), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n665), .B(G2104), .C1(G111), .C2(new_n480), .ZN(new_n666));
  INV_X1    g241(.A(G123), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n666), .B1(new_n495), .B2(new_n667), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n668), .B1(G135), .B2(new_n484), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(G2096), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n663), .A2(new_n664), .A3(new_n670), .ZN(G156));
  XOR2_X1   g246(.A(G2451), .B(G2454), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT16), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1341), .B(G1348), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT14), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2427), .B(G2438), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2430), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT15), .B(G2435), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n676), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(new_n679), .B2(new_n678), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n675), .B(new_n681), .Z(new_n682));
  XNOR2_X1  g257(.A(G2443), .B(G2446), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  AND3_X1   g260(.A1(new_n684), .A2(G14), .A3(new_n685), .ZN(G401));
  XOR2_X1   g261(.A(KEYINPUT87), .B(KEYINPUT18), .Z(new_n687));
  XOR2_X1   g262(.A(G2084), .B(G2090), .Z(new_n688));
  XNOR2_X1  g263(.A(G2067), .B(G2678), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(KEYINPUT17), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n688), .A2(new_n689), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n687), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G2072), .B(G2078), .Z(new_n694));
  INV_X1    g269(.A(new_n687), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n694), .B1(new_n690), .B2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n693), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G2096), .B(G2100), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(G227));
  XOR2_X1   g274(.A(G1961), .B(G1966), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT88), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1956), .B(G2474), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1971), .B(G1976), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT19), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT20), .Z(new_n708));
  NOR2_X1   g283(.A1(new_n701), .A2(new_n703), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n710), .A2(new_n706), .A3(new_n704), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n708), .B(new_n711), .C1(new_n706), .C2(new_n710), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(G1991), .B(G1996), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(G1981), .B(G1986), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(G229));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G20), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT23), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(new_n642), .B2(new_n719), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT102), .B(G1956), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT89), .B(G29), .Z(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n726), .A2(G35), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G162), .B2(new_n726), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT29), .ZN(new_n729));
  AND3_X1   g304(.A1(new_n729), .A2(KEYINPUT101), .A3(G2090), .ZN(new_n730));
  AOI21_X1  g305(.A(KEYINPUT101), .B1(new_n729), .B2(G2090), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n724), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n732), .A2(KEYINPUT103), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(KEYINPUT103), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n719), .A2(G19), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT93), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n571), .B2(new_n719), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT94), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(G1341), .Z(new_n739));
  INV_X1    g314(.A(G1348), .ZN(new_n740));
  NOR2_X1   g315(.A1(G4), .A2(G16), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n638), .B2(G16), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n739), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  OAI221_X1 g319(.A(new_n744), .B1(new_n740), .B2(new_n743), .C1(new_n729), .C2(G2090), .ZN(new_n745));
  INV_X1    g320(.A(G29), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n746), .A2(G33), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n511), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(new_n480), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n480), .A2(G103), .A3(G2104), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT25), .Z(new_n751));
  INV_X1    g326(.A(G139), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n751), .B1(new_n483), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT95), .Z(new_n755));
  AOI21_X1  g330(.A(new_n747), .B1(new_n755), .B2(G29), .ZN(new_n756));
  INV_X1    g331(.A(G2072), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(G168), .A2(new_n719), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n719), .B2(G21), .ZN(new_n760));
  INV_X1    g335(.A(G1966), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n719), .A2(G5), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G171), .B2(new_n719), .ZN(new_n763));
  OAI22_X1  g338(.A1(new_n760), .A2(new_n761), .B1(G1961), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n746), .A2(G32), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n496), .A2(G129), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT98), .Z(new_n767));
  NAND3_X1  g342(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT26), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n486), .A2(G105), .ZN(new_n770));
  AOI211_X1 g345(.A(new_n769), .B(new_n770), .C1(G141), .C2(new_n484), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n767), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n765), .B1(new_n772), .B2(new_n746), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT27), .B(G1996), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n669), .A2(new_n726), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT31), .B(G11), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT30), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(G28), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT99), .Z(new_n781));
  OAI211_X1 g356(.A(new_n781), .B(new_n746), .C1(new_n779), .C2(G28), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n777), .A2(new_n778), .A3(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT100), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n725), .A2(G26), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT28), .ZN(new_n786));
  OR2_X1    g361(.A1(G104), .A2(G2105), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n787), .B(G2104), .C1(G116), .C2(new_n480), .ZN(new_n788));
  INV_X1    g363(.A(G128), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(new_n495), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G140), .B2(new_n484), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n786), .B1(new_n791), .B2(new_n746), .ZN(new_n792));
  INV_X1    g367(.A(G2067), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n776), .A2(new_n784), .A3(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(G34), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT96), .B(KEYINPUT24), .Z(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n726), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  OAI22_X1  g375(.A1(new_n800), .A2(KEYINPUT97), .B1(new_n796), .B2(new_n798), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(KEYINPUT97), .B2(new_n800), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G160), .B2(G29), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n803), .A2(G2084), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n726), .A2(G27), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G164), .B2(new_n726), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(G2078), .Z(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n773), .B2(new_n775), .ZN(new_n808));
  NOR3_X1   g383(.A1(new_n795), .A2(new_n804), .A3(new_n808), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n756), .A2(new_n757), .B1(G1961), .B2(new_n763), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n760), .A2(new_n761), .B1(G2084), .B2(new_n803), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  NOR4_X1   g387(.A1(new_n745), .A2(new_n758), .A3(new_n764), .A4(new_n812), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n733), .A2(new_n734), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n719), .A2(G6), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n617), .B2(new_n719), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT91), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT32), .B(G1981), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n719), .A2(G22), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G166), .B2(new_n719), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(G1971), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n719), .A2(G23), .ZN(new_n823));
  INV_X1    g398(.A(G288), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n824), .B2(new_n719), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT33), .B(G1976), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n822), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n819), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(KEYINPUT92), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT92), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n819), .A2(new_n828), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(KEYINPUT34), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  OR2_X1    g408(.A1(G16), .A2(G24), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(G290), .B2(new_n719), .ZN(new_n835));
  INV_X1    g410(.A(G1986), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n836), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n726), .A2(G25), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n484), .A2(G131), .ZN(new_n841));
  INV_X1    g416(.A(G119), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n480), .A2(G107), .ZN(new_n843));
  OAI21_X1  g418(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n844));
  OAI22_X1  g419(.A1(new_n495), .A2(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n840), .B1(new_n846), .B2(new_n726), .ZN(new_n847));
  XNOR2_X1  g422(.A(KEYINPUT35), .B(G1991), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT90), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n847), .B(new_n849), .Z(new_n850));
  OR2_X1    g425(.A1(new_n839), .A2(new_n850), .ZN(new_n851));
  NOR3_X1   g426(.A1(new_n833), .A2(new_n837), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n830), .A2(KEYINPUT34), .A3(new_n832), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(KEYINPUT36), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT36), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n852), .A2(new_n856), .A3(new_n853), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n814), .B1(new_n855), .B2(new_n857), .ZN(G311));
  NAND2_X1  g433(.A1(new_n855), .A2(new_n857), .ZN(new_n859));
  INV_X1    g434(.A(new_n814), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(G150));
  NAND2_X1  g436(.A1(new_n638), .A2(G559), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT38), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n568), .A2(new_n570), .ZN(new_n864));
  NAND2_X1  g439(.A1(G80), .A2(G543), .ZN(new_n865));
  INV_X1    g440(.A(G67), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n865), .B1(new_n517), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(G651), .ZN(new_n868));
  INV_X1    g443(.A(G93), .ZN(new_n869));
  INV_X1    g444(.A(G55), .ZN(new_n870));
  OAI221_X1 g445(.A(new_n868), .B1(new_n534), .B2(new_n869), .C1(new_n870), .C2(new_n533), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n864), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n868), .B1(new_n533), .B2(new_n870), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n534), .A2(new_n869), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n571), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n863), .B(new_n878), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n879), .A2(KEYINPUT39), .ZN(new_n880));
  INV_X1    g455(.A(G860), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(KEYINPUT39), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n875), .A2(new_n881), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT37), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(G145));
  XNOR2_X1  g461(.A(new_n755), .B(new_n772), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n496), .A2(G130), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n480), .A2(G118), .ZN(new_n889));
  OAI21_X1  g464(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n891), .B1(G142), .B2(new_n484), .ZN(new_n892));
  XOR2_X1   g467(.A(new_n892), .B(new_n660), .Z(new_n893));
  XNOR2_X1  g468(.A(new_n887), .B(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(G140), .ZN(new_n895));
  OAI221_X1 g470(.A(new_n788), .B1(new_n483), .B2(new_n895), .C1(new_n789), .C2(new_n495), .ZN(new_n896));
  XNOR2_X1  g471(.A(G164), .B(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(new_n846), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n894), .B(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n488), .B(new_n669), .ZN(new_n900));
  XNOR2_X1  g475(.A(G162), .B(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(G37), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n899), .A2(new_n901), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT40), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n906), .B(new_n907), .ZN(G395));
  AND3_X1   g483(.A1(new_n650), .A2(new_n652), .A3(new_n878), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n878), .B1(new_n650), .B2(new_n652), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n649), .A2(G299), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n642), .A2(new_n638), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(KEYINPUT106), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT104), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(new_n914), .B2(KEYINPUT41), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n638), .B(G299), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT41), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(KEYINPUT104), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT105), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n922), .B1(new_n918), .B2(new_n919), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n914), .A2(KEYINPUT105), .A3(KEYINPUT41), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n921), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n915), .B1(new_n911), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n925), .A2(new_n927), .A3(new_n911), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT42), .B1(new_n926), .B2(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(G303), .B(G288), .ZN(new_n931));
  NAND2_X1  g506(.A1(G290), .A2(new_n617), .ZN(new_n932));
  OR2_X1    g507(.A1(G290), .A2(new_n617), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n925), .A2(new_n911), .ZN(new_n937));
  OR2_X1    g512(.A1(new_n909), .A2(new_n910), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n927), .B1(new_n938), .B2(new_n918), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT42), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(new_n941), .A3(new_n928), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n930), .A2(new_n936), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n936), .B1(new_n930), .B2(new_n942), .ZN(new_n944));
  OAI21_X1  g519(.A(G868), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n875), .A2(G868), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n945), .A2(new_n947), .ZN(G295));
  INV_X1    g523(.A(G868), .ZN(new_n949));
  OR2_X1    g524(.A1(new_n934), .A2(new_n935), .ZN(new_n950));
  INV_X1    g525(.A(new_n942), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n941), .B1(new_n940), .B2(new_n928), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n930), .A2(new_n936), .A3(new_n942), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n949), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT107), .B1(new_n955), .B2(new_n946), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n945), .A2(new_n957), .A3(new_n947), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n956), .A2(new_n958), .ZN(G331));
  INV_X1    g534(.A(KEYINPUT108), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n960), .B1(new_n559), .B2(new_n561), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n961), .B1(new_n872), .B2(new_n876), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(G286), .B1(KEYINPUT108), .B2(G171), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n872), .A2(new_n876), .A3(new_n961), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(G168), .B1(new_n960), .B2(G301), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n872), .A2(new_n876), .A3(new_n961), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n967), .B1(new_n968), .B2(new_n962), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT105), .B1(new_n914), .B2(KEYINPUT41), .ZN(new_n972));
  AOI211_X1 g547(.A(new_n922), .B(new_n919), .C1(new_n912), .C2(new_n913), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n971), .B1(new_n974), .B2(new_n921), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n966), .A2(new_n969), .A3(new_n918), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n936), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT104), .B1(new_n918), .B2(new_n919), .ZN(new_n979));
  AND4_X1   g554(.A1(KEYINPUT104), .A2(new_n912), .A3(new_n919), .A4(new_n913), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n923), .A2(new_n924), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n970), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n983), .A2(new_n950), .A3(new_n976), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n978), .A2(new_n984), .A3(new_n903), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT43), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n914), .A2(KEYINPUT41), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n919), .B1(new_n912), .B2(new_n913), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n970), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n976), .ZN(new_n990));
  AOI21_X1  g565(.A(G37), .B1(new_n990), .B2(new_n936), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n984), .A2(new_n986), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT109), .ZN(new_n993));
  AOI22_X1  g568(.A1(KEYINPUT43), .A2(new_n985), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n984), .A2(new_n991), .A3(KEYINPUT109), .A4(new_n986), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT44), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT44), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n985), .A2(new_n986), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n984), .A2(KEYINPUT43), .A3(new_n991), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n996), .A2(KEYINPUT110), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n985), .A2(KEYINPUT43), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n992), .A2(new_n993), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1003), .A2(new_n1004), .A3(new_n995), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n997), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n998), .A2(new_n999), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT44), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1002), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1001), .A2(new_n1009), .ZN(G397));
  NAND2_X1  g585(.A1(new_n791), .A2(new_n793), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n896), .A2(G2067), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g588(.A(new_n1013), .B(KEYINPUT113), .Z(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n513), .A2(new_n510), .ZN(new_n1016));
  INV_X1    g591(.A(new_n507), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1384), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT45), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n477), .A2(G40), .A3(new_n487), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1015), .A2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n1025), .B(KEYINPUT114), .ZN(new_n1026));
  INV_X1    g601(.A(new_n772), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1027), .A2(G1996), .A3(new_n1024), .ZN(new_n1028));
  INV_X1    g603(.A(G1996), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1024), .A2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n1030), .B(KEYINPUT112), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1026), .B(new_n1028), .C1(new_n1027), .C2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n846), .B(new_n849), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1032), .B1(new_n1024), .B2(new_n1033), .ZN(new_n1034));
  OR2_X1    g609(.A1(G290), .A2(G1986), .ZN(new_n1035));
  NAND2_X1  g610(.A1(G290), .A2(G1986), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(KEYINPUT111), .A3(new_n1036), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1037), .B(new_n1024), .C1(KEYINPUT111), .C2(new_n1036), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n1034), .A2(new_n1038), .ZN(new_n1039));
  XOR2_X1   g614(.A(KEYINPUT116), .B(G8), .Z(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(G286), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT115), .B1(G164), .B2(G1384), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1018), .A2(new_n1044), .A3(new_n1019), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT50), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1043), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1023), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1020), .A2(KEYINPUT50), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1050), .A2(G2084), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1044), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1052));
  AOI211_X1 g627(.A(KEYINPUT115), .B(G1384), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1021), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT119), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1054), .A2(new_n1055), .A3(new_n1048), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT45), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1057));
  OAI21_X1  g632(.A(KEYINPUT119), .B1(new_n1057), .B2(new_n1023), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1018), .A2(KEYINPUT45), .A3(new_n1019), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1056), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1051), .B1(new_n1060), .B2(new_n761), .ZN(new_n1061));
  INV_X1    g636(.A(G8), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1042), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NOR3_X1   g638(.A1(G164), .A2(new_n1021), .A3(G1384), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1023), .B1(new_n1065), .B2(new_n1021), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1064), .B1(new_n1066), .B2(new_n1055), .ZN(new_n1067));
  AOI21_X1  g642(.A(G1966), .B1(new_n1067), .B2(new_n1058), .ZN(new_n1068));
  OAI211_X1 g643(.A(G286), .B(new_n1041), .C1(new_n1068), .C2(new_n1051), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1063), .A2(new_n1069), .A3(KEYINPUT51), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT51), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1071), .B(new_n1042), .C1(new_n1061), .C2(new_n1040), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1070), .A2(KEYINPUT62), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1046), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1020), .A2(KEYINPUT50), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1076), .A2(new_n1023), .ZN(new_n1077));
  INV_X1    g652(.A(G2090), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1075), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G1971), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1022), .A2(new_n1059), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1080), .B1(new_n1081), .B2(new_n1023), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1079), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT118), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1079), .A2(new_n1085), .A3(new_n1082), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1084), .A2(new_n1041), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT55), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1088), .B1(G166), .B2(new_n1062), .ZN(new_n1089));
  NAND3_X1  g664(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1087), .A2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1047), .A2(new_n1048), .A3(new_n1078), .A4(new_n1049), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1082), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1091), .A2(new_n1095), .A3(G8), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n824), .A2(G1976), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1097), .B(new_n1041), .C1(new_n1023), .C2(new_n1065), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT52), .ZN(new_n1099));
  INV_X1    g674(.A(G86), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n534), .A2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(G1981), .B1(new_n616), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(G305), .B2(G1981), .ZN(new_n1103));
  NOR2_X1   g678(.A1(KEYINPUT117), .A2(KEYINPUT49), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI221_X1 g680(.A(new_n1102), .B1(KEYINPUT117), .B2(KEYINPUT49), .C1(G305), .C2(G1981), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1065), .A2(new_n1023), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1107), .A2(new_n1040), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1105), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(G1976), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT52), .B1(G288), .B2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1108), .A2(new_n1097), .A3(new_n1111), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1096), .A2(new_n1099), .A3(new_n1109), .A4(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT53), .ZN(new_n1115));
  AOI21_X1  g690(.A(KEYINPUT45), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1064), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n1048), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1115), .B1(new_n1118), .B2(G2078), .ZN(new_n1119));
  INV_X1    g694(.A(G1961), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1050), .A2(new_n1120), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1115), .A2(G2078), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1067), .A2(new_n1058), .A3(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(G301), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n1093), .A2(new_n1114), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1073), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(KEYINPUT62), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT126), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1113), .B1(new_n1092), .B2(new_n1087), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1122), .A2(new_n1124), .A3(G301), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT54), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1081), .A2(new_n1023), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n1123), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1119), .A2(new_n1134), .A3(new_n1121), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1132), .B1(new_n1135), .B2(G171), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1131), .A2(new_n1136), .ZN(new_n1137));
  AND4_X1   g712(.A1(new_n1070), .A2(new_n1130), .A3(new_n1137), .A4(new_n1072), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT57), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n590), .A2(new_n583), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1139), .B1(new_n1140), .B2(KEYINPUT121), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n642), .A2(new_n1141), .ZN(new_n1142));
  OR2_X1    g717(.A1(new_n642), .A2(new_n1141), .ZN(new_n1143));
  AOI21_X1  g718(.A(G1956), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1144));
  XNOR2_X1  g719(.A(KEYINPUT56), .B(G2072), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(KEYINPUT122), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1117), .A2(new_n1048), .A3(new_n1146), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1142), .B(new_n1143), .C1(new_n1144), .C2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1050), .A2(new_n740), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1107), .A2(new_n793), .ZN(new_n1150));
  AND2_X1   g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1148), .B1(new_n1151), .B2(new_n649), .ZN(new_n1152));
  INV_X1    g727(.A(G1956), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1048), .B1(KEYINPUT50), .B2(new_n1020), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1153), .B1(new_n1154), .B2(new_n1074), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1133), .A2(new_n1146), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1143), .A2(new_n1142), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1152), .A2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1151), .A2(KEYINPUT60), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1149), .A2(new_n1150), .A3(KEYINPUT60), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(KEYINPUT124), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(new_n638), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1161), .A2(KEYINPUT124), .A3(new_n649), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  OR2_X1    g740(.A1(new_n1161), .A2(KEYINPUT124), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1160), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1148), .A2(new_n1158), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT61), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1148), .A2(new_n1158), .A3(KEYINPUT61), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT59), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1117), .A2(new_n1029), .A3(new_n1048), .ZN(new_n1173));
  XOR2_X1   g748(.A(KEYINPUT58), .B(G1341), .Z(new_n1174));
  OAI21_X1  g749(.A(new_n1174), .B1(new_n1065), .B2(new_n1023), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n864), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1172), .B1(new_n1176), .B2(KEYINPUT123), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1176), .A2(KEYINPUT123), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NOR3_X1   g754(.A1(new_n1176), .A2(KEYINPUT123), .A3(new_n1172), .ZN(new_n1180));
  OAI211_X1 g755(.A(new_n1170), .B(new_n1171), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1159), .B1(new_n1167), .B2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1135), .A2(G171), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1132), .B1(new_n1125), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1184), .A2(KEYINPUT125), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT125), .ZN(new_n1186));
  OAI211_X1 g761(.A(new_n1186), .B(new_n1132), .C1(new_n1125), .C2(new_n1183), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1138), .A2(new_n1182), .A3(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT63), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1095), .A2(G8), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1190), .B1(new_n1191), .B2(new_n1092), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT120), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n1061), .A2(new_n1040), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1193), .B1(new_n1194), .B2(G168), .ZN(new_n1195));
  NOR4_X1   g770(.A1(new_n1061), .A2(KEYINPUT120), .A3(G286), .A4(new_n1040), .ZN(new_n1196));
  OAI211_X1 g771(.A(new_n1114), .B(new_n1192), .C1(new_n1195), .C2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1093), .A2(new_n1114), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1194), .A2(G168), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1199), .A2(KEYINPUT120), .ZN(new_n1200));
  INV_X1    g775(.A(new_n1196), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1198), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1197), .B1(new_n1202), .B2(KEYINPUT63), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1099), .A2(new_n1109), .A3(new_n1112), .ZN(new_n1204));
  NOR2_X1   g779(.A1(new_n1204), .A2(new_n1096), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1109), .A2(new_n1110), .A3(new_n824), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1206), .B1(G1981), .B2(G305), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1205), .B1(new_n1207), .B2(new_n1108), .ZN(new_n1208));
  NAND4_X1  g783(.A1(new_n1129), .A2(new_n1189), .A3(new_n1203), .A4(new_n1208), .ZN(new_n1209));
  NOR3_X1   g784(.A1(new_n1127), .A2(KEYINPUT126), .A3(new_n1128), .ZN(new_n1210));
  OAI21_X1  g785(.A(new_n1039), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NOR3_X1   g786(.A1(new_n1035), .A2(new_n1023), .A3(new_n1022), .ZN(new_n1212));
  XOR2_X1   g787(.A(new_n1212), .B(KEYINPUT48), .Z(new_n1213));
  NAND2_X1  g788(.A1(new_n1034), .A2(new_n1213), .ZN(new_n1214));
  OAI21_X1  g789(.A(new_n1024), .B1(new_n1015), .B2(new_n1027), .ZN(new_n1215));
  AND2_X1   g790(.A1(new_n1031), .A2(KEYINPUT46), .ZN(new_n1216));
  NOR2_X1   g791(.A1(new_n1031), .A2(KEYINPUT46), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n1215), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  XNOR2_X1  g793(.A(new_n1218), .B(KEYINPUT47), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1214), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n846), .A2(new_n849), .ZN(new_n1221));
  OAI21_X1  g796(.A(new_n1011), .B1(new_n1032), .B2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g797(.A(new_n1220), .B1(new_n1024), .B2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1211), .A2(new_n1223), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g799(.A(new_n906), .ZN(new_n1226));
  NOR3_X1   g800(.A1(G401), .A2(new_n461), .A3(G227), .ZN(new_n1227));
  XOR2_X1   g801(.A(new_n1227), .B(KEYINPUT127), .Z(new_n1228));
  NOR2_X1   g802(.A1(G229), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g803(.A1(new_n1226), .A2(new_n1005), .A3(new_n1229), .ZN(G225));
  INV_X1    g804(.A(G225), .ZN(G308));
endmodule


