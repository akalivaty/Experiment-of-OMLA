//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 1 0 1 0 1 1 0 1 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 0 1 1 0 0 0 0 1 1 1 0 0 1 0 1 1 1 1 0 0 0 1 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998;
  INV_X1    g000(.A(KEYINPUT75), .ZN(new_n187));
  NOR2_X1   g001(.A1(G472), .A2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT32), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G128), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT65), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(new_n196), .A3(G143), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n198), .B1(new_n193), .B2(G143), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n197), .A2(new_n200), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n194), .A2(new_n196), .A3(KEYINPUT66), .A4(G143), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n192), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT0), .ZN(new_n204));
  INV_X1    g018(.A(G137), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G134), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT11), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n205), .A2(KEYINPUT11), .A3(G134), .ZN(new_n209));
  INV_X1    g023(.A(G134), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G137), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n208), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G131), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT67), .B(G131), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n214), .A2(new_n208), .A3(new_n209), .A4(new_n211), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G143), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(G146), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT65), .B(G146), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n219), .B1(new_n220), .B2(G143), .ZN(new_n221));
  OR3_X1    g035(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n222));
  NAND2_X1  g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n204), .A2(new_n216), .A3(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n199), .B1(new_n220), .B2(G143), .ZN(new_n228));
  AND4_X1   g042(.A1(KEYINPUT66), .A2(new_n194), .A3(new_n196), .A4(G143), .ZN(new_n229));
  OAI211_X1 g043(.A(G128), .B(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT70), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n201), .A2(new_n202), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT70), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n232), .A2(new_n233), .A3(G128), .A4(new_n227), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT71), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT1), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT69), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT1), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n192), .B1(new_n197), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n194), .A2(new_n196), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n218), .B1(new_n242), .B2(new_n217), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n235), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n227), .B1(G143), .B2(new_n220), .ZN(new_n245));
  OAI211_X1 g059(.A(KEYINPUT71), .B(new_n221), .C1(new_n245), .C2(new_n192), .ZN(new_n246));
  AOI22_X1  g060(.A1(new_n231), .A2(new_n234), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n206), .A2(new_n211), .A3(new_n248), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n249), .B(G131), .C1(new_n248), .C2(new_n206), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(new_n215), .ZN(new_n251));
  OAI211_X1 g065(.A(KEYINPUT30), .B(new_n226), .C1(new_n247), .C2(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(G116), .B(G119), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT2), .B(G113), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n253), .B(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT72), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n204), .A2(new_n216), .A3(new_n225), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n246), .A2(new_n244), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n230), .A2(KEYINPUT70), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n233), .B1(new_n203), .B2(new_n227), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n251), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n259), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n258), .B1(new_n265), .B2(KEYINPUT30), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n226), .B1(new_n247), .B2(new_n251), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT30), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n267), .A2(KEYINPUT72), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n257), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n226), .B(new_n255), .C1(new_n247), .C2(new_n251), .ZN(new_n271));
  NOR2_X1   g085(.A1(G237), .A2(G953), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G210), .ZN(new_n273));
  XOR2_X1   g087(.A(new_n273), .B(KEYINPUT27), .Z(new_n274));
  XNOR2_X1  g088(.A(KEYINPUT26), .B(G101), .ZN(new_n275));
  XOR2_X1   g089(.A(new_n274), .B(new_n275), .Z(new_n276));
  NAND2_X1  g090(.A1(new_n271), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT73), .B1(new_n270), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n255), .B1(new_n265), .B2(KEYINPUT30), .ZN(new_n279));
  AND3_X1   g093(.A1(new_n267), .A2(KEYINPUT72), .A3(new_n268), .ZN(new_n280));
  AOI21_X1  g094(.A(KEYINPUT72), .B1(new_n267), .B2(new_n268), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT73), .ZN(new_n283));
  INV_X1    g097(.A(new_n277), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n278), .A2(new_n285), .A3(KEYINPUT31), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n263), .A2(new_n264), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n255), .B1(new_n287), .B2(new_n226), .ZN(new_n288));
  INV_X1    g102(.A(new_n271), .ZN(new_n289));
  OAI21_X1  g103(.A(KEYINPUT28), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT28), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n271), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT74), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT74), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n271), .A2(new_n294), .A3(new_n291), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n290), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n276), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT31), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n282), .A2(new_n299), .A3(new_n284), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n191), .B1(new_n286), .B2(new_n301), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n290), .A2(new_n276), .A3(new_n293), .A4(new_n295), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT29), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n276), .B1(new_n282), .B2(new_n271), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n267), .A2(new_n256), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n291), .B1(new_n308), .B2(new_n271), .ZN(new_n309));
  INV_X1    g123(.A(new_n295), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n311), .A2(KEYINPUT29), .A3(new_n276), .A4(new_n293), .ZN(new_n312));
  INV_X1    g126(.A(G902), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(G472), .B1(new_n307), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n302), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n270), .A2(new_n277), .ZN(new_n317));
  AOI22_X1  g131(.A1(new_n317), .A2(new_n299), .B1(new_n296), .B2(new_n297), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n278), .A2(new_n285), .A3(KEYINPUT31), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(KEYINPUT32), .B1(new_n320), .B2(new_n188), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n187), .B1(new_n316), .B2(new_n321), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n312), .B(new_n313), .C1(new_n305), .C2(new_n306), .ZN(new_n323));
  AOI22_X1  g137(.A1(new_n320), .A2(new_n191), .B1(new_n323), .B2(G472), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n188), .B1(new_n286), .B2(new_n301), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n190), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(new_n326), .A3(KEYINPUT75), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT76), .B(G217), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n328), .B1(G234), .B2(new_n313), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n192), .A2(G119), .ZN(new_n330));
  INV_X1    g144(.A(G119), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G128), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT24), .B(G110), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n330), .A2(KEYINPUT77), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT23), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT23), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n330), .A2(KEYINPUT77), .A3(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n337), .A2(new_n332), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n335), .B1(new_n340), .B2(G110), .ZN(new_n341));
  NOR2_X1   g155(.A1(G125), .A2(G140), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT78), .B(G125), .ZN(new_n344));
  INV_X1    g158(.A(G140), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT16), .ZN(new_n347));
  OR2_X1    g161(.A1(KEYINPUT16), .A2(G140), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n347), .A2(G146), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(G146), .B1(new_n347), .B2(new_n350), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n341), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G125), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n355), .A2(new_n345), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n220), .B1(new_n342), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G110), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n337), .A2(new_n339), .A3(new_n358), .A4(new_n332), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT79), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n333), .A2(new_n334), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n360), .B1(new_n359), .B2(new_n361), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n351), .B(new_n357), .C1(new_n362), .C2(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT22), .B(G137), .ZN(new_n365));
  INV_X1    g179(.A(G953), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(G221), .A3(G234), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n365), .B(new_n367), .ZN(new_n368));
  AND3_X1   g182(.A1(new_n354), .A2(new_n364), .A3(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n368), .B1(new_n354), .B2(new_n364), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(KEYINPUT25), .B1(new_n371), .B2(new_n313), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT25), .ZN(new_n373));
  NOR4_X1   g187(.A1(new_n369), .A2(new_n370), .A3(new_n373), .A4(G902), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n329), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n329), .A2(G902), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n371), .A2(new_n377), .ZN(new_n378));
  OR2_X1    g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n322), .A2(new_n327), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT80), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n322), .A2(new_n327), .A3(KEYINPUT80), .A4(new_n380), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(G214), .B1(G237), .B2(G902), .ZN(new_n386));
  XOR2_X1   g200(.A(new_n386), .B(KEYINPUT87), .Z(new_n387));
  XOR2_X1   g201(.A(new_n387), .B(KEYINPUT88), .Z(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G224), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n390), .A2(G953), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT7), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n344), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n204), .A2(new_n225), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n396), .B1(new_n263), .B2(new_n344), .ZN(new_n397));
  NAND2_X1  g211(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n394), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n247), .A2(new_n395), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n393), .B(new_n398), .C1(new_n401), .C2(new_n396), .ZN(new_n402));
  INV_X1    g216(.A(new_n253), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(new_n254), .ZN(new_n404));
  XOR2_X1   g218(.A(KEYINPUT89), .B(KEYINPUT5), .Z(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(G116), .A3(new_n331), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n406), .B(KEYINPUT90), .ZN(new_n407));
  INV_X1    g221(.A(G113), .ZN(new_n408));
  INV_X1    g222(.A(new_n405), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n408), .B1(new_n409), .B2(new_n253), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n404), .B1(new_n407), .B2(new_n410), .ZN(new_n411));
  OR2_X1    g225(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n412));
  INV_X1    g226(.A(G107), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G104), .ZN(new_n414));
  AND2_X1   g228(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n412), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G101), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n413), .A2(G104), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G104), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n420), .A2(G107), .ZN(new_n421));
  NOR2_X1   g235(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n416), .A2(new_n417), .A3(new_n419), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT82), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n418), .B1(new_n422), .B2(new_n421), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT82), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n426), .A2(new_n427), .A3(new_n417), .A4(new_n416), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n418), .B(KEYINPUT84), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n414), .B(KEYINPUT83), .ZN(new_n431));
  OAI21_X1  g245(.A(G101), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n411), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(G110), .B(G122), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(KEYINPUT8), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n408), .B1(new_n253), .B2(KEYINPUT5), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n404), .B1(new_n407), .B2(new_n437), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n434), .B(new_n436), .C1(new_n433), .C2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n400), .A2(new_n402), .A3(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT94), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT85), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n433), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n429), .A2(KEYINPUT85), .A3(new_n432), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(new_n411), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n426), .A2(new_n416), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(G101), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT4), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n425), .A2(new_n428), .B1(G101), .B2(new_n447), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n450), .B1(new_n451), .B2(new_n449), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n256), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n446), .A2(new_n453), .A3(new_n435), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n400), .A2(new_n402), .A3(KEYINPUT94), .A4(new_n439), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n442), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT6), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n446), .A2(new_n453), .ZN(new_n458));
  XOR2_X1   g272(.A(new_n435), .B(KEYINPUT91), .Z(new_n459));
  AOI21_X1  g273(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n454), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n397), .B(new_n391), .ZN(new_n462));
  INV_X1    g276(.A(new_n459), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n463), .B1(new_n446), .B2(new_n453), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT92), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n464), .A2(new_n465), .A3(new_n457), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n465), .B1(new_n464), .B2(new_n457), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n461), .B(new_n462), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n456), .A2(new_n468), .A3(new_n313), .ZN(new_n469));
  OAI21_X1  g283(.A(G210), .B1(G237), .B2(G902), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n456), .A2(new_n468), .A3(new_n313), .A4(new_n470), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n389), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(G234), .A2(G237), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n475), .A2(G952), .A3(new_n366), .ZN(new_n476));
  XOR2_X1   g290(.A(KEYINPUT21), .B(G898), .Z(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(KEYINPUT100), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n475), .A2(G902), .A3(G953), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n480), .B(KEYINPUT99), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n476), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n474), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n353), .ZN(new_n486));
  INV_X1    g300(.A(new_n214), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n272), .A2(G143), .A3(G214), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(G143), .B1(new_n272), .B2(G214), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n487), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT17), .ZN(new_n492));
  OR2_X1    g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n490), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(new_n214), .A3(new_n488), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n491), .A2(new_n495), .A3(new_n492), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n486), .A2(new_n351), .A3(new_n493), .A4(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(G113), .B(G122), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n498), .B(new_n420), .ZN(new_n499));
  NAND2_X1  g313(.A1(KEYINPUT18), .A2(G131), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n494), .A2(new_n488), .A3(new_n500), .ZN(new_n501));
  OAI211_X1 g315(.A(KEYINPUT18), .B(G131), .C1(new_n489), .C2(new_n490), .ZN(new_n502));
  OAI211_X1 g316(.A(G146), .B(new_n343), .C1(new_n344), .C2(new_n345), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT95), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n357), .B1(new_n503), .B2(new_n504), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n501), .B(new_n502), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n497), .A2(new_n499), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n491), .A2(new_n495), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT19), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n510), .B1(new_n356), .B2(new_n342), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n220), .B(new_n511), .C1(new_n346), .C2(new_n510), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n351), .A2(new_n509), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n507), .A2(KEYINPUT96), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n499), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(KEYINPUT96), .B1(new_n507), .B2(new_n513), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n508), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT97), .ZN(new_n519));
  NOR2_X1   g333(.A1(G475), .A2(G902), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n520), .B(KEYINPUT98), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT97), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n523), .B(new_n508), .C1(new_n516), .C2(new_n517), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n519), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n521), .A2(KEYINPUT20), .ZN(new_n526));
  AOI22_X1  g340(.A1(new_n525), .A2(KEYINPUT20), .B1(new_n518), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n497), .A2(new_n507), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n515), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n508), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n313), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(G475), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n527), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n192), .A2(G143), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n217), .A2(G128), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(new_n210), .ZN(new_n538));
  INV_X1    g352(.A(G116), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n539), .A2(KEYINPUT14), .A3(G122), .ZN(new_n540));
  XNOR2_X1  g354(.A(G116), .B(G122), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  OAI211_X1 g356(.A(G107), .B(new_n540), .C1(new_n542), .C2(KEYINPUT14), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n538), .B(new_n543), .C1(G107), .C2(new_n542), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n535), .A2(KEYINPUT13), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(new_n536), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n535), .A2(KEYINPUT13), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n210), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n541), .B(new_n413), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n537), .A2(new_n210), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n544), .B1(new_n548), .B2(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT9), .B(G234), .ZN(new_n553));
  NOR3_X1   g367(.A1(new_n328), .A2(new_n553), .A3(G953), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n552), .A2(new_n555), .ZN(new_n557));
  OR2_X1    g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n313), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT15), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n560), .A3(G478), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(G478), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n558), .A2(new_n313), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n534), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(G469), .ZN(new_n566));
  XNOR2_X1  g380(.A(G110), .B(G140), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n366), .A2(G227), .ZN(new_n568));
  XOR2_X1   g382(.A(new_n567), .B(new_n568), .Z(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n231), .A2(new_n234), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n571), .A2(new_n260), .A3(new_n433), .ZN(new_n572));
  INV_X1    g386(.A(new_n232), .ZN(new_n573));
  OAI21_X1  g387(.A(G128), .B1(new_n218), .B2(new_n236), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n433), .B1(new_n571), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n216), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT12), .ZN(new_n578));
  OR2_X1    g392(.A1(new_n578), .A2(KEYINPUT86), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(KEYINPUT86), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n577), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n247), .A2(new_n433), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n231), .A2(new_n234), .B1(new_n573), .B2(new_n574), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n582), .B1(new_n433), .B2(new_n583), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n584), .A2(KEYINPUT86), .A3(new_n578), .A4(new_n216), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n263), .A2(new_n444), .A3(KEYINPUT10), .A4(new_n445), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n452), .A2(new_n204), .A3(new_n225), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT10), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n588), .B1(new_n583), .B2(new_n433), .ZN(new_n589));
  INV_X1    g403(.A(new_n216), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n586), .A2(new_n587), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  AND4_X1   g405(.A1(new_n570), .A2(new_n581), .A3(new_n585), .A4(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n586), .A2(new_n589), .A3(new_n587), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n216), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n570), .B1(new_n594), .B2(new_n591), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n566), .B(new_n313), .C1(new_n592), .C2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n581), .A2(new_n585), .A3(new_n591), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n569), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n591), .A2(new_n570), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n594), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n598), .A2(new_n600), .A3(G469), .ZN(new_n601));
  NAND2_X1  g415(.A1(G469), .A2(G902), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n596), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(G221), .B1(new_n553), .B2(G902), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n565), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  AND2_X1   g419(.A1(new_n485), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n385), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G101), .ZN(G3));
  NAND3_X1  g422(.A1(new_n458), .A2(new_n457), .A3(new_n459), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(KEYINPUT92), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n464), .A2(new_n465), .A3(new_n457), .ZN(new_n611));
  AOI22_X1  g425(.A1(new_n610), .A2(new_n611), .B1(new_n454), .B2(new_n460), .ZN(new_n612));
  AOI21_X1  g426(.A(G902), .B1(new_n612), .B2(new_n462), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n470), .B1(new_n613), .B2(new_n456), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n473), .B1(new_n614), .B2(KEYINPUT101), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n469), .A2(KEYINPUT101), .A3(new_n471), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n387), .ZN(new_n619));
  NAND2_X1  g433(.A1(G478), .A2(G902), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n620), .B1(new_n559), .B2(G478), .ZN(new_n621));
  XOR2_X1   g435(.A(new_n558), .B(KEYINPUT33), .Z(new_n622));
  AOI21_X1  g436(.A(new_n621), .B1(new_n622), .B2(G478), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n534), .A2(new_n484), .A3(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n618), .A2(new_n619), .A3(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(G472), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n627), .B1(new_n320), .B2(new_n313), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n189), .B1(new_n318), .B2(new_n319), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n603), .A2(new_n604), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n630), .A2(new_n380), .A3(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n626), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT102), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT34), .B(G104), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  AOI21_X1  g450(.A(new_n387), .B1(new_n615), .B2(new_n617), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n519), .A2(new_n524), .A3(new_n526), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT103), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n640), .A2(new_n533), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n525), .A2(KEYINPUT20), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n642), .A2(new_n639), .A3(new_n638), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n637), .A2(new_n484), .A3(new_n564), .A4(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n645), .A2(new_n632), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT105), .B(G107), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT104), .B(KEYINPUT35), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  NAND2_X1  g464(.A1(new_n354), .A2(new_n364), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT106), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n368), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(KEYINPUT36), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n651), .B(KEYINPUT106), .ZN(new_n657));
  INV_X1    g471(.A(new_n655), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n656), .A2(new_n659), .A3(new_n377), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n376), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n485), .A2(new_n605), .A3(new_n630), .A4(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT37), .B(G110), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G12));
  NAND4_X1  g479(.A1(new_n322), .A2(new_n327), .A3(new_n631), .A4(new_n662), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n481), .A2(G900), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(KEYINPUT107), .ZN(new_n668));
  INV_X1    g482(.A(new_n476), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n667), .A2(KEYINPUT107), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  AND4_X1   g487(.A1(new_n564), .A2(new_n641), .A3(new_n643), .A4(new_n673), .ZN(new_n674));
  AND4_X1   g488(.A1(new_n313), .A2(new_n456), .A3(new_n468), .A4(new_n470), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT101), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n675), .B1(new_n676), .B2(new_n472), .ZN(new_n677));
  OAI211_X1 g491(.A(new_n619), .B(new_n674), .C1(new_n677), .C2(new_n616), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(KEYINPUT108), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT108), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n618), .A2(new_n680), .A3(new_n619), .A4(new_n674), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n666), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(new_n192), .ZN(G30));
  XOR2_X1   g497(.A(new_n672), .B(KEYINPUT39), .Z(new_n684));
  NAND2_X1  g498(.A1(new_n631), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(new_n685), .B(KEYINPUT40), .Z(new_n686));
  NAND2_X1  g500(.A1(new_n472), .A2(new_n473), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT109), .B(KEYINPUT38), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n297), .B1(new_n288), .B2(new_n289), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n278), .A2(new_n285), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n313), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(G472), .ZN(new_n693));
  OAI211_X1 g507(.A(new_n302), .B(new_n693), .C1(new_n629), .C2(KEYINPUT32), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n527), .A2(new_n533), .ZN(new_n695));
  INV_X1    g509(.A(new_n564), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AND4_X1   g511(.A1(new_n619), .A2(new_n694), .A3(new_n661), .A4(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n686), .A2(new_n689), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G143), .ZN(G45));
  NAND3_X1  g514(.A1(new_n534), .A2(new_n623), .A3(new_n673), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n702), .B(new_n619), .C1(new_n677), .C2(new_n616), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n666), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n193), .ZN(G48));
  NAND3_X1  g519(.A1(new_n599), .A2(new_n585), .A3(new_n581), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n594), .A2(new_n591), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n569), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n313), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(G469), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n596), .ZN(new_n712));
  INV_X1    g526(.A(new_n604), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n712), .A2(new_n379), .A3(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n322), .A2(new_n327), .A3(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n715), .A2(new_n626), .ZN(new_n716));
  XOR2_X1   g530(.A(KEYINPUT41), .B(G113), .Z(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G15));
  NOR2_X1   g532(.A1(new_n645), .A2(new_n715), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(new_n539), .ZN(G18));
  AND2_X1   g534(.A1(new_n322), .A2(new_n327), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n619), .B1(new_n677), .B2(new_n616), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n566), .B1(new_n709), .B2(new_n313), .ZN(new_n723));
  INV_X1    g537(.A(new_n596), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n725), .A2(new_n565), .A3(new_n484), .A4(new_n604), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT110), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n721), .A2(new_n727), .A3(new_n728), .A4(new_n662), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n322), .A2(new_n327), .A3(new_n662), .ZN(new_n730));
  NOR4_X1   g544(.A1(new_n723), .A2(new_n724), .A3(new_n483), .A4(new_n713), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n618), .A2(new_n619), .A3(new_n565), .A4(new_n731), .ZN(new_n732));
  OAI21_X1  g546(.A(KEYINPUT110), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g548(.A(KEYINPUT111), .B(G119), .Z(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G21));
  NAND4_X1  g550(.A1(new_n618), .A2(new_n731), .A3(new_n619), .A4(new_n697), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n319), .A2(new_n298), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT112), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT112), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n319), .A2(new_n740), .A3(new_n298), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n739), .A2(new_n300), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n628), .B1(new_n742), .B2(new_n188), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n380), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n737), .A2(new_n744), .ZN(new_n745));
  XOR2_X1   g559(.A(new_n745), .B(G122), .Z(G24));
  NAND2_X1  g560(.A1(new_n741), .A2(new_n300), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n740), .B1(new_n319), .B2(new_n298), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n188), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n628), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(new_n750), .A3(new_n662), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n712), .A2(new_n713), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n751), .A2(new_n703), .A3(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(new_n355), .ZN(G27));
  INV_X1    g569(.A(KEYINPUT42), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n472), .A2(new_n473), .A3(new_n619), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n602), .B(KEYINPUT113), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n596), .A2(new_n601), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n604), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n322), .A2(new_n327), .A3(new_n380), .A4(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n756), .B1(new_n762), .B2(new_n701), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n757), .A2(new_n760), .A3(new_n701), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n379), .B1(new_n324), .B2(new_n326), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(new_n765), .A3(KEYINPUT42), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G131), .ZN(G33));
  INV_X1    g582(.A(new_n674), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n762), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G134), .ZN(G36));
  XNOR2_X1  g585(.A(new_n757), .B(KEYINPUT114), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n623), .A2(new_n695), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(KEYINPUT43), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n774), .A2(new_n661), .ZN(new_n775));
  OAI21_X1  g589(.A(KEYINPUT44), .B1(new_n775), .B2(new_n630), .ZN(new_n776));
  OR4_X1    g590(.A1(KEYINPUT44), .A2(new_n774), .A3(new_n630), .A4(new_n661), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n772), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n598), .A2(new_n600), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT45), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(G469), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n779), .A2(new_n780), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n758), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT46), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n724), .B1(new_n784), .B2(new_n785), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n713), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n684), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n778), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G137), .ZN(G39));
  NOR4_X1   g606(.A1(new_n721), .A2(new_n380), .A3(new_n701), .A4(new_n757), .ZN(new_n793));
  XOR2_X1   g607(.A(KEYINPUT115), .B(KEYINPUT47), .Z(new_n794));
  NAND2_X1  g608(.A1(new_n788), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n796), .A2(KEYINPUT47), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n793), .B(new_n795), .C1(new_n788), .C2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G140), .ZN(G42));
  NOR4_X1   g613(.A1(new_n773), .A2(new_n379), .A3(new_n389), .A4(new_n713), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT49), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n800), .B1(new_n801), .B2(new_n725), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n712), .A2(KEYINPUT49), .ZN(new_n803));
  OR4_X1    g617(.A1(new_n689), .A2(new_n802), .A3(new_n694), .A4(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n757), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n752), .A2(new_n805), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n806), .A2(new_n669), .A3(new_n774), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n765), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT48), .ZN(new_n809));
  INV_X1    g623(.A(G952), .ZN(new_n810));
  NOR4_X1   g624(.A1(new_n806), .A2(new_n379), .A3(new_n669), .A4(new_n694), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n534), .A2(new_n623), .ZN(new_n812));
  AOI211_X1 g626(.A(new_n810), .B(G953), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n774), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n814), .A2(new_n743), .A3(new_n380), .A4(new_n476), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n637), .A2(new_n752), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n809), .B(new_n813), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  OR3_X1    g631(.A1(new_n689), .A2(new_n753), .A3(new_n619), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n818), .A2(new_n815), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n819), .B1(KEYINPUT118), .B2(KEYINPUT50), .ZN(new_n820));
  XOR2_X1   g634(.A(KEYINPUT118), .B(KEYINPUT50), .Z(new_n821));
  OAI21_X1  g635(.A(new_n820), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n534), .A2(new_n623), .ZN(new_n823));
  INV_X1    g637(.A(new_n751), .ZN(new_n824));
  AOI22_X1  g638(.A1(new_n811), .A2(new_n823), .B1(new_n807), .B2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n795), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n788), .A2(new_n797), .ZN(new_n827));
  OAI22_X1  g641(.A1(new_n826), .A2(new_n827), .B1(new_n604), .B2(new_n712), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n815), .A2(new_n772), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n822), .B(new_n825), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT51), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n817), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n830), .B1(new_n828), .B2(KEYINPUT120), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n834), .B1(KEYINPUT120), .B2(new_n828), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT119), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n825), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n832), .B1(new_n825), .B2(new_n836), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n835), .A2(new_n822), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n833), .A2(new_n839), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n376), .A2(new_n660), .A3(new_n672), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n759), .A2(new_n604), .A3(new_n841), .ZN(new_n842));
  AOI22_X1  g656(.A1(new_n320), .A2(new_n191), .B1(new_n692), .B2(G472), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n842), .B1(new_n326), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n637), .A2(new_n844), .A3(new_n697), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n845), .B1(new_n666), .B2(new_n703), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n847));
  NOR4_X1   g661(.A1(new_n682), .A2(new_n846), .A3(new_n847), .A4(new_n754), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n679), .A2(new_n681), .ZN(new_n849));
  AND4_X1   g663(.A1(new_n322), .A2(new_n327), .A3(new_n631), .A4(new_n662), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n703), .A2(new_n753), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n849), .A2(new_n850), .B1(new_n851), .B2(new_n824), .ZN(new_n852));
  INV_X1    g666(.A(new_n760), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n694), .A2(new_n853), .A3(new_n841), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n619), .B(new_n697), .C1(new_n677), .C2(new_n616), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n703), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n856), .B1(new_n850), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT52), .B1(new_n852), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n848), .A2(new_n859), .ZN(new_n860));
  AOI22_X1  g674(.A1(new_n385), .A2(new_n606), .B1(new_n729), .B2(new_n733), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n743), .A2(new_n764), .A3(new_n662), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n561), .A2(new_n563), .A3(new_n673), .ZN(new_n863));
  INV_X1    g677(.A(new_n660), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n863), .B1(new_n864), .B2(new_n375), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n644), .A2(new_n603), .A3(new_n604), .A4(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n866), .A2(new_n757), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n867), .A2(new_n322), .A3(new_n327), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n862), .B(new_n868), .C1(new_n762), .C2(new_n769), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n869), .B1(new_n763), .B2(new_n766), .ZN(new_n870));
  OAI22_X1  g684(.A1(new_n645), .A2(new_n715), .B1(new_n737), .B2(new_n744), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT116), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n534), .A2(new_n696), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n474), .A2(new_n872), .A3(new_n484), .A4(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n625), .A2(new_n474), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n474), .A2(new_n484), .A3(new_n873), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT116), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n632), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n663), .B1(new_n715), .B2(new_n626), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n871), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n861), .A2(new_n870), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT53), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n860), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n861), .A2(new_n870), .A3(new_n881), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n849), .A2(new_n850), .ZN(new_n886));
  INV_X1    g700(.A(new_n754), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n858), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n847), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n852), .A2(KEYINPUT52), .A3(new_n858), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(KEYINPUT53), .B1(new_n885), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(KEYINPUT54), .B1(new_n884), .B2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT117), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n883), .B1(new_n860), .B2(new_n882), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n885), .A2(new_n891), .A3(KEYINPUT53), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT54), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n893), .A2(new_n894), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n897), .B1(new_n895), .B2(new_n896), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(KEYINPUT117), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n840), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(G952), .A2(G953), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT121), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n804), .B1(new_n902), .B2(new_n904), .ZN(G75));
  NAND2_X1  g719(.A1(new_n895), .A2(new_n896), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(G210), .A3(G902), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n612), .B(new_n462), .Z(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT55), .ZN(new_n909));
  XNOR2_X1  g723(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n907), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT56), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n909), .B1(new_n907), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n366), .A2(G952), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n911), .A2(new_n913), .A3(new_n914), .ZN(G51));
  XNOR2_X1  g729(.A(new_n758), .B(KEYINPUT123), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT57), .Z(new_n917));
  AND3_X1   g731(.A1(new_n895), .A2(new_n897), .A3(new_n896), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n917), .B1(new_n918), .B2(new_n900), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n709), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n782), .A2(new_n783), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT124), .Z(new_n922));
  NAND3_X1  g736(.A1(new_n906), .A2(G902), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n914), .B1(new_n920), .B2(new_n923), .ZN(G54));
  NAND4_X1  g738(.A1(new_n906), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n519), .A2(new_n524), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n925), .A2(new_n926), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n927), .A2(new_n928), .A3(new_n914), .ZN(G60));
  XOR2_X1   g743(.A(new_n620), .B(KEYINPUT59), .Z(new_n930));
  NOR2_X1   g744(.A1(new_n622), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(new_n918), .B2(new_n900), .ZN(new_n932));
  INV_X1    g746(.A(new_n914), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n930), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n899), .A2(new_n901), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n934), .B1(new_n622), .B2(new_n936), .ZN(G63));
  AND2_X1   g751(.A1(new_n656), .A2(new_n659), .ZN(new_n938));
  NAND2_X1  g752(.A1(G217), .A2(G902), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT60), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n906), .A2(new_n938), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n940), .B1(new_n895), .B2(new_n896), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n942), .B(new_n933), .C1(new_n371), .C2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(KEYINPUT61), .B1(new_n942), .B2(KEYINPUT125), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OR2_X1    g760(.A1(new_n943), .A2(new_n371), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n914), .B1(new_n943), .B2(new_n938), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT125), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n949), .B1(new_n943), .B2(new_n938), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n947), .B(new_n948), .C1(new_n950), .C2(KEYINPUT61), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n946), .A2(new_n951), .ZN(G66));
  OAI21_X1  g766(.A(G953), .B1(new_n479), .B2(new_n390), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n861), .A2(new_n881), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n953), .B1(new_n955), .B2(G953), .ZN(new_n956));
  INV_X1    g770(.A(new_n612), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(G898), .B2(new_n366), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n956), .B(new_n958), .ZN(G69));
  NOR3_X1   g773(.A1(new_n682), .A2(new_n704), .A3(new_n754), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n699), .ZN(new_n961));
  OR2_X1    g775(.A1(new_n961), .A2(KEYINPUT62), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n805), .B1(new_n812), .B2(new_n873), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n963), .A2(new_n685), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n385), .A2(new_n964), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT126), .Z(new_n966));
  NAND2_X1  g780(.A1(new_n961), .A2(KEYINPUT62), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n791), .A2(new_n798), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n962), .A2(new_n966), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n366), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n252), .B1(new_n280), .B2(new_n281), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n511), .B1(new_n346), .B2(new_n510), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n637), .A2(new_n765), .A3(new_n697), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n770), .B1(new_n789), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(new_n763), .B2(new_n766), .ZN(new_n977));
  AND4_X1   g791(.A1(new_n791), .A2(new_n977), .A3(new_n798), .A4(new_n960), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n366), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n974), .B1(G900), .B2(G953), .ZN(new_n980));
  AOI22_X1  g794(.A1(new_n970), .A2(new_n974), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n366), .B1(G227), .B2(G900), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n968), .A2(new_n960), .A3(new_n977), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n980), .B1(new_n983), .B2(G953), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n982), .B1(new_n984), .B2(KEYINPUT127), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n981), .B(new_n985), .ZN(G72));
  OAI21_X1  g800(.A(new_n276), .B1(new_n270), .B2(new_n289), .ZN(new_n987));
  OR2_X1    g801(.A1(new_n969), .A2(new_n954), .ZN(new_n988));
  NAND2_X1  g802(.A1(G472), .A2(G902), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT63), .Z(new_n990));
  AOI21_X1  g804(.A(new_n987), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n990), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n992), .B1(new_n978), .B2(new_n955), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n270), .A2(new_n289), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n297), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n933), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n278), .B(new_n285), .C1(new_n994), .C2(new_n276), .ZN(new_n997));
  AND3_X1   g811(.A1(new_n906), .A2(new_n990), .A3(new_n997), .ZN(new_n998));
  NOR3_X1   g812(.A1(new_n991), .A2(new_n996), .A3(new_n998), .ZN(G57));
endmodule


