//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 1 1 0 1 1 0 1 0 1 0 1 0 1 0 1 0 1 1 1 0 1 1 0 1 1 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n552,
    new_n554, new_n555, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n615, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1229, new_n1230, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G120), .Z(G236));
  XNOR2_X1  g015(.A(KEYINPUT66), .B(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT67), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT68), .ZN(new_n453));
  NAND4_X1  g028(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G567), .B1(G2106), .B2(new_n455), .ZN(G319));
  NAND2_X1  g033(.A1(G101), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G137), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n461), .A2(new_n463), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n467), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n468), .A2(new_n472), .ZN(G160));
  OAI21_X1  g048(.A(G2104), .B1(new_n467), .B2(G112), .ZN(new_n474));
  INV_X1    g049(.A(G100), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n474), .B1(new_n475), .B2(new_n467), .ZN(new_n476));
  XOR2_X1   g051(.A(new_n476), .B(KEYINPUT69), .Z(new_n477));
  NOR2_X1   g052(.A1(new_n464), .A2(new_n467), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n464), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  NAND2_X1  g058(.A1(KEYINPUT71), .A2(KEYINPUT4), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n469), .A2(new_n467), .ZN(new_n485));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G126), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(new_n467), .ZN(new_n489));
  NOR3_X1   g064(.A1(new_n484), .A2(new_n486), .A3(G2105), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n469), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n493), .B(KEYINPUT70), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n494), .A2(G2104), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n487), .A2(new_n491), .A3(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  XNOR2_X1  g073(.A(KEYINPUT5), .B(G543), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n499), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n500));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g077(.A(KEYINPUT6), .B(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G50), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  OAI211_X1 g086(.A(new_n507), .B(new_n509), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT72), .B(G88), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n504), .A2(new_n505), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n502), .A2(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  NAND3_X1  g091(.A1(new_n499), .A2(G63), .A3(G651), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n503), .A2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G51), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n499), .A2(new_n503), .A3(G89), .ZN(new_n520));
  AND3_X1   g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  OR2_X1    g096(.A1(KEYINPUT73), .A2(KEYINPUT7), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT73), .A2(KEYINPUT7), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  AND2_X1   g100(.A1(KEYINPUT73), .A2(KEYINPUT7), .ZN(new_n526));
  NOR2_X1   g101(.A1(KEYINPUT73), .A2(KEYINPUT7), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n520), .A2(KEYINPUT74), .A3(new_n524), .A4(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n524), .A2(new_n528), .ZN(new_n531));
  AOI21_X1  g106(.A(KEYINPUT74), .B1(new_n531), .B2(new_n520), .ZN(new_n532));
  OAI211_X1 g107(.A(new_n517), .B(new_n519), .C1(new_n530), .C2(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n507), .A2(new_n509), .ZN(new_n536));
  INV_X1    g111(.A(G64), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(KEYINPUT75), .B(G52), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n518), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n499), .A2(new_n503), .A3(G90), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n539), .A2(new_n541), .A3(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  AOI22_X1  g119(.A1(new_n499), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n501), .ZN(new_n546));
  INV_X1    g121(.A(G43), .ZN(new_n547));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n504), .A2(new_n547), .B1(new_n512), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  AND3_X1   g126(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G36), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n552), .A2(new_n555), .ZN(G188));
  NAND2_X1  g131(.A1(new_n512), .A2(KEYINPUT77), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n499), .A2(new_n503), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G91), .ZN(new_n561));
  OAI211_X1 g136(.A(G53), .B(G543), .C1(new_n510), .C2(new_n511), .ZN(new_n562));
  NAND2_X1  g137(.A1(KEYINPUT76), .A2(KEYINPUT9), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n562), .B(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(G78), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n566), .A2(new_n506), .ZN(new_n567));
  AND3_X1   g142(.A1(new_n507), .A2(new_n509), .A3(KEYINPUT78), .ZN(new_n568));
  AOI21_X1  g143(.A(KEYINPUT78), .B1(new_n507), .B2(new_n509), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n567), .B1(new_n570), .B2(G65), .ZN(new_n571));
  OAI211_X1 g146(.A(new_n561), .B(new_n565), .C1(new_n571), .C2(new_n501), .ZN(G299));
  NAND2_X1  g147(.A1(new_n560), .A2(G87), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n499), .B2(G74), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n518), .A2(G49), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(G288));
  NAND2_X1  g151(.A1(new_n560), .A2(G86), .ZN(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT79), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n578), .B(new_n579), .ZN(new_n580));
  AND3_X1   g155(.A1(new_n507), .A2(new_n509), .A3(G61), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT80), .ZN(new_n583));
  INV_X1    g158(.A(G48), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n504), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n518), .A2(KEYINPUT80), .A3(G48), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n577), .A2(new_n582), .A3(new_n585), .A4(new_n586), .ZN(G305));
  AOI22_X1  g162(.A1(new_n499), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(new_n501), .ZN(new_n589));
  INV_X1    g164(.A(G47), .ZN(new_n590));
  INV_X1    g165(.A(G85), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n504), .A2(new_n590), .B1(new_n512), .B2(new_n591), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n589), .A2(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(G301), .A2(G868), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n512), .A2(KEYINPUT77), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n558), .B1(new_n499), .B2(new_n503), .ZN(new_n596));
  OAI21_X1  g171(.A(G92), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(KEYINPUT10), .ZN(new_n598));
  INV_X1    g173(.A(G66), .ZN(new_n599));
  NOR3_X1   g174(.A1(new_n568), .A2(new_n569), .A3(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G79), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(new_n506), .ZN(new_n602));
  OAI21_X1  g177(.A(G651), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n518), .A2(G54), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT10), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n560), .A2(new_n605), .A3(G92), .ZN(new_n606));
  NAND4_X1  g181(.A1(new_n598), .A2(new_n603), .A3(new_n604), .A4(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n594), .B1(new_n608), .B2(G868), .ZN(G284));
  XOR2_X1   g184(.A(G284), .B(KEYINPUT81), .Z(G321));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(G299), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G168), .B2(new_n611), .ZN(G297));
  OAI21_X1  g188(.A(new_n612), .B1(G168), .B2(new_n611), .ZN(G280));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n608), .B1(new_n615), .B2(G860), .ZN(G148));
  NAND2_X1  g191(.A1(new_n608), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G868), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g195(.A1(new_n480), .A2(G2104), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT12), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  INV_X1    g198(.A(G2100), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(KEYINPUT82), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n623), .B(new_n625), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n624), .A2(KEYINPUT82), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n478), .A2(G123), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n480), .A2(G135), .ZN(new_n629));
  OR2_X1    g204(.A1(G99), .A2(G2105), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n630), .B(G2104), .C1(G111), .C2(new_n467), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n628), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT83), .Z(new_n633));
  AOI21_X1  g208(.A(new_n627), .B1(new_n633), .B2(G2096), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n626), .B(new_n634), .C1(G2096), .C2(new_n633), .ZN(G156));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2435), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT84), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G2427), .B(G2430), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(KEYINPUT14), .ZN(new_n641));
  XOR2_X1   g216(.A(G2451), .B(G2454), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT85), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n641), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(G14), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(G401));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  XNOR2_X1  g227(.A(G2067), .B(G2678), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2072), .B(G2078), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT18), .Z(new_n656));
  XOR2_X1   g231(.A(new_n653), .B(KEYINPUT86), .Z(new_n657));
  OAI21_X1  g232(.A(KEYINPUT17), .B1(new_n657), .B2(new_n652), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(new_n654), .Z(new_n659));
  AND2_X1   g234(.A1(new_n657), .A2(new_n652), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n656), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(G2096), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(new_n624), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(G227));
  XOR2_X1   g239(.A(G1956), .B(G2474), .Z(new_n665));
  XOR2_X1   g240(.A(G1961), .B(G1966), .Z(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1971), .B(G1976), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n665), .A2(new_n666), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n668), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT87), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT20), .ZN(new_n675));
  AND2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  OAI221_X1 g252(.A(new_n672), .B1(new_n670), .B2(new_n668), .C1(new_n676), .C2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n680), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT22), .B(G1981), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(G229));
  NOR2_X1   g261(.A1(KEYINPUT24), .A2(G34), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(KEYINPUT24), .A2(G34), .ZN(new_n689));
  AOI21_X1  g264(.A(G29), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  AOI22_X1  g265(.A1(G160), .A2(G29), .B1(KEYINPUT99), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(KEYINPUT99), .B2(new_n690), .ZN(new_n692));
  INV_X1    g267(.A(G2084), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT30), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n695), .A2(G28), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(G28), .ZN(new_n697));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(new_n633), .B2(new_n698), .ZN(new_n700));
  NOR2_X1   g275(.A1(G27), .A2(G29), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(G164), .B2(G29), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n702), .A2(G2078), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT31), .B(G11), .Z(new_n704));
  NOR3_X1   g279(.A1(new_n700), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n478), .A2(G129), .ZN(new_n706));
  NAND3_X1  g281(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT26), .Z(new_n708));
  AOI22_X1  g283(.A1(new_n469), .A2(G141), .B1(G105), .B2(G2104), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n706), .B(new_n708), .C1(new_n709), .C2(G2105), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT100), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G29), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT27), .B(G1996), .Z(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G32), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n713), .B(new_n715), .C1(G29), .C2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G2072), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT97), .ZN(new_n719));
  INV_X1    g294(.A(G139), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n485), .B2(new_n720), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n480), .A2(KEYINPUT97), .A3(G139), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(G115), .A2(G2104), .ZN(new_n724));
  INV_X1    g299(.A(G127), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n724), .B1(new_n464), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G2105), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT25), .Z(new_n729));
  NAND3_X1  g304(.A1(new_n723), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT98), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g307(.A1(new_n723), .A2(KEYINPUT98), .A3(new_n727), .A4(new_n729), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G29), .ZN(new_n735));
  NOR2_X1   g310(.A1(G29), .A2(G33), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n718), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  AOI211_X1 g313(.A(G2072), .B(new_n736), .C1(new_n734), .C2(G29), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n705), .B(new_n717), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G16), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G21), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G168), .B2(new_n741), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G1966), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT92), .B(G1348), .Z(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n741), .A2(G4), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n608), .B2(new_n741), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(KEYINPUT93), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n749), .A2(KEYINPUT93), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n747), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(new_n752), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n754), .A2(new_n746), .A3(new_n750), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n692), .A2(new_n693), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n741), .A2(G19), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n550), .B2(new_n741), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(G1341), .Z(new_n760));
  NAND4_X1  g335(.A1(new_n745), .A2(new_n756), .A3(new_n757), .A4(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(KEYINPUT23), .B1(new_n741), .B2(G20), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G299), .B2(G16), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n741), .A2(KEYINPUT23), .A3(G20), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G1956), .ZN(new_n766));
  INV_X1    g341(.A(G35), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n767), .A2(G29), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(KEYINPUT101), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n482), .B2(G29), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT102), .B(KEYINPUT29), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n769), .A2(KEYINPUT101), .ZN(new_n773));
  OR3_X1    g348(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n772), .B1(new_n771), .B2(new_n773), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n766), .B1(new_n776), .B2(G2090), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n776), .A2(G2090), .ZN(new_n778));
  INV_X1    g353(.A(G116), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n460), .B1(new_n779), .B2(G2105), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT94), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G104), .B2(G2105), .ZN(new_n782));
  INV_X1    g357(.A(G104), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n783), .A2(new_n467), .A3(KEYINPUT94), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n780), .A2(new_n782), .A3(new_n784), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT95), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n478), .A2(G128), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n480), .A2(G140), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(G29), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT96), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n698), .A2(G26), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT28), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(G2067), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n741), .A2(G5), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G171), .B2(new_n741), .ZN(new_n798));
  INV_X1    g373(.A(G1961), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n777), .A2(new_n778), .A3(new_n796), .A4(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n761), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(G16), .A2(G23), .ZN(new_n803));
  AND3_X1   g378(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(G16), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT33), .B(G1976), .Z(new_n806));
  OR2_X1    g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(G1971), .ZN(new_n808));
  NAND2_X1  g383(.A1(G303), .A2(G16), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n741), .A2(G22), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n810), .ZN(new_n812));
  AOI211_X1 g387(.A(G1971), .B(new_n812), .C1(G303), .C2(G16), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n805), .A2(new_n806), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n807), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT32), .B(G1981), .Z(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(G305), .A2(G16), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(G6), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n821), .A2(G16), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n818), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  OAI211_X1 g398(.A(new_n819), .B(new_n817), .C1(new_n821), .C2(G16), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(KEYINPUT34), .B1(new_n816), .B2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT89), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g403(.A(KEYINPUT89), .B(KEYINPUT34), .C1(new_n816), .C2(new_n825), .ZN(new_n829));
  AND2_X1   g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT90), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n831), .A2(KEYINPUT36), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT91), .Z(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n825), .ZN(new_n835));
  INV_X1    g410(.A(new_n806), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n805), .B(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT34), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n835), .A2(new_n837), .A3(new_n838), .A4(new_n814), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n741), .A2(G24), .ZN(new_n840));
  INV_X1    g415(.A(G290), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n840), .B1(new_n841), .B2(new_n741), .ZN(new_n842));
  XOR2_X1   g417(.A(KEYINPUT88), .B(G1986), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n831), .A2(KEYINPUT36), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n478), .A2(G119), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n480), .A2(G131), .ZN(new_n847));
  NOR2_X1   g422(.A1(G95), .A2(G2105), .ZN(new_n848));
  OAI21_X1  g423(.A(G2104), .B1(new_n467), .B2(G107), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n846), .B(new_n847), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  MUX2_X1   g425(.A(G25), .B(new_n850), .S(G29), .Z(new_n851));
  XNOR2_X1  g426(.A(KEYINPUT35), .B(G1991), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n851), .B(new_n852), .Z(new_n853));
  NAND4_X1  g428(.A1(new_n839), .A2(new_n844), .A3(new_n845), .A4(new_n853), .ZN(new_n854));
  NOR3_X1   g429(.A1(new_n830), .A2(new_n834), .A3(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n854), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n828), .A2(new_n829), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n833), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n694), .B(new_n802), .C1(new_n855), .C2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n702), .A2(G2078), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n713), .B1(G29), .B2(new_n716), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(new_n714), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n860), .A2(KEYINPUT103), .A3(new_n861), .A4(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT103), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n834), .B1(new_n830), .B2(new_n854), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n856), .A2(new_n833), .A3(new_n857), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND4_X1  g443(.A1(new_n868), .A2(new_n863), .A3(new_n694), .A4(new_n802), .ZN(new_n869));
  INV_X1    g444(.A(new_n861), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n865), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n864), .A2(new_n871), .ZN(G311));
  NAND3_X1  g447(.A1(new_n860), .A2(new_n861), .A3(new_n863), .ZN(G150));
  AOI22_X1  g448(.A1(new_n499), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n874), .A2(new_n501), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n499), .A2(new_n503), .A3(G93), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT104), .ZN(new_n877));
  OAI211_X1 g452(.A(G55), .B(G543), .C1(new_n510), .C2(new_n511), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n877), .B1(new_n876), .B2(new_n878), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n875), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(G860), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n883), .B(KEYINPUT37), .Z(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n550), .ZN(new_n885));
  OAI221_X1 g460(.A(new_n875), .B1(new_n546), .B2(new_n549), .C1(new_n880), .C2(new_n881), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  XOR2_X1   g462(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n888));
  XNOR2_X1  g463(.A(new_n887), .B(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n607), .A2(new_n615), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n889), .B(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n884), .B1(new_n891), .B2(G860), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(KEYINPUT105), .ZN(G145));
  XNOR2_X1  g468(.A(new_n622), .B(new_n850), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(G164), .A2(new_n789), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n497), .A2(new_n787), .A3(new_n786), .A4(new_n788), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(new_n710), .ZN(new_n899));
  INV_X1    g474(.A(new_n710), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n896), .A2(new_n900), .A3(new_n897), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n734), .A2(new_n711), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n478), .A2(G130), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n480), .A2(G142), .ZN(new_n906));
  OR2_X1    g481(.A1(G106), .A2(G2105), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n907), .B(G2104), .C1(G118), .C2(new_n467), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n905), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n734), .A2(KEYINPUT100), .ZN(new_n910));
  INV_X1    g485(.A(new_n730), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n910), .A2(new_n899), .A3(new_n911), .A4(new_n901), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n904), .A2(new_n909), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n909), .B1(new_n904), .B2(new_n912), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n895), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n915), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n917), .A2(new_n894), .A3(new_n913), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  OR2_X1    g494(.A1(new_n633), .A2(G160), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n633), .A2(G160), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(G162), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(G162), .B1(new_n920), .B2(new_n921), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT106), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n924), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(new_n927), .A3(new_n922), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n919), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT107), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n923), .A2(new_n924), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n916), .A2(new_n918), .A3(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(G37), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n919), .A2(KEYINPUT107), .A3(new_n930), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n933), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n939), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g515(.A(new_n887), .B(KEYINPUT108), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n941), .B(new_n617), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT78), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n536), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n499), .A2(KEYINPUT78), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n944), .A2(new_n945), .A3(G65), .ZN(new_n946));
  INV_X1    g521(.A(new_n567), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n501), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G91), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n949), .B1(new_n557), .B2(new_n559), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n562), .B(new_n563), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n948), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n607), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n605), .B1(new_n560), .B2(G92), .ZN(new_n954));
  INV_X1    g529(.A(G92), .ZN(new_n955));
  AOI211_X1 g530(.A(KEYINPUT10), .B(new_n955), .C1(new_n557), .C2(new_n559), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n604), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n944), .A2(new_n945), .A3(G66), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n959), .B1(new_n601), .B2(new_n506), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n958), .B1(new_n960), .B2(G651), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n957), .A2(G299), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n953), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n942), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n953), .A2(new_n962), .A3(KEYINPUT109), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT41), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT109), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n607), .A2(new_n967), .A3(new_n952), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n965), .A2(new_n966), .A3(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n953), .A2(new_n962), .A3(KEYINPUT41), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n964), .B1(new_n972), .B2(new_n942), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT110), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n973), .A2(new_n974), .A3(KEYINPUT42), .ZN(new_n975));
  XNOR2_X1  g550(.A(G288), .B(G303), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(G305), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(G290), .ZN(new_n978));
  OR2_X1    g553(.A1(new_n976), .A2(G305), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n976), .A2(G305), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n979), .A2(new_n841), .A3(new_n980), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT42), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n982), .B1(KEYINPUT110), .B2(new_n983), .ZN(new_n984));
  OAI221_X1 g559(.A(new_n964), .B1(KEYINPUT110), .B2(new_n983), .C1(new_n942), .C2(new_n972), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n975), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n984), .B1(new_n975), .B2(new_n985), .ZN(new_n987));
  OAI21_X1  g562(.A(G868), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n882), .A2(new_n611), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(G295));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n989), .ZN(G331));
  INV_X1    g566(.A(KEYINPUT111), .ZN(new_n992));
  INV_X1    g567(.A(G89), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n524), .B(new_n528), .C1(new_n512), .C2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT74), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(new_n529), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n997), .A2(G301), .A3(new_n517), .A4(new_n519), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  AOI22_X1  g574(.A1(new_n996), .A2(new_n529), .B1(G51), .B2(new_n518), .ZN(new_n1000));
  AOI21_X1  g575(.A(G301), .B1(new_n1000), .B2(new_n517), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n887), .B(new_n992), .C1(new_n999), .C2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n887), .B1(new_n999), .B2(new_n1001), .ZN(new_n1003));
  NAND2_X1  g578(.A1(G286), .A2(G171), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1004), .A2(new_n885), .A3(new_n886), .A4(new_n998), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1003), .A2(new_n1005), .A3(KEYINPUT111), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n971), .A2(new_n1002), .A3(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1003), .A2(new_n1005), .A3(KEYINPUT112), .ZN(new_n1008));
  INV_X1    g583(.A(new_n887), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT112), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1009), .A2(new_n1010), .A3(new_n998), .A4(new_n1004), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(new_n963), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1007), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT113), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1007), .A2(new_n1013), .A3(KEYINPUT113), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1016), .A2(new_n982), .A3(new_n1017), .ZN(new_n1018));
  AND2_X1   g593(.A1(new_n1007), .A2(new_n1013), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n978), .A2(new_n981), .ZN(new_n1020));
  AOI21_X1  g595(.A(G37), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT43), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1018), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n936), .B1(new_n1014), .B2(new_n982), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n963), .A2(new_n966), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT114), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n963), .A2(new_n1027), .A3(new_n966), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n966), .B1(new_n965), .B2(new_n968), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1011), .B(new_n1008), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1006), .A2(new_n1002), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n963), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1020), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT43), .B1(new_n1024), .B2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1023), .A2(KEYINPUT44), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1007), .A2(KEYINPUT113), .A3(new_n1013), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT113), .B1(new_n1007), .B2(new_n1013), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n1038), .A2(new_n1039), .A3(new_n1020), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT43), .B1(new_n1040), .B2(new_n1024), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1034), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1042), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT44), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1037), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1022), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1047));
  NOR3_X1   g622(.A1(new_n1024), .A2(new_n1034), .A3(KEYINPUT43), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1037), .B(new_n1045), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1036), .B1(new_n1046), .B2(new_n1050), .ZN(G397));
  NOR2_X1   g626(.A1(new_n789), .A2(G2067), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n789), .A2(G2067), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n710), .A2(G1996), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G1384), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n497), .A2(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g633(.A(KEYINPUT116), .B(KEYINPUT45), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G40), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n468), .A2(new_n472), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1061), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1056), .A2(new_n1065), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n1061), .A2(new_n1064), .A3(G1996), .ZN(new_n1067));
  XNOR2_X1  g642(.A(new_n1067), .B(KEYINPUT117), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1066), .B1(new_n1068), .B2(new_n712), .ZN(new_n1069));
  OR2_X1    g644(.A1(new_n1069), .A2(KEYINPUT118), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(KEYINPUT118), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n850), .A2(new_n852), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n850), .A2(new_n852), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1065), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1070), .A2(new_n1071), .A3(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g650(.A(G290), .B(G1986), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1075), .B1(new_n1065), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G1966), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1063), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT45), .B1(new_n497), .B2(new_n1057), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1078), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n497), .A2(KEYINPUT50), .A3(new_n1057), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT50), .B1(new_n497), .B2(new_n1057), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n693), .B(new_n1063), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1081), .A2(KEYINPUT123), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT123), .B1(new_n1081), .B2(new_n1085), .ZN(new_n1087));
  NOR3_X1   g662(.A1(new_n1086), .A2(new_n1087), .A3(G286), .ZN(new_n1088));
  INV_X1    g663(.A(G8), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT51), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1087), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1081), .A2(KEYINPUT123), .A3(new_n1085), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1091), .A2(KEYINPUT51), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1081), .A2(new_n1085), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(G168), .B1(new_n1095), .B2(KEYINPUT51), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1093), .A2(new_n1096), .A3(G8), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT62), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1090), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n1057), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n1061), .A2(new_n1063), .A3(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1063), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1102));
  XNOR2_X1  g677(.A(KEYINPUT119), .B(G2090), .ZN(new_n1103));
  OAI22_X1  g678(.A1(new_n1101), .A2(G1971), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT55), .ZN(new_n1105));
  NAND3_X1  g680(.A1(G303), .A2(new_n1105), .A3(G8), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1105), .B1(G303), .B2(G8), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT120), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1108), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1110), .A2(new_n1111), .A3(new_n1106), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1109), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1104), .A2(G8), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT53), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1061), .A2(new_n1063), .A3(new_n1100), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1116), .B1(new_n1117), .B2(G2078), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1102), .A2(new_n799), .ZN(new_n1119));
  OR2_X1    g694(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1120));
  OR2_X1    g695(.A1(new_n1116), .A2(G2078), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1118), .B(new_n1119), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(G171), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1104), .A2(G8), .B1(new_n1110), .B2(new_n1106), .ZN(new_n1124));
  OR2_X1    g699(.A1(G305), .A2(G1981), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n586), .A2(new_n582), .A3(new_n585), .ZN(new_n1126));
  INV_X1    g701(.A(G86), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n512), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(G1981), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1125), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT49), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1063), .A2(new_n1057), .A3(new_n497), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(G8), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1125), .A2(KEYINPUT49), .A3(new_n1129), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1132), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(G1976), .ZN(new_n1138));
  AOI21_X1  g713(.A(KEYINPUT52), .B1(G288), .B2(new_n1138), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1135), .B(new_n1139), .C1(new_n1138), .C2(G288), .ZN(new_n1140));
  NOR2_X1   g715(.A1(G288), .A2(new_n1138), .ZN(new_n1141));
  OAI21_X1  g716(.A(KEYINPUT52), .B1(new_n1134), .B2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1137), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1143));
  NOR4_X1   g718(.A1(new_n1115), .A2(new_n1123), .A3(new_n1124), .A4(new_n1143), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1099), .A2(new_n1144), .A3(KEYINPUT126), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT126), .B1(new_n1099), .B2(new_n1144), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1098), .B1(new_n1090), .B2(new_n1097), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT63), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1124), .ZN(new_n1150));
  AND3_X1   g725(.A1(new_n1137), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1150), .A2(new_n1151), .A3(G168), .A4(new_n1114), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1095), .A2(new_n1089), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1149), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  NOR3_X1   g730(.A1(new_n1115), .A2(new_n1124), .A3(new_n1143), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1156), .A2(KEYINPUT63), .A3(G168), .A4(new_n1153), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1137), .A2(new_n1138), .A3(new_n804), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1134), .B1(new_n1159), .B2(new_n1125), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1160), .B1(new_n1115), .B2(new_n1151), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT50), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1058), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1064), .B1(new_n1163), .B2(new_n1082), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1164), .A2(G1956), .ZN(new_n1165));
  XNOR2_X1  g740(.A(KEYINPUT56), .B(G2072), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1117), .A2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1165), .A2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n948), .A2(new_n950), .ZN(new_n1170));
  AOI21_X1  g745(.A(KEYINPUT57), .B1(new_n1170), .B2(KEYINPUT121), .ZN(new_n1171));
  OR2_X1    g746(.A1(new_n1171), .A2(G299), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(G299), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1169), .A2(new_n1174), .ZN(new_n1175));
  OAI211_X1 g750(.A(new_n1172), .B(new_n1173), .C1(new_n1165), .C2(new_n1168), .ZN(new_n1176));
  OAI22_X1  g751(.A1(new_n1164), .A2(G1348), .B1(G2067), .B2(new_n1133), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(new_n608), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1175), .A2(new_n1176), .A3(KEYINPUT61), .A4(new_n1178), .ZN(new_n1179));
  AND2_X1   g754(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1180));
  XOR2_X1   g755(.A(G301), .B(KEYINPUT54), .Z(new_n1181));
  XNOR2_X1  g756(.A(KEYINPUT125), .B(G2078), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1100), .A2(KEYINPUT53), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n1184), .B(KEYINPUT124), .ZN(new_n1185));
  OAI211_X1 g760(.A(new_n1180), .B(new_n1181), .C1(new_n1183), .C2(new_n1185), .ZN(new_n1186));
  AND2_X1   g761(.A1(new_n1179), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1177), .A2(new_n607), .ZN(new_n1188));
  OAI221_X1 g763(.A(new_n608), .B1(G2067), .B2(new_n1133), .C1(new_n1164), .C2(G1348), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1188), .A2(new_n1189), .A3(KEYINPUT60), .ZN(new_n1190));
  OR3_X1    g765(.A1(new_n1177), .A2(KEYINPUT60), .A3(new_n607), .ZN(new_n1191));
  INV_X1    g766(.A(new_n1133), .ZN(new_n1192));
  XNOR2_X1  g767(.A(KEYINPUT58), .B(G1341), .ZN(new_n1193));
  OAI22_X1  g768(.A1(new_n1117), .A2(G1996), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1194), .A2(new_n550), .ZN(new_n1195));
  OR2_X1    g770(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1196));
  NAND2_X1  g771(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  NAND4_X1  g773(.A1(new_n1194), .A2(KEYINPUT122), .A3(KEYINPUT59), .A4(new_n550), .ZN(new_n1199));
  NAND4_X1  g774(.A1(new_n1190), .A2(new_n1191), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1201), .A2(new_n1175), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(new_n1181), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1122), .A2(new_n1204), .ZN(new_n1205));
  OR2_X1    g780(.A1(new_n1175), .A2(KEYINPUT61), .ZN(new_n1206));
  NAND4_X1  g781(.A1(new_n1187), .A2(new_n1203), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1090), .A2(new_n1097), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1208), .A2(new_n1156), .ZN(new_n1209));
  OAI211_X1 g784(.A(new_n1158), .B(new_n1161), .C1(new_n1207), .C2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g785(.A(new_n1077), .B1(new_n1148), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT127), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1075), .A2(new_n1212), .ZN(new_n1213));
  NOR4_X1   g788(.A1(new_n1061), .A2(new_n1064), .A3(G1986), .A4(G290), .ZN(new_n1214));
  XOR2_X1   g789(.A(new_n1214), .B(KEYINPUT48), .Z(new_n1215));
  NAND4_X1  g790(.A1(new_n1070), .A2(KEYINPUT127), .A3(new_n1071), .A4(new_n1074), .ZN(new_n1216));
  NAND3_X1  g791(.A1(new_n1213), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1054), .A2(new_n900), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n1065), .B1(new_n1052), .B2(new_n1218), .ZN(new_n1219));
  AND2_X1   g794(.A1(new_n1068), .A2(KEYINPUT46), .ZN(new_n1220));
  NOR2_X1   g795(.A1(new_n1068), .A2(KEYINPUT46), .ZN(new_n1221));
  OAI21_X1  g796(.A(new_n1219), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  XNOR2_X1  g797(.A(new_n1222), .B(KEYINPUT47), .ZN(new_n1223));
  AND3_X1   g798(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1224));
  OAI21_X1  g799(.A(new_n1065), .B1(new_n1224), .B2(new_n1052), .ZN(new_n1225));
  AND3_X1   g800(.A1(new_n1217), .A2(new_n1223), .A3(new_n1225), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1211), .A2(new_n1226), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g802(.A1(new_n685), .A2(G319), .A3(new_n1044), .ZN(new_n1229));
  NAND3_X1  g803(.A1(new_n939), .A2(new_n650), .A3(new_n663), .ZN(new_n1230));
  NOR2_X1   g804(.A1(new_n1229), .A2(new_n1230), .ZN(G308));
  NAND2_X1  g805(.A1(new_n650), .A2(new_n663), .ZN(new_n1232));
  AOI21_X1  g806(.A(KEYINPUT107), .B1(new_n919), .B2(new_n930), .ZN(new_n1233));
  AOI211_X1 g807(.A(new_n932), .B(new_n929), .C1(new_n916), .C2(new_n918), .ZN(new_n1234));
  NOR2_X1   g808(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g809(.A(new_n1232), .B1(new_n1235), .B2(new_n937), .ZN(new_n1236));
  NAND4_X1  g810(.A1(new_n1236), .A2(G319), .A3(new_n685), .A4(new_n1044), .ZN(G225));
endmodule


