

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U555 ( .A1(n654), .A2(n653), .ZN(n655) );
  AND2_X1 U556 ( .A1(n651), .A2(n526), .ZN(n652) );
  BUF_X1 U557 ( .A(n722), .Z(n723) );
  AND2_X2 U558 ( .A1(n531), .A2(G2105), .ZN(n999) );
  AND2_X2 U559 ( .A1(G2104), .A2(G2105), .ZN(n998) );
  INV_X1 U560 ( .A(KEYINPUT103), .ZN(n678) );
  NAND2_X1 U561 ( .A1(n718), .A2(n717), .ZN(n719) );
  AND2_X1 U562 ( .A1(n525), .A2(n755), .ZN(n521) );
  AND2_X1 U563 ( .A1(G113), .A2(n998), .ZN(n522) );
  AND2_X1 U564 ( .A1(G125), .A2(n999), .ZN(n523) );
  AND2_X1 U565 ( .A1(n697), .A2(n696), .ZN(n524) );
  AND2_X1 U566 ( .A1(n764), .A2(n754), .ZN(n525) );
  NAND2_X1 U567 ( .A1(n911), .A2(n650), .ZN(n526) );
  XOR2_X1 U568 ( .A(KEYINPUT97), .B(n609), .Z(n527) );
  AND2_X1 U569 ( .A1(n657), .A2(G1996), .ZN(n634) );
  INV_X1 U570 ( .A(KEYINPUT98), .ZN(n642) );
  BUF_X1 U571 ( .A(n637), .Z(n672) );
  INV_X1 U572 ( .A(KEYINPUT94), .ZN(n594) );
  NAND2_X1 U573 ( .A1(n595), .A2(n721), .ZN(n637) );
  AND2_X1 U574 ( .A1(n775), .A2(G40), .ZN(n591) );
  INV_X1 U575 ( .A(KEYINPUT74), .ZN(n625) );
  AND2_X1 U576 ( .A1(n591), .A2(n772), .ZN(n593) );
  XNOR2_X1 U577 ( .A(n625), .B(KEYINPUT13), .ZN(n626) );
  NOR2_X1 U578 ( .A1(G164), .A2(G1384), .ZN(n721) );
  XNOR2_X1 U579 ( .A(KEYINPUT67), .B(G651), .ZN(n540) );
  XNOR2_X1 U580 ( .A(n627), .B(n626), .ZN(n628) );
  XOR2_X1 U581 ( .A(G543), .B(KEYINPUT0), .Z(n578) );
  NOR2_X2 U582 ( .A1(G2104), .A2(G2105), .ZN(n528) );
  XOR2_X2 U583 ( .A(KEYINPUT17), .B(n528), .Z(n722) );
  NAND2_X1 U584 ( .A1(G138), .A2(n722), .ZN(n530) );
  INV_X1 U585 ( .A(G2104), .ZN(n531) );
  NOR2_X1 U586 ( .A1(G2105), .A2(n531), .ZN(n589) );
  BUF_X1 U587 ( .A(n589), .Z(n1003) );
  NAND2_X1 U588 ( .A1(G102), .A2(n1003), .ZN(n529) );
  NAND2_X1 U589 ( .A1(n530), .A2(n529), .ZN(n535) );
  NAND2_X1 U590 ( .A1(G114), .A2(n998), .ZN(n533) );
  NAND2_X1 U591 ( .A1(G126), .A2(n999), .ZN(n532) );
  NAND2_X1 U592 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U593 ( .A1(n535), .A2(n534), .ZN(G164) );
  NOR2_X1 U594 ( .A1(G543), .A2(n540), .ZN(n536) );
  XOR2_X1 U595 ( .A(KEYINPUT1), .B(n536), .Z(n617) );
  BUF_X1 U596 ( .A(n617), .Z(n808) );
  NAND2_X1 U597 ( .A1(n808), .A2(G61), .ZN(n537) );
  XNOR2_X1 U598 ( .A(n537), .B(KEYINPUT82), .ZN(n545) );
  NOR2_X2 U599 ( .A1(G651), .A2(n578), .ZN(n806) );
  NAND2_X1 U600 ( .A1(G48), .A2(n806), .ZN(n539) );
  NOR2_X1 U601 ( .A1(G543), .A2(G651), .ZN(n619) );
  BUF_X1 U602 ( .A(n619), .Z(n802) );
  NAND2_X1 U603 ( .A1(G86), .A2(n802), .ZN(n538) );
  NAND2_X1 U604 ( .A1(n539), .A2(n538), .ZN(n543) );
  NOR2_X2 U605 ( .A1(n578), .A2(n540), .ZN(n803) );
  NAND2_X1 U606 ( .A1(n803), .A2(G73), .ZN(n541) );
  XOR2_X1 U607 ( .A(KEYINPUT2), .B(n541), .Z(n542) );
  NOR2_X1 U608 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U609 ( .A1(n545), .A2(n544), .ZN(G305) );
  NAND2_X1 U610 ( .A1(n806), .A2(G52), .ZN(n547) );
  NAND2_X1 U611 ( .A1(G64), .A2(n808), .ZN(n546) );
  NAND2_X1 U612 ( .A1(n547), .A2(n546), .ZN(n553) );
  NAND2_X1 U613 ( .A1(n802), .A2(G90), .ZN(n549) );
  NAND2_X1 U614 ( .A1(G77), .A2(n803), .ZN(n548) );
  NAND2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U616 ( .A(KEYINPUT9), .B(n550), .ZN(n551) );
  XNOR2_X1 U617 ( .A(KEYINPUT69), .B(n551), .ZN(n552) );
  NOR2_X1 U618 ( .A1(n553), .A2(n552), .ZN(G171) );
  INV_X1 U619 ( .A(G171), .ZN(G301) );
  NAND2_X1 U620 ( .A1(n806), .A2(G51), .ZN(n555) );
  NAND2_X1 U621 ( .A1(G63), .A2(n808), .ZN(n554) );
  NAND2_X1 U622 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(KEYINPUT6), .B(n556), .ZN(n563) );
  NAND2_X1 U624 ( .A1(G89), .A2(n802), .ZN(n557) );
  XOR2_X1 U625 ( .A(KEYINPUT4), .B(n557), .Z(n558) );
  XNOR2_X1 U626 ( .A(n558), .B(KEYINPUT75), .ZN(n560) );
  NAND2_X1 U627 ( .A1(G76), .A2(n803), .ZN(n559) );
  NAND2_X1 U628 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U629 ( .A(n561), .B(KEYINPUT5), .Z(n562) );
  NOR2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U631 ( .A(KEYINPUT76), .B(n564), .Z(n565) );
  XNOR2_X1 U632 ( .A(KEYINPUT7), .B(n565), .ZN(G168) );
  XOR2_X1 U633 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U634 ( .A1(n803), .A2(G75), .ZN(n566) );
  XNOR2_X1 U635 ( .A(n566), .B(KEYINPUT84), .ZN(n573) );
  NAND2_X1 U636 ( .A1(n806), .A2(G50), .ZN(n568) );
  NAND2_X1 U637 ( .A1(G62), .A2(n808), .ZN(n567) );
  NAND2_X1 U638 ( .A1(n568), .A2(n567), .ZN(n571) );
  NAND2_X1 U639 ( .A1(G88), .A2(n802), .ZN(n569) );
  XNOR2_X1 U640 ( .A(KEYINPUT83), .B(n569), .ZN(n570) );
  NOR2_X1 U641 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U642 ( .A1(n573), .A2(n572), .ZN(G303) );
  NAND2_X1 U643 ( .A1(G49), .A2(n806), .ZN(n575) );
  NAND2_X1 U644 ( .A1(G74), .A2(G651), .ZN(n574) );
  NAND2_X1 U645 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U646 ( .A1(n808), .A2(n576), .ZN(n577) );
  XOR2_X1 U647 ( .A(KEYINPUT81), .B(n577), .Z(n580) );
  NAND2_X1 U648 ( .A1(n578), .A2(G87), .ZN(n579) );
  NAND2_X1 U649 ( .A1(n580), .A2(n579), .ZN(G288) );
  NAND2_X1 U650 ( .A1(n806), .A2(G47), .ZN(n582) );
  NAND2_X1 U651 ( .A1(G60), .A2(n808), .ZN(n581) );
  NAND2_X1 U652 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U653 ( .A(KEYINPUT68), .B(n583), .Z(n587) );
  NAND2_X1 U654 ( .A1(n803), .A2(G72), .ZN(n585) );
  NAND2_X1 U655 ( .A1(n802), .A2(G85), .ZN(n584) );
  AND2_X1 U656 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U657 ( .A1(n587), .A2(n586), .ZN(G290) );
  NOR2_X1 U658 ( .A1(G1981), .A2(G305), .ZN(n588) );
  XNOR2_X1 U659 ( .A(KEYINPUT24), .B(n588), .ZN(n597) );
  NOR2_X1 U660 ( .A1(n522), .A2(n523), .ZN(n775) );
  NAND2_X1 U661 ( .A1(G101), .A2(n589), .ZN(n590) );
  XOR2_X1 U662 ( .A(KEYINPUT23), .B(n590), .Z(n772) );
  NAND2_X1 U663 ( .A1(G137), .A2(n722), .ZN(n592) );
  XNOR2_X1 U664 ( .A(n592), .B(KEYINPUT66), .ZN(n773) );
  NAND2_X1 U665 ( .A1(n593), .A2(n773), .ZN(n720) );
  XNOR2_X1 U666 ( .A(n720), .B(n594), .ZN(n595) );
  NAND2_X1 U667 ( .A1(G8), .A2(n637), .ZN(n596) );
  XNOR2_X1 U668 ( .A(KEYINPUT95), .B(n596), .ZN(n711) );
  NAND2_X1 U669 ( .A1(n597), .A2(n711), .ZN(n697) );
  INV_X1 U670 ( .A(n711), .ZN(n695) );
  NAND2_X1 U671 ( .A1(n806), .A2(G53), .ZN(n599) );
  NAND2_X1 U672 ( .A1(G65), .A2(n808), .ZN(n598) );
  NAND2_X1 U673 ( .A1(n599), .A2(n598), .ZN(n603) );
  NAND2_X1 U674 ( .A1(n802), .A2(G91), .ZN(n601) );
  NAND2_X1 U675 ( .A1(G78), .A2(n803), .ZN(n600) );
  NAND2_X1 U676 ( .A1(n601), .A2(n600), .ZN(n602) );
  NOR2_X1 U677 ( .A1(n603), .A2(n602), .ZN(n911) );
  INV_X1 U678 ( .A(KEYINPUT96), .ZN(n604) );
  XNOR2_X1 U679 ( .A(n604), .B(n637), .ZN(n636) );
  NAND2_X1 U680 ( .A1(G2072), .A2(n636), .ZN(n605) );
  XNOR2_X1 U681 ( .A(n605), .B(KEYINPUT27), .ZN(n608) );
  INV_X1 U682 ( .A(n636), .ZN(n656) );
  INV_X1 U683 ( .A(n656), .ZN(n606) );
  INV_X1 U684 ( .A(G1956), .ZN(n910) );
  NOR2_X1 U685 ( .A1(n606), .A2(n910), .ZN(n607) );
  NOR2_X1 U686 ( .A1(n608), .A2(n607), .ZN(n650) );
  NOR2_X1 U687 ( .A1(n911), .A2(n650), .ZN(n609) );
  XNOR2_X1 U688 ( .A(KEYINPUT28), .B(n527), .ZN(n654) );
  NAND2_X1 U689 ( .A1(G54), .A2(n806), .ZN(n611) );
  NAND2_X1 U690 ( .A1(G92), .A2(n802), .ZN(n610) );
  NAND2_X1 U691 ( .A1(n611), .A2(n610), .ZN(n615) );
  NAND2_X1 U692 ( .A1(G66), .A2(n617), .ZN(n613) );
  NAND2_X1 U693 ( .A1(G79), .A2(n803), .ZN(n612) );
  NAND2_X1 U694 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X2 U695 ( .A1(n615), .A2(n614), .ZN(n616) );
  XOR2_X2 U696 ( .A(KEYINPUT15), .B(n616), .Z(n1019) );
  AND2_X1 U697 ( .A1(n637), .A2(G1341), .ZN(n632) );
  NAND2_X1 U698 ( .A1(G56), .A2(n617), .ZN(n618) );
  XOR2_X1 U699 ( .A(KEYINPUT14), .B(n618), .Z(n629) );
  NAND2_X1 U700 ( .A1(n803), .A2(G68), .ZN(n624) );
  XOR2_X1 U701 ( .A(KEYINPUT12), .B(KEYINPUT73), .Z(n621) );
  NAND2_X1 U702 ( .A1(G81), .A2(n619), .ZN(n620) );
  XNOR2_X1 U703 ( .A(n621), .B(n620), .ZN(n622) );
  XNOR2_X1 U704 ( .A(KEYINPUT72), .B(n622), .ZN(n623) );
  NAND2_X1 U705 ( .A1(n624), .A2(n623), .ZN(n627) );
  NOR2_X1 U706 ( .A1(n629), .A2(n628), .ZN(n631) );
  NAND2_X1 U707 ( .A1(n806), .A2(G43), .ZN(n630) );
  NAND2_X1 U708 ( .A1(n631), .A2(n630), .ZN(n784) );
  NOR2_X1 U709 ( .A1(n632), .A2(n784), .ZN(n644) );
  AND2_X1 U710 ( .A1(n1019), .A2(n644), .ZN(n635) );
  INV_X1 U711 ( .A(n637), .ZN(n657) );
  XNOR2_X1 U712 ( .A(KEYINPUT65), .B(KEYINPUT26), .ZN(n633) );
  XNOR2_X1 U713 ( .A(n634), .B(n633), .ZN(n645) );
  NAND2_X1 U714 ( .A1(n635), .A2(n645), .ZN(n641) );
  NAND2_X1 U715 ( .A1(n636), .A2(G2067), .ZN(n639) );
  NAND2_X1 U716 ( .A1(G1348), .A2(n672), .ZN(n638) );
  NAND2_X1 U717 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U718 ( .A1(n641), .A2(n640), .ZN(n643) );
  XNOR2_X1 U719 ( .A(n643), .B(n642), .ZN(n648) );
  AND2_X1 U720 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U721 ( .A1(n1019), .A2(n646), .ZN(n647) );
  NOR2_X1 U722 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U723 ( .A(n649), .B(KEYINPUT99), .ZN(n651) );
  XNOR2_X1 U724 ( .A(n652), .B(KEYINPUT100), .ZN(n653) );
  XNOR2_X1 U725 ( .A(n655), .B(KEYINPUT29), .ZN(n661) );
  XOR2_X1 U726 ( .A(G2078), .B(KEYINPUT25), .Z(n853) );
  NOR2_X1 U727 ( .A1(n853), .A2(n656), .ZN(n659) );
  NOR2_X1 U728 ( .A1(n657), .A2(G1961), .ZN(n658) );
  NOR2_X1 U729 ( .A1(n659), .A2(n658), .ZN(n666) );
  OR2_X1 U730 ( .A1(G301), .A2(n666), .ZN(n660) );
  NAND2_X1 U731 ( .A1(n661), .A2(n660), .ZN(n671) );
  NOR2_X1 U732 ( .A1(G2084), .A2(n672), .ZN(n686) );
  NOR2_X1 U733 ( .A1(G1966), .A2(n695), .ZN(n682) );
  NOR2_X1 U734 ( .A1(n686), .A2(n682), .ZN(n662) );
  NAND2_X1 U735 ( .A1(G8), .A2(n662), .ZN(n663) );
  XNOR2_X1 U736 ( .A(KEYINPUT30), .B(n663), .ZN(n664) );
  NOR2_X1 U737 ( .A1(G168), .A2(n664), .ZN(n665) );
  XNOR2_X1 U738 ( .A(n665), .B(KEYINPUT101), .ZN(n668) );
  NAND2_X1 U739 ( .A1(n666), .A2(G301), .ZN(n667) );
  NAND2_X1 U740 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U741 ( .A(n669), .B(KEYINPUT31), .ZN(n670) );
  NAND2_X1 U742 ( .A1(n671), .A2(n670), .ZN(n683) );
  NAND2_X1 U743 ( .A1(n683), .A2(G286), .ZN(n677) );
  NOR2_X1 U744 ( .A1(G1971), .A2(n695), .ZN(n674) );
  NOR2_X1 U745 ( .A1(G2090), .A2(n672), .ZN(n673) );
  NOR2_X1 U746 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U747 ( .A1(n675), .A2(G303), .ZN(n676) );
  NAND2_X1 U748 ( .A1(n677), .A2(n676), .ZN(n679) );
  XNOR2_X1 U749 ( .A(n679), .B(n678), .ZN(n680) );
  NAND2_X1 U750 ( .A1(n680), .A2(G8), .ZN(n681) );
  XNOR2_X1 U751 ( .A(n681), .B(KEYINPUT32), .ZN(n700) );
  BUF_X1 U752 ( .A(n700), .Z(n689) );
  INV_X1 U753 ( .A(n682), .ZN(n684) );
  AND2_X1 U754 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U755 ( .A(n685), .B(KEYINPUT102), .ZN(n688) );
  NAND2_X1 U756 ( .A1(n686), .A2(G8), .ZN(n687) );
  NAND2_X1 U757 ( .A1(n688), .A2(n687), .ZN(n698) );
  NAND2_X1 U758 ( .A1(n689), .A2(n698), .ZN(n692) );
  NOR2_X1 U759 ( .A1(G2090), .A2(G303), .ZN(n690) );
  NAND2_X1 U760 ( .A1(G8), .A2(n690), .ZN(n691) );
  NAND2_X1 U761 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U762 ( .A(KEYINPUT107), .B(n693), .Z(n694) );
  NAND2_X1 U763 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U764 ( .A1(G1976), .A2(G288), .ZN(n914) );
  AND2_X1 U765 ( .A1(n698), .A2(n914), .ZN(n699) );
  NAND2_X1 U766 ( .A1(n700), .A2(n699), .ZN(n706) );
  INV_X1 U767 ( .A(n914), .ZN(n704) );
  NOR2_X1 U768 ( .A1(G1971), .A2(G303), .ZN(n702) );
  NOR2_X1 U769 ( .A1(G288), .A2(G1976), .ZN(n701) );
  XNOR2_X1 U770 ( .A(n701), .B(KEYINPUT104), .ZN(n909) );
  NOR2_X1 U771 ( .A1(n702), .A2(n909), .ZN(n703) );
  OR2_X1 U772 ( .A1(n704), .A2(n703), .ZN(n705) );
  AND2_X1 U773 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U774 ( .A(n707), .B(KEYINPUT105), .ZN(n708) );
  NAND2_X1 U775 ( .A1(n708), .A2(n711), .ZN(n709) );
  XNOR2_X1 U776 ( .A(n709), .B(KEYINPUT64), .ZN(n710) );
  INV_X1 U777 ( .A(KEYINPUT33), .ZN(n713) );
  NAND2_X1 U778 ( .A1(n710), .A2(n713), .ZN(n718) );
  XNOR2_X1 U779 ( .A(G1981), .B(G305), .ZN(n923) );
  INV_X1 U780 ( .A(n923), .ZN(n716) );
  NAND2_X1 U781 ( .A1(n711), .A2(n909), .ZN(n712) );
  NOR2_X1 U782 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U783 ( .A(n714), .B(KEYINPUT106), .Z(n715) );
  AND2_X1 U784 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U785 ( .A1(n524), .A2(n719), .ZN(n756) );
  NOR2_X1 U786 ( .A1(n721), .A2(n720), .ZN(n767) );
  NAND2_X1 U787 ( .A1(G140), .A2(n723), .ZN(n725) );
  NAND2_X1 U788 ( .A1(G104), .A2(n1003), .ZN(n724) );
  NAND2_X1 U789 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U790 ( .A(KEYINPUT34), .B(n726), .ZN(n732) );
  NAND2_X1 U791 ( .A1(G116), .A2(n998), .ZN(n728) );
  NAND2_X1 U792 ( .A1(G128), .A2(n999), .ZN(n727) );
  NAND2_X1 U793 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U794 ( .A(KEYINPUT88), .B(n729), .Z(n730) );
  XNOR2_X1 U795 ( .A(KEYINPUT35), .B(n730), .ZN(n731) );
  NOR2_X1 U796 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U797 ( .A(KEYINPUT36), .B(n733), .ZN(n995) );
  XNOR2_X1 U798 ( .A(G2067), .B(KEYINPUT37), .ZN(n757) );
  NOR2_X1 U799 ( .A1(n995), .A2(n757), .ZN(n890) );
  NAND2_X1 U800 ( .A1(n767), .A2(n890), .ZN(n764) );
  NAND2_X1 U801 ( .A1(G131), .A2(n723), .ZN(n735) );
  NAND2_X1 U802 ( .A1(G95), .A2(n1003), .ZN(n734) );
  NAND2_X1 U803 ( .A1(n735), .A2(n734), .ZN(n739) );
  NAND2_X1 U804 ( .A1(G107), .A2(n998), .ZN(n737) );
  NAND2_X1 U805 ( .A1(G119), .A2(n999), .ZN(n736) );
  NAND2_X1 U806 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U807 ( .A1(n739), .A2(n738), .ZN(n993) );
  XNOR2_X1 U808 ( .A(G1991), .B(KEYINPUT89), .ZN(n858) );
  NOR2_X1 U809 ( .A1(n993), .A2(n858), .ZN(n752) );
  NAND2_X1 U810 ( .A1(n998), .A2(G117), .ZN(n740) );
  XNOR2_X1 U811 ( .A(KEYINPUT91), .B(n740), .ZN(n743) );
  NAND2_X1 U812 ( .A1(n999), .A2(G129), .ZN(n741) );
  XOR2_X1 U813 ( .A(KEYINPUT90), .B(n741), .Z(n742) );
  NOR2_X1 U814 ( .A1(n743), .A2(n742), .ZN(n744) );
  XOR2_X1 U815 ( .A(KEYINPUT92), .B(n744), .Z(n748) );
  NAND2_X1 U816 ( .A1(G105), .A2(n1003), .ZN(n745) );
  XNOR2_X1 U817 ( .A(n745), .B(KEYINPUT93), .ZN(n746) );
  XNOR2_X1 U818 ( .A(KEYINPUT38), .B(n746), .ZN(n747) );
  NOR2_X1 U819 ( .A1(n748), .A2(n747), .ZN(n750) );
  NAND2_X1 U820 ( .A1(n723), .A2(G141), .ZN(n749) );
  NAND2_X1 U821 ( .A1(n750), .A2(n749), .ZN(n994) );
  AND2_X1 U822 ( .A1(n994), .A2(G1996), .ZN(n751) );
  NOR2_X1 U823 ( .A1(n752), .A2(n751), .ZN(n898) );
  INV_X1 U824 ( .A(n767), .ZN(n753) );
  NOR2_X1 U825 ( .A1(n898), .A2(n753), .ZN(n760) );
  INV_X1 U826 ( .A(n760), .ZN(n754) );
  XNOR2_X1 U827 ( .A(G1986), .B(G290), .ZN(n917) );
  NAND2_X1 U828 ( .A1(n917), .A2(n767), .ZN(n755) );
  NAND2_X1 U829 ( .A1(n756), .A2(n521), .ZN(n770) );
  NAND2_X1 U830 ( .A1(n995), .A2(n757), .ZN(n900) );
  NOR2_X1 U831 ( .A1(G1996), .A2(n994), .ZN(n893) );
  AND2_X1 U832 ( .A1(n858), .A2(n993), .ZN(n887) );
  NOR2_X1 U833 ( .A1(G1986), .A2(G290), .ZN(n758) );
  NOR2_X1 U834 ( .A1(n887), .A2(n758), .ZN(n759) );
  NOR2_X1 U835 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U836 ( .A1(n893), .A2(n761), .ZN(n762) );
  XNOR2_X1 U837 ( .A(KEYINPUT39), .B(n762), .ZN(n763) );
  XNOR2_X1 U838 ( .A(n763), .B(KEYINPUT108), .ZN(n765) );
  NAND2_X1 U839 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U840 ( .A1(n900), .A2(n766), .ZN(n768) );
  NAND2_X1 U841 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U842 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U843 ( .A(n771), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U844 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U845 ( .A1(n775), .A2(n774), .ZN(G160) );
  AND2_X1 U846 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U847 ( .A1(G135), .A2(n723), .ZN(n777) );
  NAND2_X1 U848 ( .A1(G111), .A2(n998), .ZN(n776) );
  NAND2_X1 U849 ( .A1(n777), .A2(n776), .ZN(n780) );
  NAND2_X1 U850 ( .A1(n999), .A2(G123), .ZN(n778) );
  XOR2_X1 U851 ( .A(KEYINPUT18), .B(n778), .Z(n779) );
  NOR2_X1 U852 ( .A1(n780), .A2(n779), .ZN(n782) );
  NAND2_X1 U853 ( .A1(n1003), .A2(G99), .ZN(n781) );
  NAND2_X1 U854 ( .A1(n782), .A2(n781), .ZN(n1013) );
  XNOR2_X1 U855 ( .A(G2096), .B(n1013), .ZN(n783) );
  OR2_X1 U856 ( .A1(G2100), .A2(n783), .ZN(G156) );
  BUF_X1 U857 ( .A(n784), .Z(n1022) );
  INV_X1 U858 ( .A(G860), .ZN(n793) );
  OR2_X1 U859 ( .A1(n1022), .A2(n793), .ZN(G153) );
  INV_X1 U860 ( .A(G57), .ZN(G237) );
  XOR2_X1 U861 ( .A(KEYINPUT71), .B(KEYINPUT10), .Z(n786) );
  NAND2_X1 U862 ( .A1(G7), .A2(G661), .ZN(n785) );
  XNOR2_X1 U863 ( .A(n786), .B(n785), .ZN(G223) );
  INV_X1 U864 ( .A(G223), .ZN(n840) );
  NAND2_X1 U865 ( .A1(n840), .A2(G567), .ZN(n787) );
  XOR2_X1 U866 ( .A(KEYINPUT11), .B(n787), .Z(G234) );
  NAND2_X1 U867 ( .A1(G868), .A2(G301), .ZN(n789) );
  OR2_X1 U868 ( .A1(n1019), .A2(G868), .ZN(n788) );
  NAND2_X1 U869 ( .A1(n789), .A2(n788), .ZN(G284) );
  XOR2_X1 U870 ( .A(KEYINPUT70), .B(n911), .Z(G299) );
  NAND2_X1 U871 ( .A1(G868), .A2(G286), .ZN(n792) );
  INV_X1 U872 ( .A(G868), .ZN(n790) );
  NAND2_X1 U873 ( .A1(G299), .A2(n790), .ZN(n791) );
  NAND2_X1 U874 ( .A1(n792), .A2(n791), .ZN(G297) );
  NAND2_X1 U875 ( .A1(n793), .A2(G559), .ZN(n794) );
  NAND2_X1 U876 ( .A1(n794), .A2(n1019), .ZN(n795) );
  XNOR2_X1 U877 ( .A(n795), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U878 ( .A1(G868), .A2(n1022), .ZN(n798) );
  NAND2_X1 U879 ( .A1(G868), .A2(n1019), .ZN(n796) );
  NOR2_X1 U880 ( .A1(G559), .A2(n796), .ZN(n797) );
  NOR2_X1 U881 ( .A1(n798), .A2(n797), .ZN(G282) );
  NAND2_X1 U882 ( .A1(G559), .A2(n1019), .ZN(n799) );
  XNOR2_X1 U883 ( .A(n799), .B(n1022), .ZN(n821) );
  XOR2_X1 U884 ( .A(n821), .B(KEYINPUT77), .Z(n800) );
  NOR2_X1 U885 ( .A1(G860), .A2(n800), .ZN(n801) );
  XOR2_X1 U886 ( .A(KEYINPUT80), .B(n801), .Z(n814) );
  NAND2_X1 U887 ( .A1(n802), .A2(G93), .ZN(n805) );
  NAND2_X1 U888 ( .A1(G80), .A2(n803), .ZN(n804) );
  NAND2_X1 U889 ( .A1(n805), .A2(n804), .ZN(n813) );
  NAND2_X1 U890 ( .A1(n806), .A2(G55), .ZN(n807) );
  XNOR2_X1 U891 ( .A(n807), .B(KEYINPUT78), .ZN(n810) );
  NAND2_X1 U892 ( .A1(G67), .A2(n808), .ZN(n809) );
  NAND2_X1 U893 ( .A1(n810), .A2(n809), .ZN(n811) );
  XOR2_X1 U894 ( .A(KEYINPUT79), .B(n811), .Z(n812) );
  NOR2_X1 U895 ( .A1(n813), .A2(n812), .ZN(n824) );
  XOR2_X1 U896 ( .A(n814), .B(n824), .Z(G145) );
  INV_X1 U897 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U898 ( .A(G299), .B(G288), .ZN(n820) );
  XOR2_X1 U899 ( .A(KEYINPUT85), .B(KEYINPUT19), .Z(n816) );
  XNOR2_X1 U900 ( .A(G166), .B(n824), .ZN(n815) );
  XNOR2_X1 U901 ( .A(n816), .B(n815), .ZN(n817) );
  XOR2_X1 U902 ( .A(n817), .B(G290), .Z(n818) );
  XNOR2_X1 U903 ( .A(G305), .B(n818), .ZN(n819) );
  XNOR2_X1 U904 ( .A(n820), .B(n819), .ZN(n1018) );
  XNOR2_X1 U905 ( .A(n1018), .B(n821), .ZN(n822) );
  NAND2_X1 U906 ( .A1(n822), .A2(G868), .ZN(n823) );
  XNOR2_X1 U907 ( .A(n823), .B(KEYINPUT86), .ZN(n826) );
  OR2_X1 U908 ( .A1(G868), .A2(n824), .ZN(n825) );
  NAND2_X1 U909 ( .A1(n826), .A2(n825), .ZN(G295) );
  NAND2_X1 U910 ( .A1(G2084), .A2(G2078), .ZN(n827) );
  XOR2_X1 U911 ( .A(KEYINPUT20), .B(n827), .Z(n828) );
  NAND2_X1 U912 ( .A1(G2090), .A2(n828), .ZN(n829) );
  XNOR2_X1 U913 ( .A(KEYINPUT21), .B(n829), .ZN(n830) );
  NAND2_X1 U914 ( .A1(n830), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U915 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U916 ( .A(KEYINPUT22), .B(KEYINPUT87), .Z(n832) );
  NAND2_X1 U917 ( .A1(G132), .A2(G82), .ZN(n831) );
  XNOR2_X1 U918 ( .A(n832), .B(n831), .ZN(n833) );
  NOR2_X1 U919 ( .A1(n833), .A2(G218), .ZN(n834) );
  NAND2_X1 U920 ( .A1(G96), .A2(n834), .ZN(n967) );
  NAND2_X1 U921 ( .A1(n967), .A2(G2106), .ZN(n838) );
  NAND2_X1 U922 ( .A1(G69), .A2(G120), .ZN(n835) );
  NOR2_X1 U923 ( .A1(G237), .A2(n835), .ZN(n836) );
  NAND2_X1 U924 ( .A1(G108), .A2(n836), .ZN(n968) );
  NAND2_X1 U925 ( .A1(n968), .A2(G567), .ZN(n837) );
  NAND2_X1 U926 ( .A1(n838), .A2(n837), .ZN(n969) );
  NAND2_X1 U927 ( .A1(G661), .A2(G483), .ZN(n839) );
  NOR2_X1 U928 ( .A1(n969), .A2(n839), .ZN(n845) );
  NAND2_X1 U929 ( .A1(n845), .A2(G36), .ZN(G176) );
  NAND2_X1 U930 ( .A1(G2106), .A2(n840), .ZN(G217) );
  NAND2_X1 U931 ( .A1(G15), .A2(G2), .ZN(n842) );
  INV_X1 U932 ( .A(G661), .ZN(n841) );
  NOR2_X1 U933 ( .A1(n842), .A2(n841), .ZN(n843) );
  XNOR2_X1 U934 ( .A(n843), .B(KEYINPUT111), .ZN(G259) );
  NAND2_X1 U935 ( .A1(G3), .A2(G1), .ZN(n844) );
  NAND2_X1 U936 ( .A1(n845), .A2(n844), .ZN(G188) );
  NAND2_X1 U938 ( .A1(G124), .A2(n999), .ZN(n846) );
  XNOR2_X1 U939 ( .A(n846), .B(KEYINPUT44), .ZN(n848) );
  NAND2_X1 U940 ( .A1(n998), .A2(G112), .ZN(n847) );
  NAND2_X1 U941 ( .A1(n848), .A2(n847), .ZN(n852) );
  NAND2_X1 U942 ( .A1(G136), .A2(n723), .ZN(n850) );
  NAND2_X1 U943 ( .A1(G100), .A2(n1003), .ZN(n849) );
  NAND2_X1 U944 ( .A1(n850), .A2(n849), .ZN(n851) );
  NOR2_X1 U945 ( .A1(n852), .A2(n851), .ZN(G162) );
  XNOR2_X1 U946 ( .A(G1996), .B(G32), .ZN(n855) );
  XNOR2_X1 U947 ( .A(n853), .B(G27), .ZN(n854) );
  NOR2_X1 U948 ( .A1(n855), .A2(n854), .ZN(n856) );
  XNOR2_X1 U949 ( .A(KEYINPUT122), .B(n856), .ZN(n863) );
  XOR2_X1 U950 ( .A(G2072), .B(G33), .Z(n857) );
  NAND2_X1 U951 ( .A1(n857), .A2(G28), .ZN(n861) );
  XNOR2_X1 U952 ( .A(KEYINPUT121), .B(n858), .ZN(n859) );
  XNOR2_X1 U953 ( .A(G25), .B(n859), .ZN(n860) );
  NOR2_X1 U954 ( .A1(n861), .A2(n860), .ZN(n862) );
  NAND2_X1 U955 ( .A1(n863), .A2(n862), .ZN(n865) );
  XNOR2_X1 U956 ( .A(G26), .B(G2067), .ZN(n864) );
  NOR2_X1 U957 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U958 ( .A(KEYINPUT53), .B(n866), .Z(n870) );
  XNOR2_X1 U959 ( .A(KEYINPUT54), .B(KEYINPUT123), .ZN(n867) );
  XNOR2_X1 U960 ( .A(n867), .B(G34), .ZN(n868) );
  XNOR2_X1 U961 ( .A(G2084), .B(n868), .ZN(n869) );
  NAND2_X1 U962 ( .A1(n870), .A2(n869), .ZN(n872) );
  XNOR2_X1 U963 ( .A(G35), .B(G2090), .ZN(n871) );
  NOR2_X1 U964 ( .A1(n872), .A2(n871), .ZN(n961) );
  NAND2_X1 U965 ( .A1(KEYINPUT55), .A2(n961), .ZN(n873) );
  NAND2_X1 U966 ( .A1(G11), .A2(n873), .ZN(n960) );
  XNOR2_X1 U967 ( .A(G164), .B(G2078), .ZN(n883) );
  NAND2_X1 U968 ( .A1(G139), .A2(n723), .ZN(n875) );
  NAND2_X1 U969 ( .A1(G103), .A2(n1003), .ZN(n874) );
  NAND2_X1 U970 ( .A1(n875), .A2(n874), .ZN(n880) );
  NAND2_X1 U971 ( .A1(G115), .A2(n998), .ZN(n877) );
  NAND2_X1 U972 ( .A1(G127), .A2(n999), .ZN(n876) );
  NAND2_X1 U973 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U974 ( .A(KEYINPUT47), .B(n878), .Z(n879) );
  NOR2_X1 U975 ( .A1(n880), .A2(n879), .ZN(n1011) );
  XNOR2_X1 U976 ( .A(G2072), .B(n1011), .ZN(n881) );
  XNOR2_X1 U977 ( .A(n881), .B(KEYINPUT120), .ZN(n882) );
  NAND2_X1 U978 ( .A1(n883), .A2(n882), .ZN(n884) );
  XNOR2_X1 U979 ( .A(n884), .B(KEYINPUT50), .ZN(n903) );
  XNOR2_X1 U980 ( .A(G160), .B(G2084), .ZN(n885) );
  NAND2_X1 U981 ( .A1(n885), .A2(n1013), .ZN(n886) );
  NOR2_X1 U982 ( .A1(n887), .A2(n886), .ZN(n888) );
  XNOR2_X1 U983 ( .A(n888), .B(KEYINPUT117), .ZN(n889) );
  NOR2_X1 U984 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U985 ( .A(KEYINPUT118), .B(n891), .Z(n896) );
  XOR2_X1 U986 ( .A(G2090), .B(G162), .Z(n892) );
  NOR2_X1 U987 ( .A1(n893), .A2(n892), .ZN(n894) );
  XNOR2_X1 U988 ( .A(KEYINPUT51), .B(n894), .ZN(n895) );
  NOR2_X1 U989 ( .A1(n896), .A2(n895), .ZN(n897) );
  NAND2_X1 U990 ( .A1(n898), .A2(n897), .ZN(n899) );
  XNOR2_X1 U991 ( .A(n899), .B(KEYINPUT119), .ZN(n901) );
  NAND2_X1 U992 ( .A1(n901), .A2(n900), .ZN(n902) );
  NOR2_X1 U993 ( .A1(n903), .A2(n902), .ZN(n904) );
  XNOR2_X1 U994 ( .A(KEYINPUT52), .B(n904), .ZN(n906) );
  INV_X1 U995 ( .A(KEYINPUT55), .ZN(n905) );
  NAND2_X1 U996 ( .A1(n906), .A2(n905), .ZN(n907) );
  NAND2_X1 U997 ( .A1(n907), .A2(G29), .ZN(n958) );
  XOR2_X1 U998 ( .A(G16), .B(KEYINPUT56), .Z(n930) );
  XNOR2_X1 U999 ( .A(G1341), .B(n1022), .ZN(n908) );
  NOR2_X1 U1000 ( .A1(n909), .A2(n908), .ZN(n919) );
  XNOR2_X1 U1001 ( .A(n911), .B(n910), .ZN(n913) );
  XNOR2_X1 U1002 ( .A(G303), .B(G1971), .ZN(n912) );
  NOR2_X1 U1003 ( .A1(n913), .A2(n912), .ZN(n915) );
  NAND2_X1 U1004 ( .A1(n915), .A2(n914), .ZN(n916) );
  NOR2_X1 U1005 ( .A1(n917), .A2(n916), .ZN(n918) );
  NAND2_X1 U1006 ( .A1(n919), .A2(n918), .ZN(n928) );
  XOR2_X1 U1007 ( .A(n1019), .B(G1348), .Z(n921) );
  XOR2_X1 U1008 ( .A(G171), .B(G1961), .Z(n920) );
  NOR2_X1 U1009 ( .A1(n921), .A2(n920), .ZN(n926) );
  XOR2_X1 U1010 ( .A(G168), .B(G1966), .Z(n922) );
  NOR2_X1 U1011 ( .A1(n923), .A2(n922), .ZN(n924) );
  XOR2_X1 U1012 ( .A(KEYINPUT57), .B(n924), .Z(n925) );
  NAND2_X1 U1013 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1014 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1015 ( .A1(n930), .A2(n929), .ZN(n955) );
  XNOR2_X1 U1016 ( .A(G1348), .B(KEYINPUT59), .ZN(n931) );
  XNOR2_X1 U1017 ( .A(n931), .B(G4), .ZN(n935) );
  XNOR2_X1 U1018 ( .A(G1956), .B(G20), .ZN(n933) );
  XNOR2_X1 U1019 ( .A(G1981), .B(G6), .ZN(n932) );
  NOR2_X1 U1020 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1021 ( .A1(n935), .A2(n934), .ZN(n938) );
  XOR2_X1 U1022 ( .A(KEYINPUT125), .B(G1341), .Z(n936) );
  XNOR2_X1 U1023 ( .A(G19), .B(n936), .ZN(n937) );
  NOR2_X1 U1024 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1025 ( .A(KEYINPUT60), .B(n939), .ZN(n949) );
  XNOR2_X1 U1026 ( .A(G1961), .B(KEYINPUT124), .ZN(n940) );
  XNOR2_X1 U1027 ( .A(n940), .B(G5), .ZN(n947) );
  XNOR2_X1 U1028 ( .A(G1971), .B(G22), .ZN(n942) );
  XNOR2_X1 U1029 ( .A(G23), .B(G1976), .ZN(n941) );
  NOR2_X1 U1030 ( .A1(n942), .A2(n941), .ZN(n944) );
  XOR2_X1 U1031 ( .A(G1986), .B(G24), .Z(n943) );
  NAND2_X1 U1032 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1033 ( .A(KEYINPUT58), .B(n945), .ZN(n946) );
  NOR2_X1 U1034 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1035 ( .A1(n949), .A2(n948), .ZN(n951) );
  XNOR2_X1 U1036 ( .A(G21), .B(G1966), .ZN(n950) );
  NOR2_X1 U1037 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1038 ( .A(KEYINPUT61), .B(n952), .Z(n953) );
  NOR2_X1 U1039 ( .A1(G16), .A2(n953), .ZN(n954) );
  NOR2_X1 U1040 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1041 ( .A(n956), .B(KEYINPUT126), .ZN(n957) );
  NAND2_X1 U1042 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1043 ( .A1(n960), .A2(n959), .ZN(n965) );
  INV_X1 U1044 ( .A(n961), .ZN(n963) );
  NOR2_X1 U1045 ( .A1(G29), .A2(KEYINPUT55), .ZN(n962) );
  NAND2_X1 U1046 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1047 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1048 ( .A(KEYINPUT62), .B(n966), .Z(G311) );
  XNOR2_X1 U1049 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1050 ( .A(G132), .ZN(G219) );
  INV_X1 U1051 ( .A(G120), .ZN(G236) );
  INV_X1 U1052 ( .A(G96), .ZN(G221) );
  INV_X1 U1053 ( .A(G82), .ZN(G220) );
  INV_X1 U1054 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1055 ( .A1(n968), .A2(n967), .ZN(G325) );
  INV_X1 U1056 ( .A(G325), .ZN(G261) );
  INV_X1 U1057 ( .A(n969), .ZN(G319) );
  XNOR2_X1 U1058 ( .A(G1986), .B(G1981), .ZN(n979) );
  XOR2_X1 U1059 ( .A(G1971), .B(G1956), .Z(n971) );
  XNOR2_X1 U1060 ( .A(G1996), .B(G1966), .ZN(n970) );
  XNOR2_X1 U1061 ( .A(n971), .B(n970), .ZN(n975) );
  XOR2_X1 U1062 ( .A(KEYINPUT114), .B(G2474), .Z(n973) );
  XNOR2_X1 U1063 ( .A(G1991), .B(G1961), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(n973), .B(n972), .ZN(n974) );
  XOR2_X1 U1065 ( .A(n975), .B(n974), .Z(n977) );
  XNOR2_X1 U1066 ( .A(G1976), .B(KEYINPUT41), .ZN(n976) );
  XNOR2_X1 U1067 ( .A(n977), .B(n976), .ZN(n978) );
  XNOR2_X1 U1068 ( .A(n979), .B(n978), .ZN(G229) );
  XOR2_X1 U1069 ( .A(KEYINPUT43), .B(G2678), .Z(n981) );
  XNOR2_X1 U1070 ( .A(G2072), .B(G2090), .ZN(n980) );
  XNOR2_X1 U1071 ( .A(n981), .B(n980), .ZN(n985) );
  XOR2_X1 U1072 ( .A(KEYINPUT113), .B(KEYINPUT112), .Z(n983) );
  XNOR2_X1 U1073 ( .A(G2067), .B(KEYINPUT42), .ZN(n982) );
  XNOR2_X1 U1074 ( .A(n983), .B(n982), .ZN(n984) );
  XOR2_X1 U1075 ( .A(n985), .B(n984), .Z(n987) );
  XNOR2_X1 U1076 ( .A(G2096), .B(G2100), .ZN(n986) );
  XNOR2_X1 U1077 ( .A(n987), .B(n986), .ZN(n989) );
  XOR2_X1 U1078 ( .A(G2084), .B(G2078), .Z(n988) );
  XNOR2_X1 U1079 ( .A(n989), .B(n988), .ZN(G227) );
  XOR2_X1 U1080 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n991) );
  XNOR2_X1 U1081 ( .A(G160), .B(KEYINPUT116), .ZN(n990) );
  XNOR2_X1 U1082 ( .A(n991), .B(n990), .ZN(n992) );
  XNOR2_X1 U1083 ( .A(n993), .B(n992), .ZN(n997) );
  XOR2_X1 U1084 ( .A(n995), .B(n994), .Z(n996) );
  XNOR2_X1 U1085 ( .A(n997), .B(n996), .ZN(n1010) );
  NAND2_X1 U1086 ( .A1(G118), .A2(n998), .ZN(n1001) );
  NAND2_X1 U1087 ( .A1(G130), .A2(n999), .ZN(n1000) );
  NAND2_X1 U1088 ( .A1(n1001), .A2(n1000), .ZN(n1008) );
  NAND2_X1 U1089 ( .A1(n723), .A2(G142), .ZN(n1002) );
  XOR2_X1 U1090 ( .A(KEYINPUT115), .B(n1002), .Z(n1005) );
  NAND2_X1 U1091 ( .A1(n1003), .A2(G106), .ZN(n1004) );
  NAND2_X1 U1092 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1093 ( .A(n1006), .B(KEYINPUT45), .Z(n1007) );
  NOR2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1095 ( .A(n1010), .B(n1009), .Z(n1016) );
  XOR2_X1 U1096 ( .A(n1011), .B(G162), .Z(n1012) );
  XNOR2_X1 U1097 ( .A(n1013), .B(n1012), .ZN(n1014) );
  XNOR2_X1 U1098 ( .A(G164), .B(n1014), .ZN(n1015) );
  XNOR2_X1 U1099 ( .A(n1016), .B(n1015), .ZN(n1017) );
  NOR2_X1 U1100 ( .A1(G37), .A2(n1017), .ZN(G395) );
  XNOR2_X1 U1101 ( .A(G286), .B(n1018), .ZN(n1021) );
  XNOR2_X1 U1102 ( .A(G171), .B(n1019), .ZN(n1020) );
  XNOR2_X1 U1103 ( .A(n1021), .B(n1020), .ZN(n1023) );
  XOR2_X1 U1104 ( .A(n1023), .B(n1022), .Z(n1024) );
  NOR2_X1 U1105 ( .A1(G37), .A2(n1024), .ZN(G397) );
  XNOR2_X1 U1106 ( .A(G1341), .B(G2443), .ZN(n1034) );
  XOR2_X1 U1107 ( .A(G2451), .B(G2446), .Z(n1026) );
  XNOR2_X1 U1108 ( .A(G1348), .B(G2454), .ZN(n1025) );
  XNOR2_X1 U1109 ( .A(n1026), .B(n1025), .ZN(n1030) );
  XOR2_X1 U1110 ( .A(G2435), .B(KEYINPUT109), .Z(n1028) );
  XNOR2_X1 U1111 ( .A(G2438), .B(KEYINPUT110), .ZN(n1027) );
  XNOR2_X1 U1112 ( .A(n1028), .B(n1027), .ZN(n1029) );
  XOR2_X1 U1113 ( .A(n1030), .B(n1029), .Z(n1032) );
  XNOR2_X1 U1114 ( .A(G2430), .B(G2427), .ZN(n1031) );
  XNOR2_X1 U1115 ( .A(n1032), .B(n1031), .ZN(n1033) );
  XNOR2_X1 U1116 ( .A(n1034), .B(n1033), .ZN(n1035) );
  NAND2_X1 U1117 ( .A1(n1035), .A2(G14), .ZN(n1041) );
  NAND2_X1 U1118 ( .A1(G319), .A2(n1041), .ZN(n1038) );
  NOR2_X1 U1119 ( .A1(G229), .A2(G227), .ZN(n1036) );
  XNOR2_X1 U1120 ( .A(KEYINPUT49), .B(n1036), .ZN(n1037) );
  NOR2_X1 U1121 ( .A1(n1038), .A2(n1037), .ZN(n1040) );
  NOR2_X1 U1122 ( .A1(G395), .A2(G397), .ZN(n1039) );
  NAND2_X1 U1123 ( .A1(n1040), .A2(n1039), .ZN(G225) );
  INV_X1 U1124 ( .A(G225), .ZN(G308) );
  INV_X1 U1125 ( .A(G108), .ZN(G238) );
  INV_X1 U1126 ( .A(n1041), .ZN(G401) );
endmodule

