

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596;

  XNOR2_X1 U322 ( .A(n381), .B(n380), .ZN(n383) );
  XNOR2_X1 U323 ( .A(n379), .B(KEYINPUT19), .ZN(n380) );
  INV_X1 U324 ( .A(KEYINPUT17), .ZN(n379) );
  XNOR2_X1 U325 ( .A(n320), .B(n319), .ZN(n325) );
  XNOR2_X1 U326 ( .A(n585), .B(KEYINPUT41), .ZN(n568) );
  XNOR2_X1 U327 ( .A(n480), .B(n479), .ZN(n511) );
  XOR2_X1 U328 ( .A(n455), .B(n454), .Z(n539) );
  AND2_X1 U329 ( .A1(G227GAT), .A2(G233GAT), .ZN(n290) );
  XOR2_X1 U330 ( .A(n355), .B(n333), .Z(n291) );
  XNOR2_X1 U331 ( .A(n385), .B(G183GAT), .ZN(n386) );
  XNOR2_X1 U332 ( .A(KEYINPUT110), .B(KEYINPUT47), .ZN(n371) );
  XNOR2_X1 U333 ( .A(n455), .B(n386), .ZN(n387) );
  XNOR2_X1 U334 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U335 ( .A(n372), .B(n371), .ZN(n377) );
  XNOR2_X1 U336 ( .A(n439), .B(n290), .ZN(n441) );
  XNOR2_X1 U337 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U338 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U339 ( .A(n441), .B(n440), .ZN(n442) );
  NOR2_X1 U340 ( .A1(n594), .A2(n477), .ZN(n478) );
  XNOR2_X1 U341 ( .A(n451), .B(n450), .ZN(n452) );
  NOR2_X1 U342 ( .A1(n421), .A2(n481), .ZN(n580) );
  XNOR2_X1 U343 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U344 ( .A(n350), .B(n349), .ZN(n585) );
  XOR2_X1 U345 ( .A(n330), .B(n329), .Z(n589) );
  INV_X1 U346 ( .A(G43GAT), .ZN(n487) );
  XNOR2_X1 U347 ( .A(n396), .B(n395), .ZN(n508) );
  XNOR2_X1 U348 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U349 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U350 ( .A(n494), .B(n493), .ZN(G1351GAT) );
  XNOR2_X1 U351 ( .A(n490), .B(n489), .ZN(G1330GAT) );
  XOR2_X1 U352 ( .A(G29GAT), .B(KEYINPUT8), .Z(n293) );
  XNOR2_X1 U353 ( .A(KEYINPUT7), .B(KEYINPUT73), .ZN(n292) );
  XNOR2_X1 U354 ( .A(n293), .B(n292), .ZN(n358) );
  XOR2_X1 U355 ( .A(n358), .B(KEYINPUT67), .Z(n295) );
  NAND2_X1 U356 ( .A1(G229GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U357 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U358 ( .A(KEYINPUT70), .B(KEYINPUT69), .Z(n297) );
  XNOR2_X1 U359 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n296) );
  XNOR2_X1 U360 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U361 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U362 ( .A(KEYINPUT71), .B(G1GAT), .Z(n301) );
  XNOR2_X1 U363 ( .A(G169GAT), .B(G8GAT), .ZN(n300) );
  XNOR2_X1 U364 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U365 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U366 ( .A(G22GAT), .B(G43GAT), .Z(n305) );
  XNOR2_X1 U367 ( .A(G50GAT), .B(G36GAT), .ZN(n304) );
  XNOR2_X1 U368 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U369 ( .A(n307), .B(n306), .Z(n315) );
  XOR2_X1 U370 ( .A(KEYINPUT68), .B(KEYINPUT74), .Z(n309) );
  XNOR2_X1 U371 ( .A(KEYINPUT72), .B(KEYINPUT66), .ZN(n308) );
  XNOR2_X1 U372 ( .A(n309), .B(n308), .ZN(n313) );
  XOR2_X1 U373 ( .A(G15GAT), .B(G113GAT), .Z(n311) );
  XNOR2_X1 U374 ( .A(G197GAT), .B(G141GAT), .ZN(n310) );
  XNOR2_X1 U375 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U376 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U377 ( .A(n315), .B(n314), .Z(n540) );
  INV_X1 U378 ( .A(n540), .ZN(n581) );
  XOR2_X1 U379 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n317) );
  XNOR2_X1 U380 ( .A(KEYINPUT81), .B(KEYINPUT82), .ZN(n316) );
  XNOR2_X1 U381 ( .A(n317), .B(n316), .ZN(n330) );
  XNOR2_X1 U382 ( .A(G15GAT), .B(G183GAT), .ZN(n318) );
  XNOR2_X1 U383 ( .A(n318), .B(G127GAT), .ZN(n440) );
  XNOR2_X1 U384 ( .A(G1GAT), .B(n440), .ZN(n320) );
  INV_X1 U385 ( .A(KEYINPUT15), .ZN(n319) );
  XNOR2_X1 U386 ( .A(G71GAT), .B(G57GAT), .ZN(n321) );
  XNOR2_X1 U387 ( .A(n321), .B(KEYINPUT13), .ZN(n333) );
  XOR2_X1 U388 ( .A(G22GAT), .B(G155GAT), .Z(n422) );
  XNOR2_X1 U389 ( .A(n333), .B(n422), .ZN(n323) );
  AND2_X1 U390 ( .A1(G231GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U391 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U392 ( .A(G8GAT), .B(G211GAT), .Z(n384) );
  XOR2_X1 U393 ( .A(n326), .B(n384), .Z(n328) );
  XNOR2_X1 U394 ( .A(G78GAT), .B(G64GAT), .ZN(n327) );
  XNOR2_X1 U395 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U396 ( .A(n589), .B(KEYINPUT109), .ZN(n575) );
  XOR2_X1 U397 ( .A(KEYINPUT33), .B(KEYINPUT76), .Z(n332) );
  XNOR2_X1 U398 ( .A(KEYINPUT31), .B(KEYINPUT32), .ZN(n331) );
  XNOR2_X1 U399 ( .A(n332), .B(n331), .ZN(n350) );
  XOR2_X1 U400 ( .A(G99GAT), .B(G85GAT), .Z(n355) );
  NAND2_X1 U401 ( .A1(G230GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U402 ( .A(n291), .B(n334), .ZN(n336) );
  INV_X1 U403 ( .A(KEYINPUT77), .ZN(n335) );
  XNOR2_X1 U404 ( .A(n336), .B(n335), .ZN(n342) );
  XOR2_X1 U405 ( .A(G78GAT), .B(G148GAT), .Z(n338) );
  XNOR2_X1 U406 ( .A(G106GAT), .B(G204GAT), .ZN(n337) );
  XNOR2_X1 U407 ( .A(n338), .B(n337), .ZN(n435) );
  XNOR2_X1 U408 ( .A(n435), .B(KEYINPUT75), .ZN(n340) );
  XOR2_X1 U409 ( .A(G92GAT), .B(G64GAT), .Z(n395) );
  INV_X1 U410 ( .A(n395), .ZN(n339) );
  XNOR2_X1 U411 ( .A(G176GAT), .B(G120GAT), .ZN(n344) );
  NAND2_X1 U412 ( .A1(n343), .A2(n344), .ZN(n348) );
  INV_X1 U413 ( .A(n343), .ZN(n346) );
  INV_X1 U414 ( .A(n344), .ZN(n345) );
  NAND2_X1 U415 ( .A1(n346), .A2(n345), .ZN(n347) );
  AND2_X1 U416 ( .A1(n348), .A2(n347), .ZN(n349) );
  NOR2_X1 U417 ( .A1(n581), .A2(n568), .ZN(n351) );
  XNOR2_X1 U418 ( .A(n351), .B(KEYINPUT46), .ZN(n352) );
  NOR2_X1 U419 ( .A1(n575), .A2(n352), .ZN(n370) );
  XOR2_X1 U420 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n354) );
  XNOR2_X1 U421 ( .A(KEYINPUT78), .B(KEYINPUT80), .ZN(n353) );
  XNOR2_X1 U422 ( .A(n354), .B(n353), .ZN(n369) );
  XOR2_X1 U423 ( .A(KEYINPUT79), .B(KEYINPUT65), .Z(n357) );
  XOR2_X1 U424 ( .A(G36GAT), .B(G218GAT), .Z(n388) );
  XNOR2_X1 U425 ( .A(n388), .B(n355), .ZN(n356) );
  XNOR2_X1 U426 ( .A(n357), .B(n356), .ZN(n362) );
  XOR2_X1 U427 ( .A(G50GAT), .B(G162GAT), .Z(n426) );
  XOR2_X1 U428 ( .A(n426), .B(n358), .Z(n360) );
  NAND2_X1 U429 ( .A1(G232GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U430 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U431 ( .A(n362), .B(n361), .Z(n367) );
  XOR2_X1 U432 ( .A(G43GAT), .B(G134GAT), .Z(n439) );
  XOR2_X1 U433 ( .A(KEYINPUT11), .B(G92GAT), .Z(n364) );
  XNOR2_X1 U434 ( .A(G190GAT), .B(G106GAT), .ZN(n363) );
  XNOR2_X1 U435 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U436 ( .A(n439), .B(n365), .ZN(n366) );
  XNOR2_X1 U437 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U438 ( .A(n369), .B(n368), .Z(n550) );
  INV_X1 U439 ( .A(n550), .ZN(n565) );
  NAND2_X1 U440 ( .A1(n370), .A2(n565), .ZN(n372) );
  XOR2_X1 U441 ( .A(KEYINPUT36), .B(n550), .Z(n594) );
  NOR2_X1 U442 ( .A1(n594), .A2(n589), .ZN(n373) );
  XNOR2_X1 U443 ( .A(KEYINPUT45), .B(n373), .ZN(n374) );
  NAND2_X1 U444 ( .A1(n374), .A2(n581), .ZN(n375) );
  NOR2_X1 U445 ( .A1(n375), .A2(n585), .ZN(n376) );
  NOR2_X1 U446 ( .A1(n377), .A2(n376), .ZN(n378) );
  XNOR2_X1 U447 ( .A(n378), .B(KEYINPUT48), .ZN(n536) );
  INV_X1 U448 ( .A(n536), .ZN(n397) );
  XOR2_X1 U449 ( .A(G197GAT), .B(KEYINPUT21), .Z(n423) );
  INV_X1 U450 ( .A(n423), .ZN(n391) );
  XNOR2_X1 U451 ( .A(G176GAT), .B(KEYINPUT18), .ZN(n381) );
  XNOR2_X1 U452 ( .A(G169GAT), .B(G190GAT), .ZN(n382) );
  XNOR2_X1 U453 ( .A(n383), .B(n382), .ZN(n455) );
  XOR2_X1 U454 ( .A(n384), .B(G204GAT), .Z(n385) );
  XNOR2_X1 U455 ( .A(n388), .B(n387), .ZN(n390) );
  AND2_X1 U456 ( .A1(G226GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U457 ( .A(n390), .B(n389), .ZN(n392) );
  OR2_X1 U458 ( .A1(n391), .A2(n392), .ZN(n394) );
  NAND2_X1 U459 ( .A1(n391), .A2(n392), .ZN(n393) );
  NAND2_X1 U460 ( .A1(n394), .A2(n393), .ZN(n396) );
  NAND2_X1 U461 ( .A1(n397), .A2(n508), .ZN(n399) );
  XOR2_X1 U462 ( .A(KEYINPUT119), .B(KEYINPUT54), .Z(n398) );
  XNOR2_X1 U463 ( .A(n399), .B(n398), .ZN(n421) );
  XOR2_X1 U464 ( .A(G57GAT), .B(G155GAT), .Z(n401) );
  XNOR2_X1 U465 ( .A(G127GAT), .B(G148GAT), .ZN(n400) );
  XNOR2_X1 U466 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U467 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n403) );
  XNOR2_X1 U468 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n402) );
  XNOR2_X1 U469 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U470 ( .A(n405), .B(n404), .Z(n410) );
  XOR2_X1 U471 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n407) );
  NAND2_X1 U472 ( .A1(G225GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U473 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U474 ( .A(KEYINPUT1), .B(n408), .ZN(n409) );
  XNOR2_X1 U475 ( .A(n410), .B(n409), .ZN(n414) );
  XOR2_X1 U476 ( .A(G85GAT), .B(G162GAT), .Z(n412) );
  XNOR2_X1 U477 ( .A(G29GAT), .B(G134GAT), .ZN(n411) );
  XNOR2_X1 U478 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U479 ( .A(n414), .B(n413), .Z(n420) );
  XNOR2_X1 U480 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n415) );
  XNOR2_X1 U481 ( .A(n415), .B(G120GAT), .ZN(n443) );
  XOR2_X1 U482 ( .A(KEYINPUT2), .B(KEYINPUT90), .Z(n417) );
  XNOR2_X1 U483 ( .A(KEYINPUT91), .B(KEYINPUT3), .ZN(n416) );
  XNOR2_X1 U484 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U485 ( .A(G141GAT), .B(n418), .Z(n431) );
  XNOR2_X1 U486 ( .A(n443), .B(n431), .ZN(n419) );
  XOR2_X1 U487 ( .A(n420), .B(n419), .Z(n526) );
  INV_X1 U488 ( .A(n526), .ZN(n481) );
  XOR2_X1 U489 ( .A(n423), .B(n422), .Z(n425) );
  NAND2_X1 U490 ( .A1(G228GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U491 ( .A(n425), .B(n424), .ZN(n427) );
  XOR2_X1 U492 ( .A(n427), .B(n426), .Z(n433) );
  XOR2_X1 U493 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n429) );
  XNOR2_X1 U494 ( .A(G218GAT), .B(KEYINPUT92), .ZN(n428) );
  XNOR2_X1 U495 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U496 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U497 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U498 ( .A(n434), .B(KEYINPUT22), .Z(n437) );
  XNOR2_X1 U499 ( .A(n435), .B(G211GAT), .ZN(n436) );
  XNOR2_X1 U500 ( .A(n437), .B(n436), .ZN(n471) );
  NAND2_X1 U501 ( .A1(n580), .A2(n471), .ZN(n438) );
  XNOR2_X1 U502 ( .A(n438), .B(KEYINPUT55), .ZN(n456) );
  XOR2_X1 U503 ( .A(n442), .B(KEYINPUT83), .Z(n453) );
  XNOR2_X1 U504 ( .A(n443), .B(G71GAT), .ZN(n451) );
  XOR2_X1 U505 ( .A(KEYINPUT88), .B(KEYINPUT86), .Z(n445) );
  XNOR2_X1 U506 ( .A(KEYINPUT20), .B(KEYINPUT85), .ZN(n444) );
  XNOR2_X1 U507 ( .A(n445), .B(n444), .ZN(n449) );
  XOR2_X1 U508 ( .A(KEYINPUT87), .B(KEYINPUT84), .Z(n447) );
  XNOR2_X1 U509 ( .A(G99GAT), .B(KEYINPUT64), .ZN(n446) );
  XNOR2_X1 U510 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U511 ( .A(n449), .B(n448), .ZN(n450) );
  INV_X1 U512 ( .A(n539), .ZN(n486) );
  NAND2_X1 U513 ( .A1(n456), .A2(n486), .ZN(n574) );
  NOR2_X1 U514 ( .A1(n581), .A2(n574), .ZN(n459) );
  INV_X1 U515 ( .A(G169GAT), .ZN(n457) );
  XNOR2_X1 U516 ( .A(n457), .B(KEYINPUT120), .ZN(n458) );
  XNOR2_X1 U517 ( .A(n459), .B(n458), .ZN(G1348GAT) );
  NOR2_X1 U518 ( .A1(n471), .A2(n486), .ZN(n461) );
  XNOR2_X1 U519 ( .A(KEYINPUT95), .B(KEYINPUT26), .ZN(n460) );
  XOR2_X1 U520 ( .A(n461), .B(n460), .Z(n579) );
  XNOR2_X1 U521 ( .A(KEYINPUT27), .B(n508), .ZN(n469) );
  AND2_X1 U522 ( .A1(n579), .A2(n469), .ZN(n462) );
  XOR2_X1 U523 ( .A(KEYINPUT96), .B(n462), .Z(n467) );
  NAND2_X1 U524 ( .A1(n486), .A2(n508), .ZN(n463) );
  XOR2_X1 U525 ( .A(KEYINPUT97), .B(n463), .Z(n464) );
  NAND2_X1 U526 ( .A1(n464), .A2(n471), .ZN(n465) );
  XOR2_X1 U527 ( .A(KEYINPUT25), .B(n465), .Z(n466) );
  NAND2_X1 U528 ( .A1(n467), .A2(n466), .ZN(n468) );
  NAND2_X1 U529 ( .A1(n468), .A2(n526), .ZN(n474) );
  NAND2_X1 U530 ( .A1(n481), .A2(n469), .ZN(n535) );
  XNOR2_X1 U531 ( .A(KEYINPUT89), .B(n539), .ZN(n470) );
  NOR2_X1 U532 ( .A1(n535), .A2(n470), .ZN(n472) );
  XOR2_X1 U533 ( .A(n471), .B(KEYINPUT28), .Z(n510) );
  INV_X1 U534 ( .A(n510), .ZN(n537) );
  NAND2_X1 U535 ( .A1(n472), .A2(n537), .ZN(n473) );
  NAND2_X1 U536 ( .A1(n474), .A2(n473), .ZN(n496) );
  NAND2_X1 U537 ( .A1(n496), .A2(n589), .ZN(n476) );
  INV_X1 U538 ( .A(KEYINPUT101), .ZN(n475) );
  XNOR2_X1 U539 ( .A(n476), .B(n475), .ZN(n477) );
  XOR2_X1 U540 ( .A(KEYINPUT37), .B(n478), .Z(n525) );
  NOR2_X1 U541 ( .A1(n581), .A2(n585), .ZN(n499) );
  NAND2_X1 U542 ( .A1(n525), .A2(n499), .ZN(n480) );
  XOR2_X1 U543 ( .A(KEYINPUT102), .B(KEYINPUT38), .Z(n479) );
  NAND2_X1 U544 ( .A1(n511), .A2(n481), .ZN(n485) );
  XOR2_X1 U545 ( .A(G29GAT), .B(KEYINPUT100), .Z(n483) );
  XOR2_X1 U546 ( .A(KEYINPUT39), .B(KEYINPUT103), .Z(n482) );
  XNOR2_X1 U547 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U548 ( .A(n485), .B(n484), .ZN(G1328GAT) );
  NAND2_X1 U549 ( .A1(n511), .A2(n486), .ZN(n490) );
  XOR2_X1 U550 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n488) );
  NOR2_X1 U551 ( .A1(n565), .A2(n574), .ZN(n494) );
  XNOR2_X1 U552 ( .A(KEYINPUT124), .B(KEYINPUT58), .ZN(n492) );
  INV_X1 U553 ( .A(G190GAT), .ZN(n491) );
  NOR2_X1 U554 ( .A1(n550), .A2(n589), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n495), .B(KEYINPUT16), .ZN(n497) );
  NAND2_X1 U556 ( .A1(n497), .A2(n496), .ZN(n498) );
  XOR2_X1 U557 ( .A(KEYINPUT98), .B(n498), .Z(n514) );
  NAND2_X1 U558 ( .A1(n499), .A2(n514), .ZN(n506) );
  NOR2_X1 U559 ( .A1(n526), .A2(n506), .ZN(n500) );
  XOR2_X1 U560 ( .A(G1GAT), .B(n500), .Z(n501) );
  XNOR2_X1 U561 ( .A(KEYINPUT34), .B(n501), .ZN(G1324GAT) );
  INV_X1 U562 ( .A(n508), .ZN(n529) );
  NOR2_X1 U563 ( .A1(n529), .A2(n506), .ZN(n503) );
  XNOR2_X1 U564 ( .A(G8GAT), .B(KEYINPUT99), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n503), .B(n502), .ZN(G1325GAT) );
  NOR2_X1 U566 ( .A1(n539), .A2(n506), .ZN(n505) );
  XNOR2_X1 U567 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n505), .B(n504), .ZN(G1326GAT) );
  NOR2_X1 U569 ( .A1(n537), .A2(n506), .ZN(n507) );
  XOR2_X1 U570 ( .A(G22GAT), .B(n507), .Z(G1327GAT) );
  NAND2_X1 U571 ( .A1(n508), .A2(n511), .ZN(n509) );
  XNOR2_X1 U572 ( .A(n509), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U573 ( .A(G50GAT), .B(KEYINPUT105), .Z(n513) );
  NAND2_X1 U574 ( .A1(n511), .A2(n510), .ZN(n512) );
  XNOR2_X1 U575 ( .A(n513), .B(n512), .ZN(G1331GAT) );
  NOR2_X1 U576 ( .A1(n540), .A2(n568), .ZN(n524) );
  NAND2_X1 U577 ( .A1(n524), .A2(n514), .ZN(n521) );
  NOR2_X1 U578 ( .A1(n526), .A2(n521), .ZN(n516) );
  XNOR2_X1 U579 ( .A(KEYINPUT42), .B(KEYINPUT106), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U581 ( .A(G57GAT), .B(n517), .Z(G1332GAT) );
  NOR2_X1 U582 ( .A1(n529), .A2(n521), .ZN(n519) );
  XNOR2_X1 U583 ( .A(G64GAT), .B(KEYINPUT107), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n519), .B(n518), .ZN(G1333GAT) );
  NOR2_X1 U585 ( .A1(n539), .A2(n521), .ZN(n520) );
  XOR2_X1 U586 ( .A(G71GAT), .B(n520), .Z(G1334GAT) );
  NOR2_X1 U587 ( .A1(n537), .A2(n521), .ZN(n523) );
  XNOR2_X1 U588 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(G1335GAT) );
  NAND2_X1 U590 ( .A1(n525), .A2(n524), .ZN(n532) );
  NOR2_X1 U591 ( .A1(n526), .A2(n532), .ZN(n527) );
  XOR2_X1 U592 ( .A(G85GAT), .B(n527), .Z(n528) );
  XNOR2_X1 U593 ( .A(KEYINPUT108), .B(n528), .ZN(G1336GAT) );
  NOR2_X1 U594 ( .A1(n529), .A2(n532), .ZN(n530) );
  XOR2_X1 U595 ( .A(G92GAT), .B(n530), .Z(G1337GAT) );
  NOR2_X1 U596 ( .A1(n539), .A2(n532), .ZN(n531) );
  XOR2_X1 U597 ( .A(G99GAT), .B(n531), .Z(G1338GAT) );
  NOR2_X1 U598 ( .A1(n537), .A2(n532), .ZN(n533) );
  XOR2_X1 U599 ( .A(KEYINPUT44), .B(n533), .Z(n534) );
  XNOR2_X1 U600 ( .A(G106GAT), .B(n534), .ZN(G1339GAT) );
  XOR2_X1 U601 ( .A(G113GAT), .B(KEYINPUT111), .Z(n542) );
  NOR2_X1 U602 ( .A1(n536), .A2(n535), .ZN(n556) );
  NAND2_X1 U603 ( .A1(n556), .A2(n537), .ZN(n538) );
  NOR2_X1 U604 ( .A1(n539), .A2(n538), .ZN(n551) );
  NAND2_X1 U605 ( .A1(n551), .A2(n540), .ZN(n541) );
  XNOR2_X1 U606 ( .A(n542), .B(n541), .ZN(G1340GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT112), .B(KEYINPUT49), .Z(n545) );
  INV_X1 U608 ( .A(n568), .ZN(n543) );
  NAND2_X1 U609 ( .A1(n551), .A2(n543), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U611 ( .A(G120GAT), .B(n546), .ZN(G1341GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT50), .B(KEYINPUT113), .Z(n548) );
  NAND2_X1 U613 ( .A1(n551), .A2(n575), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U615 ( .A(G127GAT), .B(n549), .ZN(G1342GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n553) );
  NAND2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(n555) );
  XOR2_X1 U619 ( .A(G134GAT), .B(KEYINPUT115), .Z(n554) );
  XNOR2_X1 U620 ( .A(n555), .B(n554), .ZN(G1343GAT) );
  NAND2_X1 U621 ( .A1(n556), .A2(n579), .ZN(n564) );
  NOR2_X1 U622 ( .A1(n581), .A2(n564), .ZN(n557) );
  XOR2_X1 U623 ( .A(G141GAT), .B(n557), .Z(G1344GAT) );
  NOR2_X1 U624 ( .A1(n568), .A2(n564), .ZN(n562) );
  XOR2_X1 U625 ( .A(KEYINPUT53), .B(KEYINPUT117), .Z(n559) );
  XNOR2_X1 U626 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U628 ( .A(KEYINPUT52), .B(n560), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(G1345GAT) );
  NOR2_X1 U630 ( .A1(n589), .A2(n564), .ZN(n563) );
  XOR2_X1 U631 ( .A(G155GAT), .B(n563), .Z(G1346GAT) );
  NOR2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U633 ( .A(KEYINPUT118), .B(n566), .Z(n567) );
  XNOR2_X1 U634 ( .A(G162GAT), .B(n567), .ZN(G1347GAT) );
  NOR2_X1 U635 ( .A1(n568), .A2(n574), .ZN(n573) );
  XOR2_X1 U636 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n570) );
  XNOR2_X1 U637 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n569) );
  XNOR2_X1 U638 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U639 ( .A(KEYINPUT121), .B(n571), .ZN(n572) );
  XNOR2_X1 U640 ( .A(n573), .B(n572), .ZN(G1349GAT) );
  XOR2_X1 U641 ( .A(G183GAT), .B(KEYINPUT123), .Z(n578) );
  INV_X1 U642 ( .A(n574), .ZN(n576) );
  NAND2_X1 U643 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(G1350GAT) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n593) );
  NOR2_X1 U646 ( .A1(n581), .A2(n593), .ZN(n583) );
  XNOR2_X1 U647 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(G197GAT), .B(n584), .ZN(G1352GAT) );
  XOR2_X1 U650 ( .A(G204GAT), .B(KEYINPUT61), .Z(n588) );
  INV_X1 U651 ( .A(n593), .ZN(n586) );
  NAND2_X1 U652 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(G1353GAT) );
  NOR2_X1 U654 ( .A1(n589), .A2(n593), .ZN(n590) );
  XOR2_X1 U655 ( .A(G211GAT), .B(n590), .Z(G1354GAT) );
  XOR2_X1 U656 ( .A(KEYINPUT125), .B(KEYINPUT62), .Z(n592) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n591) );
  XNOR2_X1 U658 ( .A(n592), .B(n591), .ZN(n596) );
  NOR2_X1 U659 ( .A1(n594), .A2(n593), .ZN(n595) );
  XOR2_X1 U660 ( .A(n596), .B(n595), .Z(G1355GAT) );
endmodule

