// Benchmark "locked_c2670" written by ABC on Sat Dec 16 10:59:00 2023

module locked_c2670 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6,
    G7, G8, G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26,
    G27, G28, G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48,
    G49, G50, G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64,
    G65, G66, G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80,
    G81, G82, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96,
    G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G111, G112,
    G113, G114, G115, G116, G117, G118, G119, G120, G123, G124, G125, G126,
    G127, G128, G129, G130, G131, G132, G135, G136, G137, G138, G139, G140,
    G141, G142, G169, G174, G177, G178, G179, G180, G181, G182, G183, G184,
    G185, G186, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198,
    G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210,
    G211, G212, G213, G214, G215, G239, G240, G241, G242, G243, G244, G245,
    G246, G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
    G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272, G273,
    G274, G275, G276, G277, G278, G279, G452, G483, G543, G559, G567, G651,
    G661, G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966,
    G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078,
    G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435,
    G2438, G2443, G2446, G2451, G2454, G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3,
    G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22, G23, G24,
    G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40, G43, G44,
    G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60, G61, G62,
    G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76, G77, G78,
    G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94,
    G95, G96, G99, G100, G101, G102, G103, G104, G105, G106, G107, G108,
    G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G123, G124,
    G125, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G138,
    G139, G140, G141, G142, G169, G174, G177, G178, G179, G180, G181, G182,
    G183, G184, G185, G186, G189, G190, G191, G192, G193, G194, G195, G196,
    G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208,
    G209, G210, G211, G212, G213, G214, G215, G239, G240, G241, G242, G243,
    G244, G245, G246, G247, G248, G249, G250, G251, G252, G253, G254, G255,
    G256, G257, G262, G263, G264, G265, G266, G267, G268, G269, G270, G271,
    G272, G273, G274, G275, G276, G277, G278, G279, G452, G483, G543, G559,
    G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384, G1956, G1961,
    G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072,
    G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430,
    G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n378, new_n383, new_n387, new_n388, new_n389, new_n390, new_n393,
    new_n394, new_n395, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n408, new_n409,
    new_n410, new_n411, new_n412, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n437, new_n438, new_n439, new_n440,
    new_n441, new_n442, new_n443, new_n446, new_n447, new_n448, new_n449,
    new_n450, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n459, new_n461, new_n462, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n473, new_n474, new_n475, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n503,
    new_n504, new_n507, new_n509, new_n510, new_n511, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n593, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n942;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n378));
  NAND3_X1  g017(.A1(new_n378), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n383));
  XOR2_X1   g022(.A(new_n383), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n387));
  XOR2_X1   g026(.A(new_n387), .B(KEYINPUT2), .Z(new_n388));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n389));
  INV_X1    g028(.A(new_n389), .ZN(new_n390));
  NOR2_X1   g029(.A1(new_n388), .A2(new_n390), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n388), .A2(G2106), .ZN(new_n393));
  NAND2_X1  g032(.A1(new_n390), .A2(G567), .ZN(new_n394));
  NAND2_X1  g033(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g034(.A(new_n395), .ZN(G319));
  OR2_X1    g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n397));
  NAND2_X1  g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n398));
  AOI21_X1  g037(.A(G2105), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g038(.A1(new_n399), .A2(G137), .ZN(new_n400));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n401));
  NAND3_X1  g040(.A1(new_n401), .A2(G125), .A3(G2105), .ZN(new_n402));
  INV_X1    g041(.A(G2104), .ZN(new_n403));
  NOR2_X1   g042(.A1(new_n403), .A2(G2105), .ZN(new_n404));
  AND2_X1   g043(.A1(G113), .A2(G2104), .ZN(new_n405));
  AOI22_X1  g044(.A1(new_n404), .A2(G101), .B1(new_n405), .B2(G2105), .ZN(new_n406));
  AND3_X1   g045(.A1(new_n400), .A2(new_n402), .A3(new_n406), .ZN(G160));
  NAND2_X1  g046(.A1(new_n399), .A2(G136), .ZN(new_n408));
  NAND3_X1  g047(.A1(new_n401), .A2(G124), .A3(G2105), .ZN(new_n409));
  NAND3_X1  g048(.A1(G112), .A2(G2104), .A3(G2105), .ZN(new_n410));
  NAND2_X1  g049(.A1(new_n404), .A2(G100), .ZN(new_n411));
  NAND4_X1  g050(.A1(new_n408), .A2(new_n409), .A3(new_n410), .A4(new_n411), .ZN(new_n412));
  INV_X1    g051(.A(new_n412), .ZN(G162));
  AND2_X1   g052(.A1(G126), .A2(G2105), .ZN(new_n414));
  AND2_X1   g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n415));
  NOR2_X1   g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n416));
  OAI21_X1  g055(.A(new_n414), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g056(.A1(G114), .A2(G2104), .A3(G2105), .ZN(new_n418));
  INV_X1    g057(.A(G2105), .ZN(new_n419));
  NAND3_X1  g058(.A1(new_n419), .A2(G102), .A3(G2104), .ZN(new_n420));
  NAND3_X1  g059(.A1(new_n417), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  OAI211_X1 g060(.A(G138), .B(new_n419), .C1(new_n415), .C2(new_n416), .ZN(new_n422));
  NAND2_X1  g061(.A1(new_n422), .A2(KEYINPUT4), .ZN(new_n423));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n424));
  NAND4_X1  g063(.A1(new_n401), .A2(new_n424), .A3(G138), .A4(new_n419), .ZN(new_n425));
  AOI21_X1  g064(.A(new_n421), .B1(new_n423), .B2(new_n425), .ZN(G164));
  XNOR2_X1  g065(.A(KEYINPUT5), .B(G543), .ZN(new_n427));
  AOI22_X1  g066(.A1(new_n427), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n428));
  INV_X1    g067(.A(G651), .ZN(new_n429));
  NOR2_X1   g068(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g069(.A(KEYINPUT6), .B(G651), .ZN(new_n431));
  NAND3_X1  g070(.A1(new_n431), .A2(G50), .A3(G543), .ZN(new_n432));
  NAND2_X1  g071(.A1(new_n427), .A2(new_n431), .ZN(new_n433));
  INV_X1    g072(.A(G88), .ZN(new_n434));
  OAI21_X1  g073(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NOR2_X1   g074(.A1(new_n430), .A2(new_n435), .ZN(G166));
  AND2_X1   g075(.A1(new_n427), .A2(new_n431), .ZN(new_n437));
  AND2_X1   g076(.A1(new_n437), .A2(G89), .ZN(new_n438));
  NAND3_X1  g077(.A1(new_n427), .A2(G63), .A3(G651), .ZN(new_n439));
  NAND3_X1  g078(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n440));
  XNOR2_X1  g079(.A(new_n440), .B(KEYINPUT7), .ZN(new_n441));
  NAND3_X1  g080(.A1(new_n431), .A2(G51), .A3(G543), .ZN(new_n442));
  NAND3_X1  g081(.A1(new_n439), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  OR2_X1    g082(.A1(new_n438), .A2(new_n443), .ZN(G286));
  INV_X1    g083(.A(G286), .ZN(G168));
  AOI22_X1  g084(.A1(new_n427), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n446));
  NOR2_X1   g085(.A1(new_n446), .A2(new_n429), .ZN(new_n447));
  NAND3_X1  g086(.A1(new_n431), .A2(G52), .A3(G543), .ZN(new_n448));
  INV_X1    g087(.A(G90), .ZN(new_n449));
  OAI21_X1  g088(.A(new_n448), .B1(new_n433), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g089(.A1(new_n447), .A2(new_n450), .ZN(G171));
  AOI22_X1  g090(.A1(new_n427), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n452));
  NOR2_X1   g091(.A1(new_n452), .A2(new_n429), .ZN(new_n453));
  NAND3_X1  g092(.A1(new_n431), .A2(G43), .A3(G543), .ZN(new_n454));
  INV_X1    g093(.A(G81), .ZN(new_n455));
  OAI21_X1  g094(.A(new_n454), .B1(new_n433), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g095(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g096(.A1(new_n457), .A2(G860), .ZN(G153));
  AND3_X1   g097(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n459));
  NAND2_X1  g098(.A1(new_n459), .A2(G36), .ZN(G176));
  NAND2_X1  g099(.A1(G1), .A2(G3), .ZN(new_n461));
  XNOR2_X1  g100(.A(new_n461), .B(KEYINPUT8), .ZN(new_n462));
  NAND2_X1  g101(.A1(new_n459), .A2(new_n462), .ZN(G188));
  AOI22_X1  g102(.A1(new_n427), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n464));
  INV_X1    g103(.A(G91), .ZN(new_n465));
  OAI22_X1  g104(.A1(new_n464), .A2(new_n429), .B1(new_n433), .B2(new_n465), .ZN(new_n466));
  INV_X1    g105(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g106(.A1(new_n431), .A2(G53), .A3(G543), .ZN(new_n468));
  XNOR2_X1  g107(.A(new_n468), .B(KEYINPUT9), .ZN(new_n469));
  NAND2_X1  g108(.A1(new_n467), .A2(new_n469), .ZN(G299));
  INV_X1    g109(.A(G171), .ZN(G301));
  INV_X1    g110(.A(G166), .ZN(G303));
  OAI21_X1  g111(.A(G651), .B1(new_n427), .B2(G74), .ZN(new_n473));
  NAND3_X1  g112(.A1(new_n431), .A2(G49), .A3(G543), .ZN(new_n474));
  INV_X1    g113(.A(G87), .ZN(new_n475));
  OAI211_X1 g114(.A(new_n473), .B(new_n474), .C1(new_n475), .C2(new_n433), .ZN(G288));
  AOI22_X1  g115(.A1(new_n427), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n477));
  NOR2_X1   g116(.A1(new_n477), .A2(new_n429), .ZN(new_n478));
  NAND3_X1  g117(.A1(new_n431), .A2(G48), .A3(G543), .ZN(new_n479));
  INV_X1    g118(.A(G86), .ZN(new_n480));
  OAI21_X1  g119(.A(new_n479), .B1(new_n433), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g120(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  INV_X1    g121(.A(new_n482), .ZN(G305));
  NAND3_X1  g122(.A1(new_n431), .A2(G47), .A3(G543), .ZN(new_n484));
  INV_X1    g123(.A(G85), .ZN(new_n485));
  AOI22_X1  g124(.A1(new_n427), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n486));
  OAI221_X1 g125(.A(new_n484), .B1(new_n433), .B2(new_n485), .C1(new_n486), .C2(new_n429), .ZN(G290));
  NAND2_X1  g126(.A1(G301), .A2(G868), .ZN(new_n488));
  NAND3_X1  g127(.A1(new_n437), .A2(KEYINPUT10), .A3(G92), .ZN(new_n489));
  INV_X1    g128(.A(KEYINPUT10), .ZN(new_n490));
  INV_X1    g129(.A(G92), .ZN(new_n491));
  OAI21_X1  g130(.A(new_n490), .B1(new_n433), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g131(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g132(.A1(new_n427), .A2(G66), .ZN(new_n494));
  NAND2_X1  g133(.A1(G79), .A2(G543), .ZN(new_n495));
  NAND2_X1  g134(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AND2_X1   g135(.A1(G54), .A2(G543), .ZN(new_n497));
  AOI22_X1  g136(.A1(new_n496), .A2(G651), .B1(new_n431), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g137(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  INV_X1    g138(.A(new_n499), .ZN(new_n500));
  OAI21_X1  g139(.A(new_n488), .B1(new_n500), .B2(G868), .ZN(G284));
  OAI21_X1  g140(.A(new_n488), .B1(new_n500), .B2(G868), .ZN(G321));
  INV_X1    g141(.A(G868), .ZN(new_n503));
  NAND2_X1  g142(.A1(G299), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g143(.A(new_n504), .B1(G168), .B2(new_n503), .ZN(G297));
  OAI21_X1  g144(.A(new_n504), .B1(G168), .B2(new_n503), .ZN(G280));
  INV_X1    g145(.A(G559), .ZN(new_n507));
  OAI21_X1  g146(.A(new_n500), .B1(new_n507), .B2(G860), .ZN(G148));
  INV_X1    g147(.A(new_n457), .ZN(new_n509));
  NAND2_X1  g148(.A1(new_n509), .A2(new_n503), .ZN(new_n510));
  NOR2_X1   g149(.A1(new_n499), .A2(G559), .ZN(new_n511));
  OAI21_X1  g150(.A(new_n510), .B1(new_n511), .B2(new_n503), .ZN(G323));
  XNOR2_X1  g151(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g152(.A1(new_n399), .A2(G2104), .ZN(new_n514));
  XNOR2_X1  g153(.A(new_n514), .B(KEYINPUT12), .ZN(new_n515));
  XNOR2_X1  g154(.A(new_n515), .B(G2100), .ZN(new_n516));
  XNOR2_X1  g155(.A(new_n516), .B(KEYINPUT13), .ZN(new_n517));
  NAND2_X1  g156(.A1(new_n399), .A2(G135), .ZN(new_n518));
  NAND3_X1  g157(.A1(new_n401), .A2(G123), .A3(G2105), .ZN(new_n519));
  AND2_X1   g158(.A1(G111), .A2(G2104), .ZN(new_n520));
  AOI22_X1  g159(.A1(new_n404), .A2(G99), .B1(new_n520), .B2(G2105), .ZN(new_n521));
  NAND3_X1  g160(.A1(new_n518), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  XOR2_X1   g161(.A(new_n522), .B(G2096), .Z(new_n523));
  NAND2_X1  g162(.A1(new_n517), .A2(new_n523), .ZN(G156));
  XOR2_X1   g163(.A(G2427), .B(G2430), .Z(new_n525));
  XNOR2_X1  g164(.A(new_n525), .B(KEYINPUT15), .ZN(new_n526));
  XOR2_X1   g165(.A(G2435), .B(G2438), .Z(new_n527));
  OR2_X1    g166(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g167(.A1(new_n526), .A2(new_n527), .ZN(new_n529));
  NAND3_X1  g168(.A1(new_n528), .A2(KEYINPUT14), .A3(new_n529), .ZN(new_n530));
  XOR2_X1   g169(.A(G2443), .B(G2446), .Z(new_n531));
  XNOR2_X1  g170(.A(new_n530), .B(new_n531), .ZN(new_n532));
  XNOR2_X1  g171(.A(G2451), .B(G2454), .ZN(new_n533));
  XNOR2_X1  g172(.A(new_n533), .B(KEYINPUT16), .ZN(new_n534));
  XNOR2_X1  g173(.A(G1341), .B(G1348), .ZN(new_n535));
  XNOR2_X1  g174(.A(new_n534), .B(new_n535), .ZN(new_n536));
  XNOR2_X1  g175(.A(new_n532), .B(new_n536), .ZN(new_n537));
  AND2_X1   g176(.A1(new_n537), .A2(G14), .ZN(G401));
  XOR2_X1   g177(.A(G2067), .B(G2678), .Z(new_n539));
  INV_X1    g178(.A(new_n539), .ZN(new_n540));
  XOR2_X1   g179(.A(G2084), .B(G2090), .Z(new_n541));
  XNOR2_X1  g180(.A(G2072), .B(G2078), .ZN(new_n542));
  NAND3_X1  g181(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  XOR2_X1   g182(.A(new_n543), .B(KEYINPUT18), .Z(new_n544));
  XOR2_X1   g183(.A(new_n542), .B(KEYINPUT17), .Z(new_n545));
  NAND3_X1  g184(.A1(new_n545), .A2(new_n541), .A3(new_n539), .ZN(new_n546));
  AND2_X1   g185(.A1(new_n539), .A2(new_n542), .ZN(new_n547));
  AOI21_X1  g186(.A(new_n547), .B1(new_n545), .B2(new_n540), .ZN(new_n548));
  OAI211_X1 g187(.A(new_n544), .B(new_n546), .C1(new_n548), .C2(new_n541), .ZN(new_n549));
  XOR2_X1   g188(.A(G2096), .B(G2100), .Z(new_n550));
  XNOR2_X1  g189(.A(new_n549), .B(new_n550), .ZN(G227));
  XNOR2_X1  g190(.A(G1981), .B(G1986), .ZN(new_n552));
  XNOR2_X1  g191(.A(new_n552), .B(KEYINPUT21), .ZN(new_n553));
  XOR2_X1   g192(.A(G1991), .B(G1996), .Z(new_n554));
  XNOR2_X1  g193(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XOR2_X1   g194(.A(new_n555), .B(KEYINPUT22), .Z(new_n556));
  XNOR2_X1  g195(.A(G1971), .B(G1976), .ZN(new_n557));
  XNOR2_X1  g196(.A(new_n557), .B(KEYINPUT19), .ZN(new_n558));
  XNOR2_X1  g197(.A(G1956), .B(G2474), .ZN(new_n559));
  XNOR2_X1  g198(.A(G1961), .B(G1966), .ZN(new_n560));
  OR2_X1    g199(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g200(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  XOR2_X1   g201(.A(new_n562), .B(KEYINPUT20), .Z(new_n563));
  NAND2_X1  g202(.A1(new_n558), .A2(new_n561), .ZN(new_n564));
  NAND2_X1  g203(.A1(new_n559), .A2(new_n560), .ZN(new_n565));
  XNOR2_X1  g204(.A(new_n564), .B(new_n565), .ZN(new_n566));
  NAND2_X1  g205(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g206(.A(new_n556), .B(new_n567), .ZN(G229));
  INV_X1    g207(.A(G16), .ZN(new_n569));
  NAND2_X1  g208(.A1(new_n569), .A2(G21), .ZN(new_n570));
  OAI21_X1  g209(.A(new_n570), .B1(G168), .B2(new_n569), .ZN(new_n571));
  XOR2_X1   g210(.A(new_n571), .B(G1966), .Z(new_n572));
  XNOR2_X1  g211(.A(KEYINPUT31), .B(G11), .ZN(new_n573));
  AND2_X1   g212(.A1(new_n522), .A2(G29), .ZN(new_n574));
  INV_X1    g213(.A(G29), .ZN(new_n575));
  OAI21_X1  g214(.A(new_n575), .B1(KEYINPUT30), .B2(G28), .ZN(new_n576));
  AOI21_X1  g215(.A(new_n576), .B1(KEYINPUT30), .B2(G28), .ZN(new_n577));
  OAI21_X1  g216(.A(new_n573), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g217(.A1(new_n569), .A2(G5), .ZN(new_n579));
  OAI21_X1  g218(.A(new_n579), .B1(G171), .B2(new_n569), .ZN(new_n580));
  AOI21_X1  g219(.A(new_n578), .B1(new_n580), .B2(G1961), .ZN(new_n581));
  NAND2_X1  g220(.A1(new_n575), .A2(G35), .ZN(new_n582));
  OAI21_X1  g221(.A(new_n582), .B1(G162), .B2(new_n575), .ZN(new_n583));
  XNOR2_X1  g222(.A(new_n583), .B(KEYINPUT29), .ZN(new_n584));
  NAND2_X1  g223(.A1(new_n584), .A2(G2090), .ZN(new_n585));
  NAND2_X1  g224(.A1(new_n569), .A2(G19), .ZN(new_n586));
  OAI21_X1  g225(.A(new_n586), .B1(new_n457), .B2(new_n569), .ZN(new_n587));
  XOR2_X1   g226(.A(new_n587), .B(G1341), .Z(new_n588));
  NAND4_X1  g227(.A1(new_n572), .A2(new_n581), .A3(new_n585), .A4(new_n588), .ZN(new_n589));
  NAND2_X1  g228(.A1(new_n404), .A2(G103), .ZN(new_n590));
  INV_X1    g229(.A(KEYINPUT25), .ZN(new_n591));
  NAND2_X1  g230(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g231(.A1(new_n404), .A2(KEYINPUT25), .A3(G103), .ZN(new_n593));
  AOI22_X1  g232(.A1(new_n592), .A2(new_n593), .B1(new_n399), .B2(G139), .ZN(new_n594));
  AOI22_X1  g233(.A1(new_n401), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n595));
  OAI21_X1  g234(.A(new_n594), .B1(new_n419), .B2(new_n595), .ZN(new_n596));
  MUX2_X1   g235(.A(G33), .B(new_n596), .S(G29), .Z(new_n597));
  XOR2_X1   g236(.A(new_n597), .B(G2072), .Z(new_n598));
  NAND2_X1  g237(.A1(new_n575), .A2(G27), .ZN(new_n599));
  OAI21_X1  g238(.A(new_n599), .B1(G164), .B2(new_n575), .ZN(new_n600));
  INV_X1    g239(.A(G2078), .ZN(new_n601));
  XNOR2_X1  g240(.A(new_n600), .B(new_n601), .ZN(new_n602));
  OAI211_X1 g241(.A(new_n598), .B(new_n602), .C1(G2090), .C2(new_n584), .ZN(new_n603));
  NAND2_X1  g242(.A1(new_n569), .A2(G4), .ZN(new_n604));
  OAI21_X1  g243(.A(new_n604), .B1(new_n500), .B2(new_n569), .ZN(new_n605));
  INV_X1    g244(.A(G1348), .ZN(new_n606));
  XNOR2_X1  g245(.A(new_n605), .B(new_n606), .ZN(new_n607));
  NAND2_X1  g246(.A1(new_n569), .A2(G20), .ZN(new_n608));
  XOR2_X1   g247(.A(new_n608), .B(KEYINPUT23), .Z(new_n609));
  AOI21_X1  g248(.A(new_n609), .B1(G299), .B2(G16), .ZN(new_n610));
  XNOR2_X1  g249(.A(new_n610), .B(G1956), .ZN(new_n611));
  NAND2_X1  g250(.A1(new_n575), .A2(G26), .ZN(new_n612));
  XOR2_X1   g251(.A(new_n612), .B(KEYINPUT28), .Z(new_n613));
  NAND2_X1  g252(.A1(new_n399), .A2(G140), .ZN(new_n614));
  NAND3_X1  g253(.A1(new_n401), .A2(G128), .A3(G2105), .ZN(new_n615));
  AND2_X1   g254(.A1(G116), .A2(G2104), .ZN(new_n616));
  AOI22_X1  g255(.A1(new_n404), .A2(G104), .B1(new_n616), .B2(G2105), .ZN(new_n617));
  NAND3_X1  g256(.A1(new_n614), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g257(.A(new_n613), .B1(new_n618), .B2(G29), .ZN(new_n619));
  INV_X1    g258(.A(G2067), .ZN(new_n620));
  XNOR2_X1  g259(.A(new_n619), .B(new_n620), .ZN(new_n621));
  OAI21_X1  g260(.A(new_n575), .B1(KEYINPUT24), .B2(G34), .ZN(new_n622));
  AOI21_X1  g261(.A(new_n622), .B1(KEYINPUT24), .B2(G34), .ZN(new_n623));
  NAND3_X1  g262(.A1(new_n400), .A2(new_n402), .A3(new_n406), .ZN(new_n624));
  AOI21_X1  g263(.A(new_n623), .B1(new_n624), .B2(G29), .ZN(new_n625));
  INV_X1    g264(.A(G2084), .ZN(new_n626));
  XNOR2_X1  g265(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NOR2_X1   g266(.A1(new_n580), .A2(G1961), .ZN(new_n628));
  NOR3_X1   g267(.A1(new_n621), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND3_X1  g268(.A1(new_n607), .A2(new_n611), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g269(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n631));
  XOR2_X1   g270(.A(new_n631), .B(KEYINPUT26), .Z(new_n632));
  NAND2_X1  g271(.A1(new_n399), .A2(G141), .ZN(new_n633));
  NAND3_X1  g272(.A1(new_n401), .A2(G129), .A3(G2105), .ZN(new_n634));
  NAND2_X1  g273(.A1(new_n404), .A2(G105), .ZN(new_n635));
  NAND4_X1  g274(.A1(new_n632), .A2(new_n633), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  MUX2_X1   g275(.A(G32), .B(new_n636), .S(G29), .Z(new_n637));
  INV_X1    g276(.A(G1996), .ZN(new_n638));
  XNOR2_X1  g277(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g278(.A(new_n639), .B(KEYINPUT27), .ZN(new_n640));
  NOR4_X1   g279(.A1(new_n589), .A2(new_n603), .A3(new_n630), .A4(new_n640), .ZN(new_n641));
  INV_X1    g280(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g281(.A1(new_n569), .A2(G6), .ZN(new_n643));
  OAI21_X1  g282(.A(new_n643), .B1(new_n482), .B2(new_n569), .ZN(new_n644));
  XNOR2_X1  g283(.A(new_n644), .B(KEYINPUT32), .ZN(new_n645));
  INV_X1    g284(.A(G1981), .ZN(new_n646));
  XNOR2_X1  g285(.A(new_n645), .B(new_n646), .ZN(new_n647));
  MUX2_X1   g286(.A(G23), .B(G288), .S(G16), .Z(new_n648));
  XNOR2_X1  g287(.A(new_n648), .B(G1976), .ZN(new_n649));
  XNOR2_X1  g288(.A(new_n649), .B(KEYINPUT33), .ZN(new_n650));
  NAND2_X1  g289(.A1(new_n569), .A2(G22), .ZN(new_n651));
  OAI21_X1  g290(.A(new_n651), .B1(G166), .B2(new_n569), .ZN(new_n652));
  INV_X1    g291(.A(G1971), .ZN(new_n653));
  XNOR2_X1  g292(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NAND3_X1  g293(.A1(new_n647), .A2(new_n650), .A3(new_n654), .ZN(new_n655));
  OR2_X1    g294(.A1(new_n655), .A2(KEYINPUT34), .ZN(new_n656));
  NAND2_X1  g295(.A1(new_n655), .A2(KEYINPUT34), .ZN(new_n657));
  NAND2_X1  g296(.A1(new_n399), .A2(G131), .ZN(new_n658));
  NAND3_X1  g297(.A1(new_n401), .A2(G119), .A3(G2105), .ZN(new_n659));
  NAND3_X1  g298(.A1(G107), .A2(G2104), .A3(G2105), .ZN(new_n660));
  NAND2_X1  g299(.A1(new_n404), .A2(G95), .ZN(new_n661));
  NAND4_X1  g300(.A1(new_n658), .A2(new_n659), .A3(new_n660), .A4(new_n661), .ZN(new_n662));
  MUX2_X1   g301(.A(G25), .B(new_n662), .S(G29), .Z(new_n663));
  XNOR2_X1  g302(.A(KEYINPUT35), .B(G1991), .ZN(new_n664));
  XNOR2_X1  g303(.A(new_n663), .B(new_n664), .ZN(new_n665));
  AND2_X1   g304(.A1(new_n569), .A2(G24), .ZN(new_n666));
  AOI21_X1  g305(.A(new_n666), .B1(G290), .B2(G16), .ZN(new_n667));
  INV_X1    g306(.A(G1986), .ZN(new_n668));
  AND2_X1   g307(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g308(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  NOR3_X1   g309(.A1(new_n665), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND3_X1  g310(.A1(new_n656), .A2(new_n657), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g311(.A1(new_n672), .A2(KEYINPUT36), .ZN(new_n673));
  AND2_X1   g312(.A1(new_n657), .A2(new_n671), .ZN(new_n674));
  INV_X1    g313(.A(KEYINPUT36), .ZN(new_n675));
  NAND3_X1  g314(.A1(new_n674), .A2(new_n675), .A3(new_n656), .ZN(new_n676));
  AOI21_X1  g315(.A(new_n642), .B1(new_n673), .B2(new_n676), .ZN(G311));
  AOI21_X1  g316(.A(new_n675), .B1(new_n674), .B2(new_n656), .ZN(new_n678));
  AND4_X1   g317(.A1(new_n675), .A2(new_n656), .A3(new_n657), .A4(new_n671), .ZN(new_n679));
  OAI21_X1  g318(.A(new_n641), .B1(new_n678), .B2(new_n679), .ZN(G150));
  AOI22_X1  g319(.A1(new_n427), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n681));
  NOR2_X1   g320(.A1(new_n681), .A2(new_n429), .ZN(new_n682));
  NAND3_X1  g321(.A1(new_n431), .A2(G55), .A3(G543), .ZN(new_n683));
  INV_X1    g322(.A(G93), .ZN(new_n684));
  OAI21_X1  g323(.A(new_n683), .B1(new_n433), .B2(new_n684), .ZN(new_n685));
  NOR2_X1   g324(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  INV_X1    g325(.A(G860), .ZN(new_n687));
  NOR2_X1   g326(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g327(.A(new_n688), .B(KEYINPUT37), .ZN(new_n689));
  NOR2_X1   g328(.A1(new_n499), .A2(new_n507), .ZN(new_n690));
  XNOR2_X1  g329(.A(new_n690), .B(new_n509), .ZN(new_n691));
  XNOR2_X1  g330(.A(new_n691), .B(KEYINPUT38), .ZN(new_n692));
  XNOR2_X1  g331(.A(new_n692), .B(new_n686), .ZN(new_n693));
  INV_X1    g332(.A(KEYINPUT39), .ZN(new_n694));
  AND2_X1   g333(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g334(.A(new_n687), .B1(new_n693), .B2(new_n694), .ZN(new_n696));
  OAI21_X1  g335(.A(new_n689), .B1(new_n695), .B2(new_n696), .ZN(G145));
  INV_X1    g336(.A(G37), .ZN(new_n698));
  NAND2_X1  g337(.A1(new_n423), .A2(new_n425), .ZN(new_n699));
  INV_X1    g338(.A(new_n421), .ZN(new_n700));
  NAND2_X1  g339(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g340(.A(new_n596), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g341(.A(new_n636), .B(new_n618), .ZN(new_n703));
  XNOR2_X1  g342(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g343(.A1(new_n399), .A2(G142), .ZN(new_n705));
  NAND3_X1  g344(.A1(new_n401), .A2(G130), .A3(G2105), .ZN(new_n706));
  NAND3_X1  g345(.A1(G118), .A2(G2104), .A3(G2105), .ZN(new_n707));
  NAND2_X1  g346(.A1(new_n404), .A2(G106), .ZN(new_n708));
  NAND4_X1  g347(.A1(new_n705), .A2(new_n706), .A3(new_n707), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g348(.A(new_n662), .B(new_n709), .ZN(new_n710));
  XNOR2_X1  g349(.A(new_n704), .B(new_n710), .ZN(new_n711));
  XNOR2_X1  g350(.A(new_n515), .B(new_n522), .ZN(new_n712));
  XNOR2_X1  g351(.A(G160), .B(new_n412), .ZN(new_n713));
  XNOR2_X1  g352(.A(new_n712), .B(new_n713), .ZN(new_n714));
  AND2_X1   g353(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g354(.A1(new_n711), .A2(new_n714), .ZN(new_n716));
  OAI21_X1  g355(.A(new_n698), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  XNOR2_X1  g356(.A(new_n717), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g357(.A(new_n482), .B(G290), .ZN(new_n719));
  XNOR2_X1  g358(.A(G166), .B(G288), .ZN(new_n720));
  XOR2_X1   g359(.A(new_n719), .B(new_n720), .Z(new_n721));
  XNOR2_X1  g360(.A(new_n457), .B(new_n686), .ZN(new_n722));
  NAND2_X1  g361(.A1(G299), .A2(new_n499), .ZN(new_n723));
  NAND4_X1  g362(.A1(new_n467), .A2(new_n493), .A3(new_n469), .A4(new_n498), .ZN(new_n724));
  AOI21_X1  g363(.A(KEYINPUT41), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g364(.A(new_n725), .ZN(new_n726));
  NAND3_X1  g365(.A1(new_n723), .A2(KEYINPUT41), .A3(new_n724), .ZN(new_n727));
  AOI21_X1  g366(.A(new_n722), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g367(.A1(new_n723), .A2(new_n724), .ZN(new_n729));
  NAND2_X1  g368(.A1(new_n729), .A2(new_n722), .ZN(new_n730));
  INV_X1    g369(.A(new_n730), .ZN(new_n731));
  OAI22_X1  g370(.A1(new_n728), .A2(new_n731), .B1(G559), .B2(new_n499), .ZN(new_n732));
  INV_X1    g371(.A(new_n722), .ZN(new_n733));
  AOI21_X1  g372(.A(new_n733), .B1(new_n726), .B2(new_n727), .ZN(new_n734));
  NAND2_X1  g373(.A1(new_n733), .A2(new_n729), .ZN(new_n735));
  INV_X1    g374(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g375(.A(new_n511), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  INV_X1    g376(.A(KEYINPUT42), .ZN(new_n738));
  AND3_X1   g377(.A1(new_n732), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g378(.A(new_n738), .B1(new_n732), .B2(new_n737), .ZN(new_n740));
  OAI21_X1  g379(.A(new_n721), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g380(.A1(new_n741), .A2(G868), .ZN(new_n742));
  NOR3_X1   g381(.A1(new_n739), .A2(new_n740), .A3(new_n721), .ZN(new_n743));
  OAI22_X1  g382(.A1(new_n742), .A2(new_n743), .B1(G868), .B2(new_n686), .ZN(G295));
  OAI22_X1  g383(.A1(new_n742), .A2(new_n743), .B1(G868), .B2(new_n686), .ZN(G331));
  INV_X1    g384(.A(KEYINPUT44), .ZN(new_n746));
  INV_X1    g385(.A(KEYINPUT43), .ZN(new_n747));
  XNOR2_X1  g386(.A(G286), .B(G171), .ZN(new_n748));
  INV_X1    g387(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g388(.A(new_n749), .B1(new_n734), .B2(new_n736), .ZN(new_n750));
  OAI21_X1  g389(.A(new_n748), .B1(new_n728), .B2(new_n731), .ZN(new_n751));
  NAND2_X1  g390(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g391(.A(new_n721), .ZN(new_n753));
  AOI21_X1  g392(.A(G37), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g393(.A1(new_n750), .A2(new_n751), .A3(new_n721), .ZN(new_n755));
  AOI21_X1  g394(.A(new_n747), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g395(.A(new_n727), .ZN(new_n757));
  OAI21_X1  g396(.A(new_n722), .B1(new_n757), .B2(new_n725), .ZN(new_n758));
  AOI21_X1  g397(.A(new_n748), .B1(new_n758), .B2(new_n735), .ZN(new_n759));
  OAI21_X1  g398(.A(new_n733), .B1(new_n757), .B2(new_n725), .ZN(new_n760));
  AOI21_X1  g399(.A(new_n749), .B1(new_n760), .B2(new_n730), .ZN(new_n761));
  OAI21_X1  g400(.A(new_n753), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  AND4_X1   g401(.A1(new_n747), .A2(new_n762), .A3(new_n755), .A4(new_n698), .ZN(new_n763));
  OAI21_X1  g402(.A(new_n746), .B1(new_n756), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g403(.A1(new_n754), .A2(new_n747), .A3(new_n755), .ZN(new_n765));
  NAND3_X1  g404(.A1(new_n762), .A2(new_n755), .A3(new_n698), .ZN(new_n766));
  NAND2_X1  g405(.A1(new_n766), .A2(KEYINPUT43), .ZN(new_n767));
  NAND3_X1  g406(.A1(new_n765), .A2(new_n767), .A3(KEYINPUT44), .ZN(new_n768));
  NAND2_X1  g407(.A1(new_n764), .A2(new_n768), .ZN(G397));
  INV_X1    g408(.A(G40), .ZN(new_n770));
  NOR2_X1   g409(.A1(new_n624), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g410(.A(G1384), .B1(new_n699), .B2(new_n700), .ZN(new_n772));
  INV_X1    g411(.A(KEYINPUT50), .ZN(new_n773));
  OAI21_X1  g412(.A(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR3_X1   g413(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n775));
  OAI21_X1  g414(.A(new_n606), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g415(.A1(new_n772), .A2(new_n771), .ZN(new_n777));
  INV_X1    g416(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g417(.A1(new_n778), .A2(new_n620), .ZN(new_n779));
  NAND3_X1  g418(.A1(new_n776), .A2(new_n779), .A3(new_n500), .ZN(new_n780));
  INV_X1    g419(.A(KEYINPUT60), .ZN(new_n781));
  NAND2_X1  g420(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g421(.A1(new_n776), .A2(new_n779), .ZN(new_n783));
  NAND2_X1  g422(.A1(new_n783), .A2(new_n499), .ZN(new_n784));
  NAND4_X1  g423(.A1(new_n776), .A2(new_n779), .A3(KEYINPUT60), .A4(new_n500), .ZN(new_n785));
  NAND3_X1  g424(.A1(new_n782), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  XNOR2_X1  g425(.A(KEYINPUT58), .B(G1341), .ZN(new_n787));
  AOI21_X1  g426(.A(new_n787), .B1(new_n772), .B2(new_n771), .ZN(new_n788));
  NAND2_X1  g427(.A1(G160), .A2(G40), .ZN(new_n789));
  INV_X1    g428(.A(KEYINPUT45), .ZN(new_n790));
  INV_X1    g429(.A(G1384), .ZN(new_n791));
  NAND3_X1  g430(.A1(new_n701), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  OAI21_X1  g431(.A(KEYINPUT45), .B1(G164), .B2(G1384), .ZN(new_n793));
  AOI21_X1  g432(.A(new_n789), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g433(.A(new_n788), .B1(new_n794), .B2(new_n638), .ZN(new_n795));
  OAI21_X1  g434(.A(KEYINPUT59), .B1(new_n795), .B2(new_n509), .ZN(new_n796));
  INV_X1    g435(.A(KEYINPUT59), .ZN(new_n797));
  AOI211_X1 g436(.A(G1996), .B(new_n789), .C1(new_n792), .C2(new_n793), .ZN(new_n798));
  OAI211_X1 g437(.A(new_n797), .B(new_n457), .C1(new_n798), .C2(new_n788), .ZN(new_n799));
  NAND2_X1  g438(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  INV_X1    g439(.A(KEYINPUT61), .ZN(new_n801));
  INV_X1    g440(.A(G1956), .ZN(new_n802));
  OAI21_X1  g441(.A(new_n802), .B1(new_n774), .B2(new_n775), .ZN(new_n803));
  XOR2_X1   g442(.A(KEYINPUT56), .B(G2072), .Z(new_n804));
  INV_X1    g443(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g444(.A(new_n790), .B1(new_n701), .B2(new_n791), .ZN(new_n806));
  AOI211_X1 g445(.A(KEYINPUT45), .B(G1384), .C1(new_n699), .C2(new_n700), .ZN(new_n807));
  OAI211_X1 g446(.A(new_n771), .B(new_n805), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  INV_X1    g447(.A(KEYINPUT9), .ZN(new_n809));
  XNOR2_X1  g448(.A(new_n468), .B(new_n809), .ZN(new_n810));
  NOR3_X1   g449(.A1(new_n810), .A2(new_n466), .A3(KEYINPUT57), .ZN(new_n811));
  INV_X1    g450(.A(KEYINPUT57), .ZN(new_n812));
  AOI21_X1  g451(.A(new_n812), .B1(new_n467), .B2(new_n469), .ZN(new_n813));
  NOR2_X1   g452(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  AND3_X1   g453(.A1(new_n803), .A2(new_n808), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g454(.A(new_n814), .B1(new_n803), .B2(new_n808), .ZN(new_n816));
  OAI21_X1  g455(.A(new_n801), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g456(.A1(new_n803), .A2(new_n808), .ZN(new_n818));
  INV_X1    g457(.A(new_n814), .ZN(new_n819));
  NAND2_X1  g458(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g459(.A1(new_n803), .A2(new_n808), .A3(new_n814), .ZN(new_n821));
  NAND3_X1  g460(.A1(new_n820), .A2(KEYINPUT61), .A3(new_n821), .ZN(new_n822));
  NAND4_X1  g461(.A1(new_n786), .A2(new_n800), .A3(new_n817), .A4(new_n822), .ZN(new_n823));
  AOI21_X1  g462(.A(new_n499), .B1(new_n776), .B2(new_n779), .ZN(new_n824));
  AOI21_X1  g463(.A(new_n816), .B1(new_n824), .B2(new_n821), .ZN(new_n825));
  NAND2_X1  g464(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g465(.A1(new_n772), .A2(new_n773), .ZN(new_n827));
  OAI21_X1  g466(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n828));
  NAND4_X1  g467(.A1(new_n827), .A2(new_n828), .A3(new_n626), .A4(new_n771), .ZN(new_n829));
  OAI21_X1  g468(.A(new_n829), .B1(new_n794), .B2(G1966), .ZN(new_n830));
  AND3_X1   g469(.A1(new_n830), .A2(G8), .A3(G286), .ZN(new_n831));
  NAND2_X1  g470(.A1(new_n830), .A2(G8), .ZN(new_n832));
  INV_X1    g471(.A(KEYINPUT51), .ZN(new_n833));
  NAND2_X1  g472(.A1(G286), .A2(G8), .ZN(new_n834));
  NAND3_X1  g473(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  OAI211_X1 g474(.A(KEYINPUT51), .B(G8), .C1(new_n830), .C2(G286), .ZN(new_n836));
  AOI21_X1  g475(.A(new_n831), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g476(.A1(new_n794), .A2(G1971), .ZN(new_n838));
  NOR3_X1   g477(.A1(new_n774), .A2(G2090), .A3(new_n775), .ZN(new_n839));
  OAI21_X1  g478(.A(G8), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g479(.A1(G303), .A2(G8), .ZN(new_n841));
  INV_X1    g480(.A(KEYINPUT55), .ZN(new_n842));
  XNOR2_X1  g481(.A(new_n841), .B(new_n842), .ZN(new_n843));
  INV_X1    g482(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g483(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  INV_X1    g484(.A(G8), .ZN(new_n846));
  AOI21_X1  g485(.A(new_n846), .B1(new_n772), .B2(new_n771), .ZN(new_n847));
  INV_X1    g486(.A(G1976), .ZN(new_n848));
  OR2_X1    g487(.A1(G288), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g488(.A1(G288), .A2(new_n848), .ZN(new_n850));
  INV_X1    g489(.A(KEYINPUT52), .ZN(new_n851));
  NAND2_X1  g490(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AND3_X1   g491(.A1(new_n847), .A2(new_n849), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g492(.A(KEYINPUT52), .B1(new_n847), .B2(new_n849), .ZN(new_n854));
  NOR2_X1   g493(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OR2_X1    g494(.A1(new_n477), .A2(new_n429), .ZN(new_n856));
  NAND2_X1  g495(.A1(new_n437), .A2(G86), .ZN(new_n857));
  NAND4_X1  g496(.A1(new_n856), .A2(new_n646), .A3(new_n857), .A4(new_n479), .ZN(new_n858));
  OAI21_X1  g497(.A(G1981), .B1(new_n478), .B2(new_n481), .ZN(new_n859));
  NAND2_X1  g498(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g499(.A(KEYINPUT49), .ZN(new_n861));
  NAND2_X1  g500(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g501(.A1(new_n858), .A2(KEYINPUT49), .A3(new_n859), .ZN(new_n863));
  AND3_X1   g502(.A1(new_n862), .A2(new_n847), .A3(new_n863), .ZN(new_n864));
  NOR2_X1   g503(.A1(new_n855), .A2(new_n864), .ZN(new_n865));
  OAI211_X1 g504(.A(new_n843), .B(G8), .C1(new_n838), .C2(new_n839), .ZN(new_n866));
  NAND3_X1  g505(.A1(new_n845), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NOR2_X1   g506(.A1(new_n837), .A2(new_n867), .ZN(new_n868));
  INV_X1    g507(.A(KEYINPUT54), .ZN(new_n869));
  NAND2_X1  g508(.A1(new_n701), .A2(new_n791), .ZN(new_n870));
  AOI21_X1  g509(.A(new_n789), .B1(new_n870), .B2(KEYINPUT50), .ZN(new_n871));
  NAND2_X1  g510(.A1(new_n871), .A2(new_n827), .ZN(new_n872));
  INV_X1    g511(.A(G1961), .ZN(new_n873));
  NAND2_X1  g512(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g513(.A(KEYINPUT53), .ZN(new_n875));
  NAND3_X1  g514(.A1(new_n794), .A2(new_n875), .A3(new_n601), .ZN(new_n876));
  INV_X1    g515(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g516(.A(new_n875), .B1(new_n794), .B2(new_n601), .ZN(new_n878));
  OAI21_X1  g517(.A(new_n874), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g518(.A1(new_n879), .A2(G171), .ZN(new_n880));
  OAI21_X1  g519(.A(new_n771), .B1(new_n806), .B2(new_n807), .ZN(new_n881));
  OAI21_X1  g520(.A(KEYINPUT53), .B1(new_n881), .B2(G2078), .ZN(new_n882));
  AOI22_X1  g521(.A1(new_n882), .A2(new_n876), .B1(new_n873), .B2(new_n872), .ZN(new_n883));
  NOR2_X1   g522(.A1(new_n883), .A2(G301), .ZN(new_n884));
  OAI21_X1  g523(.A(new_n869), .B1(new_n880), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g524(.A1(new_n879), .A2(G171), .ZN(new_n886));
  NAND2_X1  g525(.A1(new_n883), .A2(G301), .ZN(new_n887));
  NAND3_X1  g526(.A1(new_n886), .A2(new_n887), .A3(KEYINPUT54), .ZN(new_n888));
  NAND4_X1  g527(.A1(new_n826), .A2(new_n868), .A3(new_n885), .A4(new_n888), .ZN(new_n889));
  NOR2_X1   g528(.A1(new_n867), .A2(new_n886), .ZN(new_n890));
  INV_X1    g529(.A(KEYINPUT62), .ZN(new_n891));
  AOI211_X1 g530(.A(new_n891), .B(new_n831), .C1(new_n835), .C2(new_n836), .ZN(new_n892));
  NAND2_X1  g531(.A1(new_n835), .A2(new_n836), .ZN(new_n893));
  INV_X1    g532(.A(new_n831), .ZN(new_n894));
  AOI21_X1  g533(.A(KEYINPUT62), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g534(.A(new_n890), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g535(.A1(new_n862), .A2(new_n847), .A3(new_n863), .ZN(new_n897));
  OAI21_X1  g536(.A(new_n897), .B1(new_n854), .B2(new_n853), .ZN(new_n898));
  NOR2_X1   g537(.A1(G288), .A2(G1976), .ZN(new_n899));
  AOI22_X1  g538(.A1(new_n897), .A2(new_n899), .B1(new_n646), .B2(new_n482), .ZN(new_n900));
  INV_X1    g539(.A(new_n847), .ZN(new_n901));
  OAI22_X1  g540(.A1(new_n866), .A2(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g541(.A1(new_n832), .A2(G286), .ZN(new_n903));
  NAND4_X1  g542(.A1(new_n845), .A2(new_n903), .A3(new_n865), .A4(new_n866), .ZN(new_n904));
  INV_X1    g543(.A(KEYINPUT63), .ZN(new_n905));
  NAND2_X1  g544(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g545(.A(new_n839), .ZN(new_n907));
  NAND2_X1  g546(.A1(new_n881), .A2(new_n653), .ZN(new_n908));
  AOI21_X1  g547(.A(new_n846), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g548(.A(new_n898), .B1(new_n909), .B2(new_n843), .ZN(new_n910));
  NAND4_X1  g549(.A1(new_n910), .A2(KEYINPUT63), .A3(new_n845), .A4(new_n903), .ZN(new_n911));
  AOI21_X1  g550(.A(new_n902), .B1(new_n906), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g551(.A1(new_n889), .A2(new_n896), .A3(new_n912), .ZN(new_n913));
  NOR3_X1   g552(.A1(new_n806), .A2(new_n807), .A3(new_n789), .ZN(new_n914));
  NAND3_X1  g553(.A1(new_n914), .A2(new_n668), .A3(new_n777), .ZN(new_n915));
  NAND3_X1  g554(.A1(new_n914), .A2(G290), .A3(new_n777), .ZN(new_n916));
  XNOR2_X1  g555(.A(new_n915), .B(new_n916), .ZN(new_n917));
  INV_X1    g556(.A(new_n914), .ZN(new_n918));
  NOR4_X1   g557(.A1(new_n918), .A2(new_n662), .A3(new_n664), .A4(new_n778), .ZN(new_n919));
  AND4_X1   g558(.A1(new_n662), .A2(new_n914), .A3(new_n664), .A4(new_n777), .ZN(new_n920));
  NOR2_X1   g559(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g560(.A1(new_n914), .A2(new_n618), .A3(new_n777), .ZN(new_n922));
  NAND3_X1  g561(.A1(new_n914), .A2(new_n620), .A3(new_n777), .ZN(new_n923));
  XNOR2_X1  g562(.A(new_n922), .B(new_n923), .ZN(new_n924));
  NAND3_X1  g563(.A1(new_n914), .A2(new_n636), .A3(new_n777), .ZN(new_n925));
  NAND3_X1  g564(.A1(new_n914), .A2(new_n638), .A3(new_n777), .ZN(new_n926));
  XNOR2_X1  g565(.A(new_n925), .B(new_n926), .ZN(new_n927));
  AND4_X1   g566(.A1(new_n917), .A2(new_n921), .A3(new_n924), .A4(new_n927), .ZN(new_n928));
  NAND2_X1  g567(.A1(new_n913), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g568(.A1(new_n927), .A2(new_n924), .A3(new_n919), .ZN(new_n930));
  NAND3_X1  g569(.A1(new_n924), .A2(new_n927), .A3(new_n921), .ZN(new_n931));
  NOR2_X1   g570(.A1(new_n915), .A2(G290), .ZN(new_n932));
  XNOR2_X1  g571(.A(new_n932), .B(KEYINPUT48), .ZN(new_n933));
  OAI221_X1 g572(.A(new_n930), .B1(new_n618), .B2(new_n923), .C1(new_n931), .C2(new_n933), .ZN(new_n934));
  XNOR2_X1  g573(.A(new_n926), .B(KEYINPUT46), .ZN(new_n935));
  NAND3_X1  g574(.A1(new_n924), .A2(new_n935), .A3(new_n925), .ZN(new_n936));
  NAND2_X1  g575(.A1(new_n936), .A2(KEYINPUT47), .ZN(new_n937));
  OR2_X1    g576(.A1(new_n936), .A2(KEYINPUT47), .ZN(new_n938));
  AOI21_X1  g577(.A(new_n934), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g578(.A1(new_n929), .A2(new_n939), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g579(.A1(G401), .A2(new_n395), .A3(G227), .A4(G229), .ZN(new_n942));
  OAI211_X1 g580(.A(new_n717), .B(new_n942), .C1(new_n756), .C2(new_n763), .ZN(G225));
  INV_X1    g581(.A(G225), .ZN(G308));
endmodule


