//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 1 1 0 1 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 0 1 0 0 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n801, new_n802, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n974, new_n975, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1031, new_n1032;
  INV_X1    g000(.A(G183gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT27), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT27), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G183gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT69), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT69), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n203), .A2(new_n205), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT28), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(G190gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n207), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT70), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AND2_X1   g013(.A1(new_n207), .A2(new_n209), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n215), .A2(KEYINPUT70), .A3(new_n211), .ZN(new_n216));
  INV_X1    g015(.A(G190gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n204), .A2(G183gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT67), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(KEYINPUT67), .B1(new_n203), .B2(new_n205), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n210), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n222), .A2(KEYINPUT68), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT68), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n224), .B(new_n210), .C1(new_n220), .C2(new_n221), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n214), .B(new_n216), .C1(new_n223), .C2(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n202), .A2(new_n217), .ZN(new_n228));
  NAND2_X1  g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(G169gat), .A2(G176gat), .ZN(new_n231));
  NOR3_X1   g030(.A1(new_n230), .A2(new_n231), .A3(KEYINPUT26), .ZN(new_n232));
  AOI211_X1 g031(.A(new_n228), .B(new_n232), .C1(KEYINPUT26), .C2(new_n231), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n227), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n231), .A2(KEYINPUT23), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT23), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n236), .B1(G169gat), .B2(G176gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n235), .A2(new_n229), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT24), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n239), .A2(G183gat), .A3(G190gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(G183gat), .B(G190gat), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n240), .B1(new_n241), .B2(new_n239), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT64), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n238), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  OAI211_X1 g043(.A(KEYINPUT64), .B(new_n240), .C1(new_n241), .C2(new_n239), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT25), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n242), .A2(KEYINPUT65), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n250), .B(new_n240), .C1(new_n241), .C2(new_n239), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  AND3_X1   g051(.A1(new_n235), .A2(new_n229), .A3(new_n237), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n252), .A2(KEYINPUT25), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT66), .B1(new_n248), .B2(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT25), .B1(new_n244), .B2(new_n245), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n253), .A2(KEYINPUT25), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n257), .B1(new_n249), .B2(new_n251), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n259));
  NOR3_X1   g058(.A1(new_n256), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n234), .B1(new_n255), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(G113gat), .ZN(new_n262));
  INV_X1    g061(.A(G120gat), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT1), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G127gat), .B(G134gat), .ZN(new_n265));
  XOR2_X1   g064(.A(KEYINPUT71), .B(G120gat), .Z(new_n266));
  OAI211_X1 g065(.A(new_n264), .B(new_n265), .C1(new_n266), .C2(new_n262), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n264), .B1(new_n262), .B2(new_n263), .ZN(new_n268));
  INV_X1    g067(.A(new_n265), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n261), .A2(new_n272), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n234), .B(new_n271), .C1(new_n255), .C2(new_n260), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G227gat), .ZN(new_n276));
  INV_X1    g075(.A(G233gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  AND2_X1   g079(.A1(new_n280), .A2(KEYINPUT34), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(KEYINPUT34), .ZN(new_n282));
  OR2_X1    g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT32), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n273), .A2(new_n278), .A3(new_n274), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT72), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n273), .A2(KEYINPUT72), .A3(new_n278), .A4(new_n274), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n284), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT33), .B1(new_n287), .B2(new_n288), .ZN(new_n290));
  XOR2_X1   g089(.A(G15gat), .B(G43gat), .Z(new_n291));
  XNOR2_X1  g090(.A(G71gat), .B(G99gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NOR3_X1   g093(.A1(new_n289), .A2(new_n290), .A3(new_n294), .ZN(new_n295));
  AOI221_X4 g094(.A(new_n284), .B1(KEYINPUT33), .B2(new_n293), .C1(new_n287), .C2(new_n288), .ZN(new_n296));
  NOR3_X1   g095(.A1(new_n295), .A2(KEYINPUT73), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT73), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n287), .A2(new_n288), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT32), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT33), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n300), .A2(new_n302), .A3(new_n293), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n289), .B1(new_n290), .B2(new_n294), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n298), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n283), .B1(new_n297), .B2(new_n305), .ZN(new_n306));
  NOR3_X1   g105(.A1(new_n295), .A2(new_n283), .A3(new_n296), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT36), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT74), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n283), .B1(new_n295), .B2(new_n296), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n281), .A2(new_n282), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n303), .A2(new_n313), .A3(new_n304), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n311), .B1(new_n315), .B2(new_n308), .ZN(new_n316));
  AOI211_X1 g115(.A(KEYINPUT74), .B(KEYINPUT36), .C1(new_n312), .C2(new_n314), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n310), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G1gat), .B(G29gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n319), .B(KEYINPUT0), .ZN(new_n320));
  XNOR2_X1  g119(.A(G57gat), .B(G85gat), .ZN(new_n321));
  XOR2_X1   g120(.A(new_n320), .B(new_n321), .Z(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT2), .ZN(new_n324));
  INV_X1    g123(.A(G141gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n325), .A2(G148gat), .ZN(new_n326));
  INV_X1    g125(.A(G148gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n327), .A2(G141gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n324), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G155gat), .A2(G162gat), .ZN(new_n330));
  INV_X1    g129(.A(G155gat), .ZN(new_n331));
  INV_X1    g130(.A(G162gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n329), .A2(new_n330), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT76), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n335), .B1(new_n325), .B2(G148gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n327), .A2(KEYINPUT76), .A3(G141gat), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n336), .B(new_n337), .C1(G141gat), .C2(new_n327), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n330), .B1(new_n333), .B2(KEYINPUT2), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n334), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n271), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n334), .A2(new_n340), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n344), .A2(KEYINPUT3), .ZN(new_n345));
  OR2_X1    g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G225gat), .A2(G233gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT4), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n272), .A2(new_n349), .A3(new_n341), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT4), .B1(new_n271), .B2(new_n344), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NOR3_X1   g153(.A1(new_n348), .A2(new_n354), .A3(KEYINPUT5), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT5), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n271), .B(new_n344), .ZN(new_n357));
  INV_X1    g156(.A(new_n347), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n350), .A2(KEYINPUT77), .A3(new_n352), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT77), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n361), .B(KEYINPUT4), .C1(new_n271), .C2(new_n344), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n362), .B(new_n347), .C1(new_n343), .C2(new_n345), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n359), .B1(new_n360), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT78), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT78), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n359), .B(new_n366), .C1(new_n360), .C2(new_n363), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n355), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n323), .B1(new_n368), .B2(KEYINPUT83), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(KEYINPUT83), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT82), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n346), .B1(new_n353), .B2(new_n351), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(new_n358), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n322), .B1(new_n374), .B2(KEYINPUT39), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT39), .B1(new_n357), .B2(new_n358), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n376), .B1(new_n373), .B2(new_n358), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n372), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT40), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n372), .B(KEYINPUT40), .C1(new_n375), .C2(new_n377), .ZN(new_n381));
  AOI22_X1  g180(.A1(new_n370), .A2(new_n371), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n248), .A2(new_n254), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n234), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G226gat), .A2(G233gat), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n387), .A2(KEYINPUT29), .ZN(new_n388));
  AOI22_X1  g187(.A1(new_n385), .A2(new_n387), .B1(new_n261), .B2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G197gat), .B(G204gat), .ZN(new_n390));
  INV_X1    g189(.A(G211gat), .ZN(new_n391));
  INV_X1    g190(.A(G218gat), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n390), .B1(KEYINPUT22), .B2(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(G211gat), .B(G218gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n389), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n261), .ZN(new_n399));
  AOI22_X1  g198(.A1(new_n399), .A2(new_n387), .B1(new_n388), .B2(new_n384), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n400), .A2(new_n396), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT75), .B1(new_n398), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT75), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n397), .B(new_n403), .C1(new_n396), .C2(new_n400), .ZN(new_n404));
  XNOR2_X1  g203(.A(G8gat), .B(G36gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(G64gat), .B(G92gat), .ZN(new_n406));
  XOR2_X1   g205(.A(new_n405), .B(new_n406), .Z(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n402), .A2(new_n404), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n397), .B(new_n407), .C1(new_n396), .C2(new_n400), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT30), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n382), .B1(new_n410), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT80), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n368), .A2(new_n322), .ZN(new_n416));
  XNOR2_X1  g215(.A(KEYINPUT79), .B(KEYINPUT6), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n415), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NOR4_X1   g218(.A1(new_n368), .A2(KEYINPUT80), .A3(new_n322), .A4(new_n417), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n384), .A2(new_n388), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n422), .B(new_n396), .C1(new_n386), .C2(new_n261), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n423), .B(KEYINPUT84), .C1(new_n389), .C2(new_n396), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n424), .B(KEYINPUT37), .C1(KEYINPUT84), .C2(new_n423), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT38), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT37), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n397), .B(new_n427), .C1(new_n396), .C2(new_n400), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n425), .A2(new_n426), .A3(new_n408), .A4(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n418), .B1(new_n368), .B2(new_n322), .ZN(new_n430));
  INV_X1    g229(.A(new_n371), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n430), .B1(new_n431), .B2(new_n369), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n421), .A2(new_n429), .A3(new_n411), .A4(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n402), .A2(KEYINPUT37), .A3(new_n404), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n428), .A2(new_n408), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n426), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n414), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT81), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n342), .B1(new_n396), .B2(KEYINPUT29), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n344), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n396), .B1(new_n345), .B2(KEYINPUT29), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(G228gat), .A2(G233gat), .ZN(new_n443));
  AND2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n442), .A2(new_n443), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n438), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(G78gat), .B(G106gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(KEYINPUT31), .B(G50gat), .ZN(new_n448));
  XOR2_X1   g247(.A(new_n447), .B(new_n448), .Z(new_n449));
  NAND2_X1  g248(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(G22gat), .ZN(new_n451));
  NOR3_X1   g250(.A1(new_n444), .A2(new_n445), .A3(new_n438), .ZN(new_n452));
  INV_X1    g251(.A(G22gat), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n446), .A2(new_n453), .A3(new_n449), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n451), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n452), .B1(new_n451), .B2(new_n454), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n437), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n411), .B(KEYINPUT30), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n409), .ZN(new_n460));
  INV_X1    g259(.A(new_n368), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n461), .A2(new_n323), .A3(new_n418), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT80), .ZN(new_n463));
  INV_X1    g262(.A(new_n420), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n430), .B1(new_n322), .B2(new_n368), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NOR3_X1   g265(.A1(new_n460), .A2(new_n466), .A3(new_n457), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n458), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n460), .A2(new_n466), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n314), .A2(new_n457), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n306), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT35), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n463), .A2(new_n464), .ZN(new_n475));
  INV_X1    g274(.A(new_n432), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT35), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n457), .A2(new_n478), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n477), .A2(new_n479), .A3(new_n460), .ZN(new_n480));
  INV_X1    g279(.A(new_n315), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n318), .A2(new_n469), .B1(new_n474), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(G50gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(G43gat), .ZN(new_n485));
  INV_X1    g284(.A(G43gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(G50gat), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n485), .A2(new_n487), .A3(KEYINPUT15), .ZN(new_n488));
  INV_X1    g287(.A(G29gat), .ZN(new_n489));
  INV_X1    g288(.A(G36gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT85), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT85), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(G36gat), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n489), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n489), .A2(new_n490), .A3(KEYINPUT14), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT14), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n496), .B1(G29gat), .B2(G36gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NOR3_X1   g297(.A1(new_n488), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(G43gat), .B(G50gat), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT86), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT15), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n486), .A2(KEYINPUT86), .A3(G50gat), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n488), .B1(new_n494), .B2(new_n498), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n499), .A2(new_n505), .B1(new_n506), .B2(KEYINPUT87), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n495), .A2(new_n497), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n492), .A2(G36gat), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n490), .A2(KEYINPUT85), .ZN(new_n510));
  OAI21_X1  g309(.A(G29gat), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n485), .A2(new_n487), .A3(KEYINPUT15), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n508), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n504), .A2(new_n503), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n514), .B1(new_n501), .B2(new_n500), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT87), .ZN(new_n516));
  NOR3_X1   g315(.A1(new_n513), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT88), .B1(new_n507), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT17), .ZN(new_n519));
  XNOR2_X1  g318(.A(G15gat), .B(G22gat), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n520), .A2(G1gat), .ZN(new_n521));
  INV_X1    g320(.A(G1gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT16), .ZN(new_n523));
  INV_X1    g322(.A(G15gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(G22gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n453), .A2(G15gat), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(G8gat), .B1(new_n521), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n520), .A2(new_n523), .ZN(new_n529));
  INV_X1    g328(.A(G8gat), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n529), .B(new_n530), .C1(G1gat), .C2(new_n520), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n499), .A2(KEYINPUT87), .A3(new_n505), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n513), .A2(new_n515), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n508), .A2(new_n511), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n516), .B1(new_n535), .B2(new_n488), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n533), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT17), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n537), .A2(KEYINPUT88), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n519), .A2(new_n532), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G229gat), .A2(G233gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n506), .A2(KEYINPUT87), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n542), .B1(new_n515), .B2(new_n513), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n532), .B1(new_n543), .B2(new_n533), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n540), .A2(new_n541), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT18), .ZN(new_n547));
  XOR2_X1   g346(.A(new_n541), .B(KEYINPUT13), .Z(new_n548));
  AND3_X1   g347(.A1(new_n543), .A2(new_n532), .A3(new_n533), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n548), .B1(new_n549), .B2(new_n544), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT90), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT90), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n552), .B(new_n548), .C1(new_n549), .C2(new_n544), .ZN(new_n553));
  AOI22_X1  g352(.A1(new_n546), .A2(new_n547), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n540), .A2(KEYINPUT18), .A3(new_n541), .A4(new_n545), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT89), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n555), .A2(new_n556), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n554), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G113gat), .B(G141gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(G197gat), .ZN(new_n561));
  XOR2_X1   g360(.A(KEYINPUT11), .B(G169gat), .Z(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(KEYINPUT12), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n546), .A2(new_n547), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n553), .ZN(new_n567));
  AND3_X1   g366(.A1(new_n566), .A2(new_n567), .A3(new_n564), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n555), .B(new_n556), .ZN(new_n569));
  AOI22_X1  g368(.A1(new_n559), .A2(new_n565), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n483), .A2(new_n570), .ZN(new_n571));
  AND2_X1   g370(.A1(G232gat), .A2(G233gat), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n572), .A2(KEYINPUT41), .ZN(new_n573));
  XNOR2_X1  g372(.A(G134gat), .B(G162gat), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n573), .B(new_n574), .Z(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(G85gat), .A2(G92gat), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT7), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(G99gat), .A2(G106gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(KEYINPUT8), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT95), .ZN(new_n585));
  OR2_X1    g384(.A1(G85gat), .A2(G92gat), .ZN(new_n586));
  AND3_X1   g385(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n585), .B1(new_n584), .B2(new_n586), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n582), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  XOR2_X1   g388(.A(G99gat), .B(G106gat), .Z(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT8), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n592), .B1(G99gat), .B2(G106gat), .ZN(new_n593));
  NOR2_X1   g392(.A1(G85gat), .A2(G92gat), .ZN(new_n594));
  OAI21_X1  g393(.A(KEYINPUT95), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n584), .A2(new_n586), .A3(new_n585), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n590), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n597), .A2(new_n598), .A3(new_n582), .ZN(new_n599));
  AND3_X1   g398(.A1(new_n591), .A2(new_n599), .A3(KEYINPUT96), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT96), .B1(new_n591), .B2(new_n599), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n519), .A2(new_n602), .A3(new_n539), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT96), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n598), .B1(new_n597), .B2(new_n582), .ZN(new_n605));
  AOI211_X1 g404(.A(new_n590), .B(new_n581), .C1(new_n595), .C2(new_n596), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n591), .A2(new_n599), .A3(KEYINPUT96), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI22_X1  g408(.A1(new_n609), .A2(new_n537), .B1(KEYINPUT41), .B2(new_n572), .ZN(new_n610));
  AND3_X1   g409(.A1(new_n603), .A2(new_n610), .A3(KEYINPUT97), .ZN(new_n611));
  AOI21_X1  g410(.A(KEYINPUT97), .B1(new_n603), .B2(new_n610), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n217), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n603), .A2(new_n610), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT97), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n603), .A2(new_n610), .A3(KEYINPUT97), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n616), .A2(G190gat), .A3(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n613), .A2(new_n618), .A3(G218gat), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT94), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(G218gat), .B1(new_n613), .B2(new_n618), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n576), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G127gat), .B(G155gat), .ZN(new_n624));
  AND2_X1   g423(.A1(G71gat), .A2(G78gat), .ZN(new_n625));
  NOR2_X1   g424(.A1(G71gat), .A2(G78gat), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G57gat), .B(G64gat), .ZN(new_n628));
  AOI21_X1  g427(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(G57gat), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(G64gat), .ZN(new_n632));
  INV_X1    g431(.A(G64gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(G57gat), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G71gat), .B(G78gat), .ZN(new_n636));
  INV_X1    g435(.A(new_n629), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  AND3_X1   g437(.A1(new_n630), .A2(new_n638), .A3(KEYINPUT91), .ZN(new_n639));
  AOI21_X1  g438(.A(KEYINPUT91), .B1(new_n630), .B2(new_n638), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT21), .ZN(new_n642));
  INV_X1    g441(.A(G231gat), .ZN(new_n643));
  OAI211_X1 g442(.A(new_n641), .B(new_n642), .C1(new_n643), .C2(new_n277), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n643), .A2(new_n277), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n638), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT91), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n630), .A2(new_n638), .A3(KEYINPUT91), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n645), .B1(new_n650), .B2(KEYINPUT21), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n644), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n652), .B1(new_n644), .B2(new_n651), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n624), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n655), .ZN(new_n657));
  INV_X1    g456(.A(new_n624), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n657), .A2(new_n653), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g458(.A(G183gat), .B(G211gat), .Z(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  AND3_X1   g460(.A1(new_n656), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n661), .B1(new_n656), .B2(new_n659), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n532), .B1(new_n641), .B2(new_n642), .ZN(new_n664));
  XOR2_X1   g463(.A(KEYINPUT92), .B(KEYINPUT93), .Z(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  OR3_X1    g466(.A1(new_n662), .A2(new_n663), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n667), .B1(new_n662), .B2(new_n663), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n613), .A2(new_n618), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n392), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n672), .A2(new_n620), .A3(new_n619), .A4(new_n575), .ZN(new_n673));
  XNOR2_X1  g472(.A(G120gat), .B(G148gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(G176gat), .B(G204gat), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n674), .B(new_n675), .Z(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  OAI22_X1  g476(.A1(new_n605), .A2(new_n606), .B1(new_n639), .B2(new_n640), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n591), .A2(new_n599), .A3(new_n646), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  AND2_X1   g480(.A1(G230gat), .A2(G233gat), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n677), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT10), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n641), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n609), .A2(new_n685), .ZN(new_n686));
  AOI22_X1  g485(.A1(new_n599), .A2(new_n591), .B1(new_n648), .B2(new_n649), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n591), .A2(new_n599), .A3(new_n646), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n684), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(KEYINPUT98), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT98), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n680), .A2(new_n691), .A3(new_n684), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n686), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n683), .B1(new_n693), .B2(new_n682), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n609), .A2(new_n685), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n691), .B1(new_n680), .B2(new_n684), .ZN(new_n696));
  AOI211_X1 g495(.A(KEYINPUT98), .B(KEYINPUT10), .C1(new_n678), .C2(new_n679), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n695), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  XOR2_X1   g497(.A(new_n682), .B(KEYINPUT99), .Z(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  AOI22_X1  g499(.A1(new_n698), .A2(new_n700), .B1(new_n682), .B2(new_n681), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n694), .B1(new_n701), .B2(new_n676), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n623), .A2(new_n670), .A3(new_n673), .A4(new_n703), .ZN(new_n704));
  XOR2_X1   g503(.A(new_n704), .B(KEYINPUT100), .Z(new_n705));
  INV_X1    g504(.A(new_n466), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n706), .A2(KEYINPUT101), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(KEYINPUT101), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n571), .A2(new_n705), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g510(.A(KEYINPUT16), .B(G8gat), .Z(new_n712));
  NAND4_X1  g511(.A1(new_n571), .A2(new_n460), .A3(new_n705), .A4(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n571), .A2(new_n705), .ZN(new_n714));
  INV_X1    g513(.A(new_n460), .ZN(new_n715));
  OAI21_X1  g514(.A(G8gat), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n713), .ZN(new_n717));
  MUX2_X1   g516(.A(new_n713), .B(new_n717), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g517(.A(G15gat), .B1(new_n714), .B2(new_n318), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n571), .A2(new_n524), .A3(new_n481), .A4(new_n705), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(G1326gat));
  NOR2_X1   g520(.A1(new_n714), .A2(new_n457), .ZN(new_n722));
  XOR2_X1   g521(.A(KEYINPUT43), .B(G22gat), .Z(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1327gat));
  NAND2_X1  g523(.A1(new_n623), .A2(new_n673), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n726), .A2(new_n670), .A3(new_n702), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n571), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n728), .A2(new_n489), .A3(new_n709), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT45), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(new_n483), .B2(new_n726), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n313), .B1(new_n303), .B2(new_n304), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n308), .B1(new_n307), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(KEYINPUT74), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n315), .A2(new_n311), .A3(new_n308), .ZN(new_n736));
  AOI22_X1  g535(.A1(new_n735), .A2(new_n736), .B1(new_n306), .B2(new_n309), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n467), .B1(new_n437), .B2(new_n457), .ZN(new_n738));
  OAI21_X1  g537(.A(KEYINPUT73), .B1(new_n295), .B2(new_n296), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n303), .A2(new_n298), .A3(new_n304), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n471), .B1(new_n741), .B2(new_n283), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n478), .B1(new_n742), .B2(new_n470), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n480), .A2(new_n481), .ZN(new_n744));
  OAI22_X1  g543(.A1(new_n737), .A2(new_n738), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n745), .A2(KEYINPUT44), .A3(new_n725), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n732), .A2(new_n746), .ZN(new_n747));
  XOR2_X1   g546(.A(new_n670), .B(KEYINPUT102), .Z(new_n748));
  NOR3_X1   g547(.A1(new_n748), .A2(new_n570), .A3(new_n702), .ZN(new_n749));
  AND3_X1   g548(.A1(new_n747), .A2(new_n709), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n730), .B1(new_n489), .B2(new_n750), .ZN(G1328gat));
  XNOR2_X1  g550(.A(KEYINPUT85), .B(G36gat), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n460), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n571), .A2(new_n727), .A3(new_n753), .ZN(new_n754));
  OR2_X1    g553(.A1(new_n754), .A2(KEYINPUT103), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(KEYINPUT103), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT46), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n755), .A2(KEYINPUT46), .A3(new_n756), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n747), .A2(new_n460), .A3(new_n749), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n759), .B(new_n760), .C1(new_n752), .C2(new_n761), .ZN(G1329gat));
  NAND3_X1  g561(.A1(new_n728), .A2(new_n486), .A3(new_n481), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n732), .A2(new_n746), .A3(new_n737), .A4(new_n749), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(G43gat), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT47), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n766), .B(new_n767), .ZN(G1330gat));
  INV_X1    g567(.A(new_n457), .ZN(new_n769));
  AND4_X1   g568(.A1(new_n484), .A2(new_n571), .A3(new_n769), .A4(new_n727), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n732), .A2(new_n746), .A3(new_n769), .A4(new_n749), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G50gat), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n771), .A2(new_n773), .A3(KEYINPUT48), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT105), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n772), .A2(new_n775), .A3(G50gat), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n775), .B1(new_n772), .B2(G50gat), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n776), .A2(new_n777), .A3(new_n770), .ZN(new_n778));
  XOR2_X1   g577(.A(KEYINPUT104), .B(KEYINPUT48), .Z(new_n779));
  OAI21_X1  g578(.A(new_n774), .B1(new_n778), .B2(new_n779), .ZN(G1331gat));
  NAND4_X1  g579(.A1(new_n726), .A2(new_n570), .A3(new_n670), .A4(new_n702), .ZN(new_n781));
  OR3_X1    g580(.A1(new_n483), .A2(KEYINPUT106), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(KEYINPUT106), .B1(new_n483), .B2(new_n781), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n707), .A2(new_n708), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(new_n631), .ZN(G1332gat));
  NOR2_X1   g586(.A1(new_n784), .A2(new_n715), .ZN(new_n788));
  NOR2_X1   g587(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n789));
  AND2_X1   g588(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n791), .B1(new_n788), .B2(new_n789), .ZN(G1333gat));
  OAI21_X1  g591(.A(G71gat), .B1(new_n784), .B2(new_n318), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n315), .A2(G71gat), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n782), .A2(new_n783), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT50), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n793), .A2(KEYINPUT50), .A3(new_n795), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(G1334gat));
  NOR2_X1   g599(.A1(new_n784), .A2(new_n457), .ZN(new_n801));
  XNOR2_X1  g600(.A(KEYINPUT107), .B(G78gat), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n801), .B(new_n802), .ZN(G1335gat));
  NAND2_X1  g602(.A1(new_n559), .A2(new_n565), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n554), .B(new_n564), .C1(new_n557), .C2(new_n558), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n670), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT108), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n745), .A2(new_n725), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n745), .A2(KEYINPUT51), .A3(new_n725), .A4(new_n808), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n785), .A2(G85gat), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n813), .A2(new_n702), .A3(new_n814), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n808), .A2(new_n702), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n747), .A2(new_n709), .A3(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT109), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(G85gat), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n817), .A2(new_n818), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n815), .B1(new_n820), .B2(new_n821), .ZN(G1336gat));
  NAND4_X1  g621(.A1(new_n732), .A2(new_n746), .A3(new_n460), .A4(new_n816), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(G92gat), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n715), .A2(G92gat), .A3(new_n703), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT110), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n826), .B1(new_n811), .B2(new_n812), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n824), .B1(new_n827), .B2(KEYINPUT111), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT111), .ZN(new_n829));
  AOI211_X1 g628(.A(new_n829), .B(new_n826), .C1(new_n811), .C2(new_n812), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT52), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(KEYINPUT52), .B1(new_n813), .B2(new_n825), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n824), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(G1337gat));
  NAND3_X1  g633(.A1(new_n747), .A2(new_n737), .A3(new_n816), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(G99gat), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n315), .A2(G99gat), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n813), .A2(new_n702), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(G1338gat));
  NOR2_X1   g638(.A1(new_n457), .A2(G106gat), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n813), .A2(new_n702), .A3(new_n840), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n732), .A2(new_n746), .A3(new_n769), .A4(new_n816), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(G106gat), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(KEYINPUT53), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n841), .A2(new_n846), .A3(new_n843), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(new_n847), .ZN(G1339gat));
  NOR2_X1   g647(.A1(new_n704), .A2(new_n806), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n699), .B(new_n695), .C1(new_n696), .C2(new_n697), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n851), .B(KEYINPUT54), .C1(new_n693), .C2(new_n682), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n698), .A2(new_n853), .A3(new_n700), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n852), .A2(KEYINPUT55), .A3(new_n677), .A4(new_n854), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n855), .A2(new_n694), .ZN(new_n856));
  OR3_X1    g655(.A1(new_n549), .A2(new_n544), .A3(new_n548), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n541), .B1(new_n540), .B2(new_n545), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT112), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AOI211_X1 g659(.A(KEYINPUT112), .B(new_n541), .C1(new_n540), .C2(new_n545), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n563), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n805), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n852), .A2(new_n677), .A3(new_n854), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT55), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AND3_X1   g665(.A1(new_n856), .A2(new_n863), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n725), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n805), .A2(new_n702), .A3(new_n862), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT113), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n805), .A2(new_n702), .A3(new_n862), .A4(KEYINPUT113), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n806), .A2(new_n856), .A3(new_n866), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT114), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n725), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n874), .A2(new_n875), .A3(KEYINPUT114), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n869), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n850), .B1(new_n880), .B2(new_n748), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n315), .A2(new_n769), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n785), .A2(new_n460), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(G113gat), .B1(new_n885), .B2(new_n570), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT115), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n881), .A2(new_n709), .ZN(new_n888));
  INV_X1    g687(.A(new_n742), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n888), .A2(new_n460), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n890), .A2(new_n262), .A3(new_n806), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n887), .A2(new_n891), .ZN(G1340gat));
  NAND3_X1  g691(.A1(new_n890), .A2(new_n266), .A3(new_n702), .ZN(new_n893));
  OAI21_X1  g692(.A(G120gat), .B1(new_n885), .B2(new_n703), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT116), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n894), .A2(new_n895), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n893), .B1(new_n896), .B2(new_n897), .ZN(G1341gat));
  INV_X1    g697(.A(G127gat), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n890), .A2(new_n899), .A3(new_n670), .ZN(new_n900));
  AND3_X1   g699(.A1(new_n883), .A2(new_n748), .A3(new_n884), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n900), .B1(new_n899), .B2(new_n901), .ZN(G1342gat));
  INV_X1    g701(.A(G134gat), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n890), .A2(new_n903), .A3(new_n725), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n904), .A2(KEYINPUT56), .ZN(new_n905));
  OAI21_X1  g704(.A(G134gat), .B1(new_n885), .B2(new_n726), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(KEYINPUT56), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(G1343gat));
  NAND2_X1  g707(.A1(new_n888), .A2(KEYINPUT121), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n881), .A2(new_n910), .A3(new_n709), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n318), .A2(new_n769), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n912), .A2(new_n460), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n909), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n806), .A2(new_n325), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n737), .A2(new_n460), .A3(new_n785), .ZN(new_n917));
  XOR2_X1   g716(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n919), .B1(new_n881), .B2(new_n769), .ZN(new_n920));
  INV_X1    g719(.A(new_n870), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT118), .ZN(new_n922));
  AND3_X1   g721(.A1(new_n864), .A2(new_n922), .A3(new_n865), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n922), .B1(new_n864), .B2(new_n865), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n855), .A2(new_n694), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n570), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n921), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n868), .B1(new_n928), .B2(new_n725), .ZN(new_n929));
  INV_X1    g728(.A(new_n670), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n849), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT57), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n457), .A2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(KEYINPUT119), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT119), .ZN(new_n936));
  INV_X1    g735(.A(new_n924), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n864), .A2(new_n922), .A3(new_n865), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n806), .A2(new_n856), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n870), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(new_n726), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n670), .B1(new_n942), .B2(new_n868), .ZN(new_n943));
  OAI211_X1 g742(.A(new_n936), .B(new_n933), .C1(new_n943), .C2(new_n849), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n935), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n917), .B1(new_n920), .B2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT120), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI211_X1 g747(.A(KEYINPUT120), .B(new_n917), .C1(new_n920), .C2(new_n945), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n948), .A2(new_n806), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n916), .B1(new_n950), .B2(G141gat), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT58), .ZN(new_n952));
  INV_X1    g751(.A(new_n946), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n325), .B1(new_n953), .B2(new_n806), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n952), .B1(new_n914), .B2(new_n915), .ZN(new_n955));
  OAI22_X1  g754(.A1(new_n951), .A2(new_n952), .B1(new_n954), .B2(new_n955), .ZN(G1344gat));
  INV_X1    g755(.A(KEYINPUT59), .ZN(new_n957));
  INV_X1    g756(.A(new_n914), .ZN(new_n958));
  AOI211_X1 g757(.A(new_n957), .B(G148gat), .C1(new_n958), .C2(new_n702), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n948), .A2(new_n702), .A3(new_n949), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(new_n957), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n881), .A2(new_n769), .A3(new_n919), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n705), .A2(new_n570), .ZN(new_n963));
  OR2_X1    g762(.A1(new_n963), .A2(KEYINPUT122), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n943), .B1(new_n963), .B2(KEYINPUT122), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n457), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n962), .B1(new_n966), .B2(KEYINPUT57), .ZN(new_n967));
  NAND4_X1  g766(.A1(new_n967), .A2(KEYINPUT59), .A3(new_n702), .A4(new_n917), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n961), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n959), .B1(new_n969), .B2(G148gat), .ZN(G1345gat));
  NAND3_X1  g769(.A1(new_n958), .A2(new_n331), .A3(new_n670), .ZN(new_n971));
  AND3_X1   g770(.A1(new_n948), .A2(new_n748), .A3(new_n949), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n971), .B1(new_n972), .B2(new_n331), .ZN(G1346gat));
  NAND4_X1  g772(.A1(new_n948), .A2(G162gat), .A3(new_n725), .A4(new_n949), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n332), .B1(new_n914), .B2(new_n726), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n974), .A2(new_n975), .ZN(G1347gat));
  AND2_X1   g775(.A1(new_n881), .A2(new_n785), .ZN(new_n977));
  AND3_X1   g776(.A1(new_n977), .A2(new_n460), .A3(new_n742), .ZN(new_n978));
  INV_X1    g777(.A(G169gat), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n978), .A2(new_n979), .A3(new_n806), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n709), .A2(new_n715), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n883), .A2(new_n806), .A3(new_n981), .ZN(new_n982));
  AND3_X1   g781(.A1(new_n982), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n983));
  AOI21_X1  g782(.A(KEYINPUT123), .B1(new_n982), .B2(G169gat), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n980), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(KEYINPUT124), .ZN(G1348gat));
  INV_X1    g785(.A(G176gat), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n978), .A2(new_n987), .A3(new_n702), .ZN(new_n988));
  AND2_X1   g787(.A1(new_n883), .A2(new_n981), .ZN(new_n989));
  AND2_X1   g788(.A1(new_n989), .A2(new_n702), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n988), .B1(new_n990), .B2(new_n987), .ZN(G1349gat));
  NAND4_X1  g790(.A1(new_n981), .A2(new_n881), .A3(new_n748), .A4(new_n882), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT125), .ZN(new_n993));
  OR2_X1    g792(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n202), .B1(new_n992), .B2(new_n993), .ZN(new_n995));
  AND2_X1   g794(.A1(new_n670), .A2(new_n215), .ZN(new_n996));
  AOI22_X1  g795(.A1(new_n994), .A2(new_n995), .B1(new_n978), .B2(new_n996), .ZN(new_n997));
  AND3_X1   g796(.A1(new_n997), .A2(KEYINPUT126), .A3(KEYINPUT60), .ZN(new_n998));
  NOR2_X1   g797(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n999));
  AND2_X1   g798(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n1000));
  NOR3_X1   g799(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  NOR2_X1   g800(.A1(new_n998), .A2(new_n1001), .ZN(G1350gat));
  AOI21_X1  g801(.A(new_n217), .B1(new_n989), .B2(new_n725), .ZN(new_n1003));
  INV_X1    g802(.A(KEYINPUT61), .ZN(new_n1004));
  XNOR2_X1  g803(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n978), .A2(new_n217), .A3(new_n725), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1005), .A2(new_n1006), .ZN(G1351gat));
  NOR3_X1   g806(.A1(new_n737), .A2(new_n709), .A3(new_n715), .ZN(new_n1008));
  INV_X1    g807(.A(new_n1008), .ZN(new_n1009));
  INV_X1    g808(.A(KEYINPUT127), .ZN(new_n1010));
  AOI21_X1  g809(.A(new_n1009), .B1(new_n967), .B2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g810(.A(KEYINPUT127), .B(new_n962), .C1(new_n966), .C2(KEYINPUT57), .ZN(new_n1012));
  NAND4_X1  g811(.A1(new_n1011), .A2(G197gat), .A3(new_n806), .A4(new_n1012), .ZN(new_n1013));
  INV_X1    g812(.A(G197gat), .ZN(new_n1014));
  NAND4_X1  g813(.A1(new_n977), .A2(new_n460), .A3(new_n769), .A4(new_n318), .ZN(new_n1015));
  OAI21_X1  g814(.A(new_n1014), .B1(new_n1015), .B2(new_n570), .ZN(new_n1016));
  AND2_X1   g815(.A1(new_n1013), .A2(new_n1016), .ZN(G1352gat));
  NAND2_X1  g816(.A1(new_n967), .A2(new_n1010), .ZN(new_n1018));
  NAND4_X1  g817(.A1(new_n1018), .A2(new_n702), .A3(new_n1012), .A4(new_n1008), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n1019), .A2(G204gat), .ZN(new_n1020));
  NOR3_X1   g819(.A1(new_n1015), .A2(G204gat), .A3(new_n703), .ZN(new_n1021));
  XNOR2_X1  g820(.A(new_n1021), .B(KEYINPUT62), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n1020), .A2(new_n1022), .ZN(G1353gat));
  NOR2_X1   g822(.A1(new_n1009), .A2(new_n930), .ZN(new_n1024));
  NAND2_X1  g823(.A1(new_n967), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g824(.A(KEYINPUT63), .B1(new_n1025), .B2(G211gat), .ZN(new_n1026));
  INV_X1    g825(.A(KEYINPUT63), .ZN(new_n1027));
  AOI211_X1 g826(.A(new_n1027), .B(new_n391), .C1(new_n967), .C2(new_n1024), .ZN(new_n1028));
  NAND2_X1  g827(.A1(new_n670), .A2(new_n391), .ZN(new_n1029));
  OAI22_X1  g828(.A1(new_n1026), .A2(new_n1028), .B1(new_n1015), .B2(new_n1029), .ZN(G1354gat));
  NAND4_X1  g829(.A1(new_n1011), .A2(G218gat), .A3(new_n725), .A4(new_n1012), .ZN(new_n1031));
  OAI21_X1  g830(.A(new_n392), .B1(new_n1015), .B2(new_n726), .ZN(new_n1032));
  AND2_X1   g831(.A1(new_n1031), .A2(new_n1032), .ZN(G1355gat));
endmodule


