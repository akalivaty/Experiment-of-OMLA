//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 0 1 0 1 0 0 1 0 1 1 1 1 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n187));
  INV_X1    g001(.A(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(G210), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT27), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n192), .B(KEYINPUT26), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G101), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT26), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n192), .B(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G101), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n194), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT28), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT64), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G143), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(new_n204), .A3(G146), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G143), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(KEYINPUT1), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n205), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n206), .A2(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n202), .A2(new_n204), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n211), .B1(new_n212), .B2(new_n206), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n208), .B1(new_n207), .B2(KEYINPUT1), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n210), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  XOR2_X1   g029(.A(KEYINPUT66), .B(G131), .Z(new_n216));
  INV_X1    g030(.A(KEYINPUT65), .ZN(new_n217));
  INV_X1    g031(.A(G137), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(KEYINPUT65), .A2(G137), .ZN(new_n220));
  AND2_X1   g034(.A1(KEYINPUT11), .A2(G134), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(KEYINPUT11), .A2(G134), .ZN(new_n223));
  NOR2_X1   g037(.A1(KEYINPUT11), .A2(G134), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n223), .B1(new_n224), .B2(G137), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n216), .A2(new_n222), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G134), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n219), .A2(new_n227), .A3(new_n220), .ZN(new_n228));
  INV_X1    g042(.A(G131), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n229), .B1(G134), .B2(G137), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n215), .A2(new_n226), .A3(new_n231), .ZN(new_n232));
  OR2_X1    g046(.A1(KEYINPUT2), .A2(G113), .ZN(new_n233));
  NAND2_X1  g047(.A1(KEYINPUT2), .A2(G113), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G116), .ZN(new_n236));
  INV_X1    g050(.A(G119), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(G116), .A2(G119), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n235), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n239), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(new_n233), .A3(new_n234), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n226), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n222), .A2(new_n225), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n229), .B1(new_n246), .B2(KEYINPUT67), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT67), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n222), .A2(new_n225), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n245), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  AND2_X1   g064(.A1(KEYINPUT0), .A2(G128), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n205), .A2(new_n207), .A3(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(KEYINPUT0), .A2(G128), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n252), .B1(new_n213), .B2(new_n255), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n232), .B(new_n244), .C1(new_n250), .C2(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n199), .B1(new_n200), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n246), .A2(KEYINPUT67), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(G131), .A3(new_n249), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n256), .B1(new_n261), .B2(new_n226), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n226), .A2(new_n231), .ZN(new_n263));
  INV_X1    g077(.A(new_n211), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT64), .B(G143), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n264), .B1(new_n265), .B2(G146), .ZN(new_n266));
  INV_X1    g080(.A(new_n214), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n263), .B1(new_n268), .B2(new_n210), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n243), .B1(new_n262), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n257), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT28), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT69), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n271), .A2(KEYINPUT69), .A3(KEYINPUT28), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n259), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT29), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT30), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n278), .B1(new_n262), .B2(new_n269), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n232), .B(KEYINPUT30), .C1(new_n250), .C2(new_n256), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n279), .A2(new_n243), .A3(new_n280), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n281), .A2(new_n257), .ZN(new_n282));
  INV_X1    g096(.A(new_n199), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n277), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n187), .B1(new_n276), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT69), .B1(new_n271), .B2(KEYINPUT28), .ZN(new_n286));
  AOI211_X1 g100(.A(new_n273), .B(new_n200), .C1(new_n270), .C2(new_n257), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n258), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n281), .A2(new_n257), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT29), .B1(new_n289), .B2(new_n199), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n288), .A2(KEYINPUT71), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n272), .A2(new_n258), .A3(KEYINPUT29), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT72), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT72), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n272), .A2(new_n258), .A3(new_n294), .A4(KEYINPUT29), .ZN(new_n295));
  AOI21_X1  g109(.A(G902), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n285), .A2(new_n291), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G472), .ZN(new_n298));
  INV_X1    g112(.A(G472), .ZN(new_n299));
  INV_X1    g113(.A(G902), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n257), .A2(new_n200), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n302), .B1(new_n286), .B2(new_n287), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n199), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT68), .ZN(new_n305));
  NOR3_X1   g119(.A1(new_n199), .A2(new_n305), .A3(KEYINPUT31), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n194), .A2(new_n198), .A3(KEYINPUT68), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n281), .A2(new_n257), .A3(new_n307), .ZN(new_n308));
  AOI22_X1  g122(.A1(new_n282), .A2(new_n306), .B1(new_n308), .B2(KEYINPUT31), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n301), .B1(new_n304), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(KEYINPUT70), .B1(new_n310), .B2(KEYINPUT32), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT70), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT32), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n308), .A2(KEYINPUT31), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n306), .A2(new_n257), .A3(new_n281), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n316), .B1(new_n303), .B2(new_n199), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n312), .B(new_n313), .C1(new_n317), .C2(new_n301), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n310), .A2(KEYINPUT32), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n298), .A2(new_n311), .A3(new_n318), .A4(new_n319), .ZN(new_n320));
  XOR2_X1   g134(.A(KEYINPUT9), .B(G234), .Z(new_n321));
  XNOR2_X1  g135(.A(new_n321), .B(KEYINPUT79), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n322), .A2(G217), .A3(new_n189), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT89), .B(G122), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G116), .ZN(new_n325));
  INV_X1    g139(.A(G107), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n236), .A2(G122), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n265), .A2(G128), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n208), .A2(G143), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n329), .A2(new_n227), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n227), .B1(new_n329), .B2(new_n330), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n328), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT90), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n334), .B1(new_n327), .B2(KEYINPUT14), .ZN(new_n335));
  INV_X1    g149(.A(G122), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n334), .B(KEYINPUT14), .C1(new_n336), .C2(G116), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n325), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT91), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n336), .A2(G116), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT14), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n325), .B(KEYINPUT91), .C1(new_n335), .C2(new_n338), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n341), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n333), .B1(new_n346), .B2(G107), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n329), .A2(KEYINPUT13), .A3(new_n330), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n348), .B(G134), .C1(KEYINPUT13), .C2(new_n329), .ZN(new_n349));
  OR2_X1    g163(.A1(KEYINPUT89), .A2(G122), .ZN(new_n350));
  NAND2_X1  g164(.A1(KEYINPUT89), .A2(G122), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n236), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(G107), .B1(new_n352), .B2(new_n342), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n328), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n331), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n349), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n323), .B1(new_n347), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT92), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n349), .A2(new_n354), .A3(new_n355), .ZN(new_n359));
  INV_X1    g173(.A(new_n323), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT90), .B1(new_n342), .B2(new_n343), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n352), .B1(new_n361), .B2(new_n337), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n362), .A2(KEYINPUT91), .B1(new_n343), .B2(new_n342), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n326), .B1(new_n363), .B2(new_n341), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n359), .B(new_n360), .C1(new_n364), .C2(new_n333), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n357), .A2(new_n358), .A3(new_n365), .ZN(new_n366));
  OAI211_X1 g180(.A(KEYINPUT92), .B(new_n323), .C1(new_n347), .C2(new_n356), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n300), .A3(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT93), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n366), .A2(KEYINPUT93), .A3(new_n300), .A4(new_n367), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT15), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G478), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(G113), .B(G122), .ZN(new_n377));
  INV_X1    g191(.A(G104), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n377), .B(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n188), .A2(new_n189), .A3(G214), .ZN(new_n380));
  OR2_X1    g194(.A1(new_n380), .A2(new_n201), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n265), .A2(new_n380), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n381), .A2(new_n382), .A3(new_n216), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n216), .B1(new_n381), .B2(new_n382), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT16), .ZN(new_n387));
  INV_X1    g201(.A(G140), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n388), .A3(G125), .ZN(new_n389));
  XNOR2_X1  g203(.A(G125), .B(G140), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  OAI211_X1 g205(.A(G146), .B(new_n389), .C1(new_n391), .C2(new_n387), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n390), .B(KEYINPUT75), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT19), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n391), .A2(KEYINPUT19), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n386), .B(new_n392), .C1(new_n397), .C2(G146), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n393), .A2(new_n206), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n390), .A2(new_n206), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n381), .A2(new_n382), .ZN(new_n403));
  NAND2_X1  g217(.A1(KEYINPUT18), .A2(G131), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n403), .A2(new_n404), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n402), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n379), .B1(new_n398), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n384), .A2(KEYINPUT17), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n389), .B1(new_n391), .B2(new_n387), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n206), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(new_n411), .A3(new_n392), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT17), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n412), .A2(KEYINPUT87), .B1(new_n413), .B2(new_n385), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT87), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n409), .A2(new_n415), .A3(new_n411), .A4(new_n392), .ZN(new_n416));
  OR2_X1    g230(.A1(new_n405), .A2(new_n406), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n414), .A2(new_n416), .B1(new_n402), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n408), .B1(new_n418), .B2(new_n379), .ZN(new_n419));
  NOR2_X1   g233(.A1(G475), .A2(G902), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(KEYINPUT20), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n412), .A2(KEYINPUT87), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n385), .A2(new_n413), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n424), .A3(new_n416), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(new_n379), .A3(new_n407), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n397), .A2(G146), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n392), .B1(new_n383), .B2(new_n384), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n407), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n379), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(new_n433), .A3(new_n420), .ZN(new_n434));
  INV_X1    g248(.A(new_n426), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n379), .B1(new_n425), .B2(new_n407), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n300), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(KEYINPUT88), .B(G475), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n422), .A2(new_n434), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n368), .A2(new_n375), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n376), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  XOR2_X1   g256(.A(KEYINPUT82), .B(KEYINPUT4), .Z(new_n443));
  NAND2_X1  g257(.A1(new_n326), .A2(G104), .ZN(new_n444));
  AND2_X1   g258(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n445));
  NOR2_X1   g259(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(G104), .A3(new_n326), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n378), .A2(G107), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI211_X1 g266(.A(G101), .B(new_n443), .C1(new_n448), .C2(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT81), .B(G101), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n447), .A2(new_n454), .A3(new_n450), .A4(new_n451), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT4), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n450), .A2(new_n451), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n197), .B1(new_n457), .B2(new_n447), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n243), .B(new_n453), .C1(new_n456), .C2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT5), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n460), .B1(new_n238), .B2(new_n239), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n460), .A2(new_n237), .A3(G116), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(G113), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n235), .ZN(new_n466));
  AOI22_X1  g280(.A1(new_n462), .A2(new_n465), .B1(new_n466), .B2(new_n241), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT85), .ZN(new_n468));
  OAI21_X1  g282(.A(KEYINPUT83), .B1(new_n326), .B2(G104), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT83), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(new_n378), .A3(G107), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n469), .A2(new_n471), .A3(new_n444), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G101), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n467), .A2(new_n468), .A3(new_n455), .A4(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n455), .A2(new_n473), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n242), .B1(new_n461), .B2(new_n464), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT85), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n459), .A2(new_n474), .A3(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(G110), .B(G122), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n459), .A2(new_n474), .A3(new_n477), .A4(new_n479), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n481), .A2(KEYINPUT6), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(G125), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n215), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n485), .B1(new_n484), .B2(new_n256), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n189), .A2(G224), .ZN(new_n487));
  XOR2_X1   g301(.A(new_n487), .B(KEYINPUT86), .Z(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n486), .B(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT6), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n478), .A2(new_n491), .A3(new_n480), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n483), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n487), .A2(KEYINPUT7), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n256), .A2(new_n484), .ZN(new_n495));
  AOI21_X1  g309(.A(G125), .B1(new_n268), .B2(new_n210), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n494), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n485), .B(new_n498), .C1(new_n484), .C2(new_n256), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n475), .B(new_n476), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n479), .B(KEYINPUT8), .ZN(new_n501));
  AOI22_X1  g315(.A1(new_n497), .A2(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(G902), .B1(new_n502), .B2(new_n482), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n493), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(G210), .B1(G237), .B2(G902), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n493), .A2(new_n505), .A3(new_n503), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(G234), .A2(G237), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(G952), .A3(new_n189), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n511), .A2(G902), .A3(G953), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT21), .B(G898), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n513), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(G214), .B1(G237), .B2(G902), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NOR3_X1   g334(.A1(new_n442), .A2(new_n510), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(G234), .ZN(new_n522));
  OAI21_X1  g336(.A(G217), .B1(new_n522), .B2(G902), .ZN(new_n523));
  XOR2_X1   g337(.A(KEYINPUT22), .B(G137), .Z(new_n524));
  NAND3_X1  g338(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n524), .B(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n526), .B(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n399), .A2(new_n392), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n237), .A2(G128), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n208), .A2(KEYINPUT23), .A3(G119), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n237), .A2(G128), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n530), .B(new_n531), .C1(new_n532), .C2(KEYINPUT23), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n533), .A2(G110), .ZN(new_n534));
  OR2_X1    g348(.A1(new_n534), .A2(KEYINPUT74), .ZN(new_n535));
  OR2_X1    g349(.A1(new_n532), .A2(KEYINPUT73), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n532), .A2(KEYINPUT73), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(new_n530), .A3(new_n537), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT24), .B(G110), .ZN(new_n539));
  AOI22_X1  g353(.A1(new_n534), .A2(KEYINPUT74), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n529), .B1(new_n535), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n411), .A2(new_n392), .ZN(new_n542));
  OR2_X1    g356(.A1(new_n538), .A2(new_n539), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n533), .A2(G110), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n528), .B1(new_n541), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n535), .A2(new_n540), .ZN(new_n548));
  INV_X1    g362(.A(new_n529), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n528), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n550), .A2(new_n551), .A3(new_n545), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n547), .A2(new_n552), .A3(new_n300), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n523), .B1(new_n553), .B2(KEYINPUT25), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT25), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n547), .A2(new_n552), .A3(new_n555), .A4(new_n300), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n523), .A2(new_n300), .ZN(new_n558));
  XOR2_X1   g372(.A(new_n558), .B(KEYINPUT78), .Z(new_n559));
  NAND3_X1  g373(.A1(new_n547), .A2(new_n552), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(G469), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT12), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n455), .A2(new_n473), .ZN(new_n565));
  INV_X1    g379(.A(new_n207), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n566), .B1(new_n265), .B2(G146), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT1), .B1(new_n265), .B2(G146), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n567), .B1(G128), .B2(new_n568), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n205), .A2(new_n207), .A3(new_n209), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n565), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n475), .A2(new_n268), .A3(new_n210), .ZN(new_n572));
  AOI211_X1 g386(.A(new_n564), .B(new_n250), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n567), .ZN(new_n574));
  AOI21_X1  g388(.A(G146), .B1(new_n202), .B2(new_n204), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT1), .ZN(new_n576));
  OAI21_X1  g390(.A(G128), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n570), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n572), .B1(new_n578), .B2(new_n475), .ZN(new_n579));
  INV_X1    g393(.A(new_n250), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT12), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n573), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT10), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n583), .B1(new_n578), .B2(new_n475), .ZN(new_n584));
  OAI21_X1  g398(.A(G101), .B1(new_n448), .B2(new_n452), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n585), .A2(KEYINPUT4), .A3(new_n455), .ZN(new_n586));
  AOI22_X1  g400(.A1(new_n266), .A2(new_n254), .B1(new_n567), .B2(new_n251), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n586), .A2(new_n587), .A3(new_n453), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n565), .A2(KEYINPUT10), .A3(new_n215), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n584), .A2(new_n250), .A3(new_n588), .A4(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(G110), .B(G140), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n189), .A2(G227), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n591), .B(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n582), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n584), .A2(new_n588), .A3(new_n589), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n580), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n594), .B1(new_n598), .B2(new_n590), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n563), .B(new_n300), .C1(new_n596), .C2(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n590), .B1(new_n573), .B2(new_n581), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n593), .ZN(new_n602));
  AOI21_X1  g416(.A(KEYINPUT84), .B1(new_n590), .B2(new_n594), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT84), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n598), .B1(new_n595), .B2(new_n604), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n602), .B(G469), .C1(new_n603), .C2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n563), .A2(new_n300), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n600), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n322), .A2(new_n300), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n610), .A2(G221), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n320), .A2(new_n521), .A3(new_n562), .A4(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(new_n615), .B(new_n454), .Z(G3));
  INV_X1    g430(.A(new_n519), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n493), .A2(new_n505), .A3(new_n503), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n617), .B1(new_n618), .B2(KEYINPUT94), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n619), .B(new_n518), .C1(new_n509), .C2(KEYINPUT94), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n433), .B1(new_n432), .B2(new_n420), .ZN(new_n621));
  AOI211_X1 g435(.A(KEYINPUT20), .B(new_n421), .C1(new_n426), .C2(new_n431), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n425), .A2(new_n407), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n430), .ZN(new_n624));
  AOI21_X1  g438(.A(G902), .B1(new_n624), .B2(new_n426), .ZN(new_n625));
  INV_X1    g439(.A(new_n438), .ZN(new_n626));
  OAI22_X1  g440(.A1(new_n621), .A2(new_n622), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(G478), .B1(new_n370), .B2(new_n371), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT33), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n366), .A2(new_n629), .A3(new_n367), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n357), .A2(KEYINPUT33), .A3(new_n365), .ZN(new_n631));
  AND4_X1   g445(.A1(G478), .A2(new_n630), .A3(new_n300), .A4(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n627), .B1(new_n628), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(KEYINPUT95), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT95), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n627), .B(new_n635), .C1(new_n628), .C2(new_n632), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n620), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(G902), .B1(new_n304), .B2(new_n309), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n310), .B1(new_n639), .B2(G472), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n613), .A2(new_n561), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n637), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT34), .B(G104), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  AOI21_X1  g458(.A(new_n374), .B1(new_n370), .B2(new_n371), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n439), .B1(new_n645), .B2(new_n440), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n620), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n647), .A2(new_n640), .A3(new_n641), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT35), .B(G107), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  INV_X1    g464(.A(KEYINPUT96), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n550), .A2(new_n651), .A3(new_n545), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n651), .B1(new_n550), .B2(new_n545), .ZN(new_n654));
  OAI22_X1  g468(.A1(new_n653), .A2(new_n654), .B1(KEYINPUT36), .B2(new_n528), .ZN(new_n655));
  INV_X1    g469(.A(new_n654), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n528), .A2(KEYINPUT36), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n656), .A2(new_n657), .A3(new_n652), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n655), .A2(new_n658), .A3(new_n559), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n557), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n521), .A2(new_n614), .A3(new_n640), .A4(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT37), .B(G110), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G12));
  INV_X1    g477(.A(G900), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n513), .B1(new_n515), .B2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  OAI211_X1 g480(.A(new_n439), .B(new_n666), .C1(new_n645), .C2(new_n440), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n609), .A2(new_n660), .A3(new_n612), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n619), .B1(new_n509), .B2(KEYINPUT94), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n320), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G128), .ZN(G30));
  NOR2_X1   g486(.A1(new_n271), .A2(new_n283), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(G902), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n289), .A2(new_n283), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n299), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n676), .B1(new_n310), .B2(KEYINPUT32), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n311), .A2(new_n677), .A3(new_n318), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(KEYINPUT97), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT97), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n311), .A2(new_n677), .A3(new_n318), .A4(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(new_n509), .B(KEYINPUT38), .Z(new_n683));
  OAI21_X1  g497(.A(new_n627), .B1(new_n645), .B2(new_n440), .ZN(new_n684));
  NOR4_X1   g498(.A1(new_n683), .A2(new_n617), .A3(new_n684), .A4(new_n660), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT98), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n682), .A2(KEYINPUT98), .A3(new_n685), .ZN(new_n689));
  XOR2_X1   g503(.A(new_n665), .B(KEYINPUT39), .Z(new_n690));
  NAND2_X1  g504(.A1(new_n614), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(new_n691), .B(KEYINPUT40), .Z(new_n692));
  NAND3_X1  g506(.A1(new_n688), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(new_n212), .ZN(G45));
  OAI211_X1 g508(.A(new_n627), .B(new_n666), .C1(new_n628), .C2(new_n632), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n695), .A2(new_n668), .A3(new_n669), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n320), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G146), .ZN(G48));
  NOR2_X1   g512(.A1(new_n596), .A2(new_n599), .ZN(new_n699));
  OAI21_X1  g513(.A(G469), .B1(new_n699), .B2(G902), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n700), .A2(new_n612), .A3(new_n600), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n637), .A2(new_n320), .A3(new_n562), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT41), .B(G113), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G15));
  NAND4_X1  g519(.A1(new_n320), .A2(new_n562), .A3(new_n647), .A4(new_n702), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G116), .ZN(G18));
  AOI21_X1  g521(.A(new_n442), .B1(new_n557), .B2(new_n659), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n669), .A2(new_n701), .A3(new_n517), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n320), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G119), .ZN(G21));
  NOR2_X1   g525(.A1(new_n684), .A2(new_n669), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n272), .A2(new_n302), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n199), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n301), .B1(new_n309), .B2(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n715), .B1(new_n639), .B2(G472), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n701), .A2(new_n517), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n712), .A2(new_n716), .A3(new_n562), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G122), .ZN(G24));
  INV_X1    g533(.A(new_n715), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n720), .B(new_n660), .C1(new_n638), .C2(new_n299), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n721), .A2(new_n695), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n669), .A2(new_n701), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G125), .ZN(G27));
  AOI21_X1  g539(.A(new_n505), .B1(new_n493), .B2(new_n503), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n618), .A2(new_n726), .A3(new_n617), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(new_n609), .A3(new_n612), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(KEYINPUT99), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT99), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n727), .A2(new_n609), .A3(new_n730), .A4(new_n612), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n695), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n320), .A2(new_n732), .A3(new_n562), .A4(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT42), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT100), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n319), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n310), .A2(KEYINPUT100), .A3(KEYINPUT32), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n310), .ZN(new_n741));
  AOI22_X1  g555(.A1(new_n313), .A2(new_n741), .B1(new_n297), .B2(G472), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n561), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  AOI211_X1 g557(.A(new_n735), .B(new_n695), .C1(new_n729), .C2(new_n731), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n736), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(KEYINPUT101), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT101), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n736), .A2(new_n745), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(KEYINPUT102), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(new_n229), .ZN(G33));
  INV_X1    g566(.A(new_n667), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n320), .A2(new_n732), .A3(new_n562), .A4(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G134), .ZN(G36));
  OR2_X1    g569(.A1(new_n628), .A2(new_n632), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n439), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT43), .ZN(new_n758));
  INV_X1    g572(.A(new_n640), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT43), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n756), .A2(new_n760), .A3(new_n439), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n758), .A2(new_n759), .A3(new_n660), .A4(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT44), .ZN(new_n763));
  OAI211_X1 g577(.A(KEYINPUT103), .B(new_n727), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  INV_X1    g579(.A(new_n600), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n602), .B1(new_n605), .B2(new_n603), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT45), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n563), .B1(new_n767), .B2(new_n768), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n608), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT46), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n766), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n771), .A2(KEYINPUT46), .A3(new_n608), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n611), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n764), .A2(new_n690), .A3(new_n765), .A4(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT103), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n727), .B1(new_n762), .B2(new_n763), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(new_n218), .ZN(G39));
  INV_X1    g595(.A(KEYINPUT47), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT104), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n776), .A2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n776), .A2(new_n783), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n782), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n786), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n788), .A2(KEYINPUT47), .A3(new_n784), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n727), .ZN(new_n791));
  NOR4_X1   g605(.A1(new_n320), .A2(new_n562), .A3(new_n695), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G140), .ZN(G42));
  INV_X1    g608(.A(new_n682), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n702), .A2(new_n727), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n796), .A2(new_n561), .A3(new_n512), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n756), .A2(new_n627), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n795), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT114), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT113), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n758), .A2(new_n761), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n716), .A2(new_n562), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n513), .A3(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n702), .A2(KEYINPUT112), .A3(new_n617), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT112), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n806), .B1(new_n701), .B2(new_n519), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n805), .A2(new_n683), .A3(new_n807), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n801), .B(KEYINPUT50), .C1(new_n804), .C2(new_n808), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n802), .A2(new_n513), .ZN(new_n810));
  INV_X1    g624(.A(new_n796), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n810), .A2(new_n660), .A3(new_n716), .A4(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n801), .B1(new_n804), .B2(new_n808), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT50), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AND4_X1   g629(.A1(new_n800), .A2(new_n809), .A3(new_n812), .A4(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n804), .A2(new_n791), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(KEYINPUT111), .ZN(new_n818));
  INV_X1    g632(.A(new_n700), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(new_n766), .ZN(new_n820));
  XOR2_X1   g634(.A(new_n820), .B(KEYINPUT106), .Z(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n822), .A2(new_n612), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n818), .B1(new_n790), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT51), .B1(new_n816), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n810), .A2(new_n743), .A3(new_n811), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(KEYINPUT48), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n810), .A2(new_n723), .A3(new_n803), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n634), .A2(new_n636), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n795), .A2(new_n829), .A3(new_n797), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n827), .A2(new_n828), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n825), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n703), .A2(new_n706), .A3(new_n710), .A4(new_n718), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n646), .A2(new_n633), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n510), .A2(new_n520), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n640), .A2(new_n834), .A3(new_n835), .A4(new_n641), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n615), .A2(new_n661), .A3(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n722), .A2(new_n732), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n754), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT107), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n728), .A2(new_n665), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n320), .A2(new_n708), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n320), .A2(new_n708), .A3(new_n842), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT107), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n840), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n747), .A2(new_n838), .A3(new_n846), .A4(new_n749), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n671), .A2(new_n697), .A3(new_n724), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT108), .B1(new_n660), .B2(new_n665), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT108), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n557), .A2(new_n659), .A3(new_n850), .A4(new_n666), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n712), .A2(new_n614), .A3(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n682), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n848), .A2(KEYINPUT52), .A3(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT52), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n671), .A2(new_n697), .A3(new_n724), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n853), .B1(new_n679), .B2(new_n681), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT53), .B1(new_n847), .B2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT109), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n856), .A2(new_n863), .A3(new_n860), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n863), .B1(new_n856), .B2(new_n860), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n736), .A2(new_n748), .A3(new_n745), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n748), .B1(new_n736), .B2(new_n745), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT53), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n869), .A2(new_n870), .A3(new_n838), .A4(new_n846), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n862), .B(KEYINPUT54), .C1(new_n866), .C2(new_n871), .ZN(new_n872));
  AND4_X1   g686(.A1(new_n703), .A2(new_n706), .A3(new_n710), .A4(new_n718), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT110), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n873), .A2(new_n746), .A3(new_n874), .ZN(new_n875));
  AOI22_X1  g689(.A1(new_n735), .A2(new_n734), .B1(new_n743), .B2(new_n744), .ZN(new_n876));
  OAI21_X1  g690(.A(KEYINPUT110), .B1(new_n876), .B2(new_n833), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n837), .A2(new_n870), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n846), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n878), .B(new_n880), .C1(new_n864), .C2(new_n865), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n870), .B1(new_n847), .B2(new_n861), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n872), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n815), .A2(new_n809), .A3(new_n812), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n824), .A2(KEYINPUT51), .A3(new_n800), .A4(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT115), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n888), .A2(new_n889), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n832), .B(new_n886), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT116), .ZN(new_n893));
  OAI211_X1 g707(.A(G952), .B(new_n189), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(G953), .B1(new_n892), .B2(KEYINPUT116), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT49), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n683), .B1(new_n821), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n822), .A2(KEYINPUT49), .ZN(new_n898));
  OR4_X1    g712(.A1(new_n561), .A2(new_n757), .A3(new_n617), .A4(new_n611), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  AOI211_X1 g714(.A(new_n897), .B(new_n898), .C1(KEYINPUT105), .C2(new_n900), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n901), .B(new_n795), .C1(KEYINPUT105), .C2(new_n900), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n894), .A2(new_n895), .A3(new_n902), .ZN(G75));
  OR2_X1    g717(.A1(new_n189), .A2(G952), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT118), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n300), .B1(new_n881), .B2(new_n882), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(G210), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT117), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n909), .A2(KEYINPUT56), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(KEYINPUT55), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT55), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n908), .A2(new_n913), .A3(new_n910), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n483), .A2(new_n492), .ZN(new_n916));
  INV_X1    g730(.A(new_n490), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n918), .A2(new_n493), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n915), .A2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n919), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n912), .A2(new_n921), .A3(new_n914), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n906), .B1(new_n920), .B2(new_n922), .ZN(G51));
  NAND2_X1  g737(.A1(new_n881), .A2(new_n882), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(KEYINPUT54), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n884), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n607), .B(KEYINPUT57), .Z(new_n928));
  OAI22_X1  g742(.A1(new_n927), .A2(new_n928), .B1(new_n599), .B2(new_n596), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n907), .A2(new_n769), .A3(new_n770), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n906), .B1(new_n929), .B2(new_n930), .ZN(G54));
  NAND3_X1  g745(.A1(new_n907), .A2(KEYINPUT58), .A3(G475), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n932), .A2(KEYINPUT119), .A3(new_n419), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n905), .B1(new_n932), .B2(new_n419), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT119), .B1(new_n932), .B2(new_n419), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(G60));
  NAND2_X1  g750(.A1(G478), .A2(G902), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT59), .Z(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n885), .A2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT120), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n630), .A2(new_n631), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n938), .B1(new_n872), .B2(new_n884), .ZN(new_n944));
  INV_X1    g758(.A(new_n942), .ZN(new_n945));
  OAI21_X1  g759(.A(KEYINPUT120), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n942), .A2(new_n938), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n906), .B1(new_n926), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n943), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT121), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n943), .A2(new_n948), .A3(new_n946), .A4(KEYINPUT121), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(G63));
  AND2_X1   g767(.A1(new_n655), .A2(new_n658), .ZN(new_n954));
  NAND2_X1  g768(.A1(G217), .A2(G902), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT60), .Z(new_n956));
  NAND3_X1  g770(.A1(new_n924), .A2(KEYINPUT122), .A3(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT122), .B1(new_n924), .B2(new_n956), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n954), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n959), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n547), .A2(new_n552), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n961), .A2(new_n962), .A3(new_n957), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n960), .A2(new_n963), .A3(new_n905), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT61), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n960), .A2(new_n963), .A3(KEYINPUT61), .A4(new_n905), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(G66));
  INV_X1    g782(.A(G224), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n516), .A2(new_n969), .A3(new_n189), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n970), .B1(new_n838), .B2(new_n189), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n916), .B1(G898), .B2(new_n189), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(G69));
  INV_X1    g787(.A(new_n777), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n779), .A2(new_n778), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n320), .A2(new_n562), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  AOI211_X1 g791(.A(new_n791), .B(new_n691), .C1(new_n633), .C2(new_n646), .ZN(new_n978));
  AOI22_X1  g792(.A1(new_n974), .A2(new_n975), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n693), .A2(new_n848), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(KEYINPUT62), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n979), .A2(new_n981), .A3(new_n793), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n980), .A2(KEYINPUT62), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n189), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n279), .A2(new_n280), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(new_n397), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(new_n754), .ZN(new_n988));
  OAI21_X1  g802(.A(KEYINPUT123), .B1(new_n750), .B2(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT123), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n869), .A2(new_n990), .A3(new_n754), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n776), .A2(new_n690), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n743), .A2(new_n712), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n848), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n780), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n992), .A2(new_n189), .A3(new_n996), .A4(new_n793), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n987), .B1(G900), .B2(G953), .ZN(new_n998));
  AOI22_X1  g812(.A1(new_n984), .A2(new_n987), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n1001));
  AOI21_X1  g815(.A(KEYINPUT125), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT125), .ZN(new_n1003));
  INV_X1    g817(.A(new_n1001), .ZN(new_n1004));
  NOR3_X1   g818(.A1(new_n999), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  AND3_X1   g819(.A1(new_n999), .A2(KEYINPUT124), .A3(new_n1004), .ZN(new_n1006));
  AOI21_X1  g820(.A(KEYINPUT124), .B1(new_n999), .B2(new_n1004), .ZN(new_n1007));
  OAI22_X1  g821(.A1(new_n1002), .A2(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(G72));
  NOR2_X1   g822(.A1(new_n982), .A2(new_n983), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(new_n838), .ZN(new_n1010));
  XNOR2_X1  g824(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1011));
  NAND2_X1  g825(.A1(G472), .A2(G902), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1011), .B(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n675), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n289), .A2(new_n283), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n1015), .B(KEYINPUT127), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n992), .A2(new_n793), .A3(new_n996), .A4(new_n838), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1016), .B1(new_n1017), .B2(new_n1013), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n862), .B1(new_n866), .B2(new_n871), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1015), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n1020), .A2(new_n675), .A3(new_n1013), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n905), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  NOR3_X1   g836(.A1(new_n1014), .A2(new_n1018), .A3(new_n1022), .ZN(G57));
endmodule


