//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 0 0 0 0 0 0 0 1 0 1 1 0 0 1 1 0 1 1 0 1 1 1 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n762, new_n763, new_n764,
    new_n765, new_n767, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n843, new_n844, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951;
  INV_X1    g000(.A(G50gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G43gat), .ZN(new_n203));
  INV_X1    g002(.A(G43gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G50gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(new_n205), .A3(KEYINPUT15), .ZN(new_n206));
  NAND2_X1  g005(.A1(G29gat), .A2(G36gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n209));
  OR3_X1    g008(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT15), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n203), .A2(KEYINPUT89), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(new_n205), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n203), .A2(KEYINPUT89), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n212), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n211), .B1(new_n216), .B2(KEYINPUT90), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n216), .A2(KEYINPUT90), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n209), .A2(KEYINPUT88), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n209), .A2(KEYINPUT88), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(new_n220), .A3(new_n210), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n221), .A2(new_n207), .ZN(new_n222));
  OAI22_X1  g021(.A1(new_n217), .A2(new_n218), .B1(new_n206), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G85gat), .A2(G92gat), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n224), .B(KEYINPUT7), .ZN(new_n225));
  NAND2_X1  g024(.A1(G99gat), .A2(G106gat), .ZN(new_n226));
  INV_X1    g025(.A(G85gat), .ZN(new_n227));
  INV_X1    g026(.A(G92gat), .ZN(new_n228));
  AOI22_X1  g027(.A1(KEYINPUT8), .A2(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT98), .ZN(new_n230));
  XNOR2_X1  g029(.A(G99gat), .B(G106gat), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n225), .B(new_n229), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n230), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n232), .B(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n223), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  XOR2_X1   g037(.A(new_n238), .B(KEYINPUT99), .Z(new_n239));
  XNOR2_X1  g038(.A(new_n223), .B(KEYINPUT17), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(new_n234), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G190gat), .B(G218gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n243), .B(KEYINPUT100), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n242), .B(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT97), .ZN(new_n246));
  XNOR2_X1  g045(.A(G134gat), .B(G162gat), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(new_n249), .B(KEYINPUT101), .Z(new_n250));
  XNOR2_X1  g049(.A(new_n246), .B(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT16), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n253), .A2(G1gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(G15gat), .B(G22gat), .ZN(new_n255));
  MUX2_X1   g054(.A(G1gat), .B(new_n254), .S(new_n255), .Z(new_n256));
  XOR2_X1   g055(.A(new_n256), .B(G8gat), .Z(new_n257));
  INV_X1    g056(.A(G71gat), .ZN(new_n258));
  INV_X1    g057(.A(G78gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g059(.A1(G71gat), .A2(G78gat), .ZN(new_n261));
  XOR2_X1   g060(.A(G57gat), .B(G64gat), .Z(new_n262));
  AOI211_X1 g061(.A(new_n260), .B(new_n261), .C1(new_n262), .C2(KEYINPUT9), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(KEYINPUT9), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n264), .B1(new_n258), .B2(new_n259), .ZN(new_n265));
  XNOR2_X1  g064(.A(G57gat), .B(G64gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(KEYINPUT94), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n263), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT95), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n257), .B1(new_n270), .B2(KEYINPUT21), .ZN(new_n271));
  XNOR2_X1  g070(.A(G127gat), .B(G155gat), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT21), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n275), .B(KEYINPUT96), .ZN(new_n276));
  INV_X1    g075(.A(G231gat), .ZN(new_n277));
  INV_X1    g076(.A(G233gat), .ZN(new_n278));
  NOR3_X1   g077(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G231gat), .A2(G233gat), .ZN(new_n280));
  AND2_X1   g079(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n273), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NOR3_X1   g082(.A1(new_n279), .A2(new_n281), .A3(new_n273), .ZN(new_n284));
  XOR2_X1   g083(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n285));
  NOR3_X1   g084(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n285), .ZN(new_n287));
  OR3_X1    g086(.A1(new_n279), .A2(new_n281), .A3(new_n273), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n287), .B1(new_n288), .B2(new_n282), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n271), .B1(new_n286), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n285), .B1(new_n283), .B2(new_n284), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n288), .A2(new_n282), .A3(new_n287), .ZN(new_n292));
  INV_X1    g091(.A(new_n271), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  XOR2_X1   g093(.A(G183gat), .B(G211gat), .Z(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n290), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n296), .B1(new_n290), .B2(new_n294), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n252), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT102), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI211_X1 g100(.A(KEYINPUT102), .B(new_n252), .C1(new_n297), .C2(new_n298), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  XOR2_X1   g102(.A(G113gat), .B(G141gat), .Z(new_n304));
  XNOR2_X1  g103(.A(new_n304), .B(KEYINPUT11), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n305), .B(KEYINPUT87), .ZN(new_n306));
  XOR2_X1   g105(.A(G169gat), .B(G197gat), .Z(new_n307));
  XNOR2_X1  g106(.A(new_n306), .B(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n308), .B(KEYINPUT12), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n257), .A2(new_n223), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT91), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n310), .B(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n257), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n240), .A2(new_n313), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(G229gat), .A2(G233gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n315), .A2(KEYINPUT18), .A3(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n312), .B1(new_n257), .B2(new_n223), .ZN(new_n318));
  XOR2_X1   g117(.A(new_n316), .B(KEYINPUT13), .Z(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AND2_X1   g119(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n315), .A2(new_n316), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT18), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n309), .B1(new_n321), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT92), .ZN(new_n326));
  OR2_X1    g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n326), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT93), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n324), .B(new_n329), .ZN(new_n330));
  AND2_X1   g129(.A1(new_n321), .A2(new_n309), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n327), .A2(new_n328), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n269), .A2(new_n234), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT10), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n235), .A2(new_n268), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n270), .A2(KEYINPUT10), .A3(new_n235), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(KEYINPUT103), .ZN(new_n340));
  NAND2_X1  g139(.A1(G230gat), .A2(G233gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n334), .A2(new_n336), .ZN(new_n343));
  INV_X1    g142(.A(new_n341), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  XOR2_X1   g144(.A(G120gat), .B(G148gat), .Z(new_n346));
  XNOR2_X1  g145(.A(new_n346), .B(KEYINPUT104), .ZN(new_n347));
  XOR2_X1   g146(.A(G176gat), .B(G204gat), .Z(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(KEYINPUT105), .ZN(new_n349));
  XOR2_X1   g148(.A(new_n347), .B(new_n349), .Z(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n342), .A2(new_n345), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n339), .A2(new_n341), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(new_n345), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(new_n350), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n333), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n303), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G228gat), .A2(G233gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(G141gat), .B(G148gat), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(G155gat), .ZN(new_n364));
  INV_X1    g163(.A(G162gat), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT2), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n364), .B(new_n365), .C1(new_n366), .C2(KEYINPUT78), .ZN(new_n367));
  NAND2_X1  g166(.A1(G155gat), .A2(G162gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT78), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n366), .B1(G155gat), .B2(G162gat), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n363), .B(new_n369), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n364), .A2(new_n365), .A3(KEYINPUT77), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT77), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n374), .B1(G155gat), .B2(G162gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n376), .B(new_n368), .C1(KEYINPUT2), .C2(new_n362), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n372), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G197gat), .B(G204gat), .ZN(new_n379));
  INV_X1    g178(.A(G211gat), .ZN(new_n380));
  OR2_X1    g179(.A1(KEYINPUT73), .A2(G218gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(KEYINPUT73), .A2(G218gat), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n380), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n379), .B1(new_n383), .B2(KEYINPUT22), .ZN(new_n384));
  XOR2_X1   g183(.A(G211gat), .B(G218gat), .Z(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n385), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n387), .B(new_n379), .C1(KEYINPUT22), .C2(new_n383), .ZN(new_n388));
  AOI21_X1  g187(.A(KEYINPUT29), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n378), .B1(new_n389), .B2(KEYINPUT3), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT81), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n361), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n386), .A2(new_n388), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT3), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n372), .A2(new_n395), .A3(new_n377), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT29), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n390), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n392), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(G22gat), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n390), .B(new_n399), .C1(new_n391), .C2(new_n361), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT82), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n402), .B1(new_n401), .B2(new_n403), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n406), .A2(KEYINPUT82), .A3(new_n404), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n407), .A2(new_n404), .ZN(new_n410));
  XNOR2_X1  g209(.A(G78gat), .B(G106gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT31), .B(G50gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT80), .ZN(new_n414));
  AOI22_X1  g213(.A1(new_n408), .A2(new_n409), .B1(new_n410), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n413), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT80), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n410), .A2(new_n414), .ZN(new_n418));
  OAI22_X1  g217(.A1(new_n415), .A2(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT70), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT68), .ZN(new_n421));
  INV_X1    g220(.A(G127gat), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n422), .A2(G134gat), .ZN(new_n423));
  INV_X1    g222(.A(G134gat), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n424), .A2(G127gat), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n421), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(G127gat), .B(G134gat), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT68), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(G113gat), .ZN(new_n431));
  INV_X1    g230(.A(G120gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT1), .ZN(new_n434));
  NAND2_X1  g233(.A1(G113gat), .A2(G120gat), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n427), .B1(new_n430), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n433), .A2(new_n435), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT69), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n433), .A2(KEYINPUT69), .A3(new_n435), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n440), .B1(new_n428), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n434), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n437), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT66), .ZN(new_n445));
  NOR2_X1   g244(.A1(G169gat), .A2(G176gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(G169gat), .A2(G176gat), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n446), .B1(KEYINPUT23), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT25), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT23), .ZN(new_n450));
  NOR3_X1   g249(.A1(new_n450), .A2(G169gat), .A3(G176gat), .ZN(new_n451));
  NOR3_X1   g250(.A1(new_n448), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(G183gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT64), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT64), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(G183gat), .ZN(new_n456));
  INV_X1    g255(.A(G190gat), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n454), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(G183gat), .A2(G190gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT24), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT24), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n461), .A2(G183gat), .A3(G190gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n458), .A2(new_n463), .A3(KEYINPUT65), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n452), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(KEYINPUT64), .B(G183gat), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n466), .A2(new_n457), .B1(new_n460), .B2(new_n462), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n467), .A2(KEYINPUT65), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n445), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n458), .A2(new_n463), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT65), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n472), .A2(KEYINPUT66), .A3(new_n464), .A4(new_n452), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n446), .A2(KEYINPUT23), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n450), .B1(G169gat), .B2(G176gat), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n474), .B1(new_n475), .B2(new_n446), .ZN(new_n476));
  AOI22_X1  g275(.A1(new_n460), .A2(new_n462), .B1(new_n453), .B2(new_n457), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n449), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n469), .A2(new_n473), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT28), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT27), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n466), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n480), .B(new_n457), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n446), .A2(KEYINPUT26), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n459), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n446), .A2(KEYINPUT26), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n486), .B1(new_n447), .B2(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(KEYINPUT27), .B(G183gat), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT67), .ZN(new_n490));
  OR2_X1    g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n490), .ZN(new_n492));
  AOI21_X1  g291(.A(G190gat), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n484), .B(new_n488), .C1(new_n493), .C2(new_n480), .ZN(new_n494));
  AOI211_X1 g293(.A(new_n420), .B(new_n444), .C1(new_n479), .C2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n473), .A2(new_n478), .ZN(new_n496));
  OAI211_X1 g295(.A(KEYINPUT25), .B(new_n474), .C1(new_n475), .C2(new_n446), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n497), .B1(new_n467), .B2(KEYINPUT65), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT66), .B1(new_n498), .B2(new_n472), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n494), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n436), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n426), .B1(new_n501), .B2(new_n429), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n502), .B1(new_n434), .B2(new_n442), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT70), .B1(new_n500), .B2(new_n503), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n495), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(G227gat), .A2(G233gat), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT32), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT33), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n509), .B1(new_n506), .B2(new_n507), .ZN(new_n510));
  XOR2_X1   g309(.A(G15gat), .B(G43gat), .Z(new_n511));
  XNOR2_X1  g310(.A(G71gat), .B(G99gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n508), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n513), .ZN(new_n515));
  OAI221_X1 g314(.A(KEYINPUT32), .B1(new_n509), .B2(new_n515), .C1(new_n506), .C2(new_n507), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n506), .A2(new_n507), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT34), .ZN(new_n519));
  INV_X1    g318(.A(new_n495), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n504), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT34), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n520), .A2(new_n521), .A3(new_n522), .A4(new_n507), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT71), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT71), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n506), .A2(new_n525), .A3(new_n522), .A4(new_n507), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n519), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n517), .A2(new_n527), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n519), .A2(new_n524), .A3(new_n526), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n529), .A2(new_n516), .A3(new_n514), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n419), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G1gat), .B(G29gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(KEYINPUT0), .ZN(new_n533));
  XNOR2_X1  g332(.A(G57gat), .B(G85gat), .ZN(new_n534));
  XOR2_X1   g333(.A(new_n533), .B(new_n534), .Z(new_n535));
  INV_X1    g334(.A(KEYINPUT4), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n536), .B1(new_n503), .B2(new_n378), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n378), .A2(KEYINPUT3), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n503), .A2(new_n538), .A3(new_n396), .ZN(new_n539));
  INV_X1    g338(.A(new_n378), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n444), .A2(KEYINPUT4), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G225gat), .A2(G233gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(KEYINPUT79), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n537), .A2(new_n539), .A3(new_n541), .A4(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT5), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n444), .A2(new_n540), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n503), .A2(new_n378), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n543), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n546), .B1(new_n545), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n535), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT6), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n545), .A2(new_n551), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT5), .ZN(new_n558));
  INV_X1    g357(.A(new_n535), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n558), .A2(new_n559), .A3(new_n547), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n560), .A2(new_n554), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G8gat), .B(G36gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(G64gat), .B(G92gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT74), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT29), .B1(new_n479), .B2(new_n494), .ZN(new_n569));
  NAND2_X1  g368(.A1(G226gat), .A2(G233gat), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n568), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n500), .A2(new_n397), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n573), .A2(KEYINPUT74), .A3(new_n570), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n500), .A2(new_n571), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n572), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(new_n394), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n575), .B(new_n393), .C1(new_n569), .C2(new_n571), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT75), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n573), .A2(new_n570), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n581), .A2(KEYINPUT75), .A3(new_n393), .A4(new_n575), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n567), .B1(new_n577), .B2(new_n583), .ZN(new_n584));
  AND3_X1   g383(.A1(new_n577), .A2(new_n583), .A3(new_n567), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n584), .B1(new_n585), .B2(KEYINPUT30), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n577), .A2(new_n583), .A3(new_n567), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT76), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT30), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n588), .B1(new_n587), .B2(new_n589), .ZN(new_n591));
  OAI211_X1 g390(.A(new_n563), .B(new_n586), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT35), .B1(new_n531), .B2(new_n592), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n519), .A2(new_n526), .ZN(new_n594));
  AOI22_X1  g393(.A1(new_n594), .A2(new_n524), .B1(new_n514), .B2(new_n516), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT72), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n596), .B1(new_n517), .B2(new_n527), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n529), .A2(KEYINPUT72), .A3(new_n516), .A4(new_n514), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n595), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(new_n419), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n577), .A2(new_n583), .A3(KEYINPUT30), .A4(new_n567), .ZN(new_n601));
  AOI22_X1  g400(.A1(new_n394), .A2(new_n576), .B1(new_n580), .B2(new_n582), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n601), .B1(new_n602), .B2(new_n567), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n589), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(KEYINPUT76), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n603), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT35), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT84), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n609), .B1(new_n548), .B2(new_n552), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n558), .A2(KEYINPUT84), .A3(new_n547), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n535), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n562), .B1(new_n612), .B2(new_n555), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n607), .A2(new_n608), .A3(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n593), .B1(new_n600), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT37), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n581), .A2(new_n575), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n616), .B1(new_n617), .B2(new_n394), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n576), .A2(new_n393), .ZN(new_n619));
  AOI211_X1 g418(.A(KEYINPUT38), .B(new_n567), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT86), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n621), .B1(new_n602), .B2(new_n616), .ZN(new_n622));
  AND4_X1   g421(.A1(new_n621), .A2(new_n577), .A3(new_n583), .A4(new_n616), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n620), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI211_X1 g423(.A(new_n562), .B(new_n587), .C1(new_n612), .C2(new_n555), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT38), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n577), .A2(new_n583), .A3(new_n616), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(KEYINPUT86), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n602), .A2(new_n621), .A3(new_n616), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n577), .A2(new_n583), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n567), .B1(new_n633), .B2(KEYINPUT37), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n628), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n419), .B1(new_n627), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n586), .B1(new_n590), .B2(new_n591), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT39), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n549), .A2(new_n550), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n544), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT83), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n638), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n537), .A2(new_n539), .A3(new_n541), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n543), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n639), .A2(KEYINPUT83), .A3(new_n544), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n642), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n643), .A2(new_n638), .A3(new_n543), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n646), .A2(new_n535), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT40), .ZN(new_n649));
  OR2_X1    g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n612), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n648), .A2(new_n649), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(KEYINPUT85), .B1(new_n637), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n637), .A2(new_n653), .A3(KEYINPUT85), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n636), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n530), .A2(new_n528), .A3(KEYINPUT36), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n658), .B1(new_n599), .B2(KEYINPUT36), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n418), .A2(new_n417), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n408), .A2(new_n409), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(new_n418), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n660), .B1(new_n662), .B2(new_n413), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n592), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n659), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n615), .B1(new_n657), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n359), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n563), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g470(.A(KEYINPUT16), .B(G8gat), .Z(new_n672));
  NAND3_X1  g471(.A1(new_n668), .A2(new_n637), .A3(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n673), .A2(KEYINPUT42), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n668), .A2(new_n637), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n675), .B1(new_n676), .B2(G8gat), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n674), .B1(new_n673), .B2(new_n677), .ZN(G1325gat));
  INV_X1    g477(.A(new_n599), .ZN(new_n679));
  OR3_X1    g478(.A1(new_n667), .A2(G15gat), .A3(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(G15gat), .B1(new_n667), .B2(new_n659), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT106), .ZN(G1326gat));
  NOR2_X1   g482(.A1(new_n667), .A2(new_n419), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT107), .ZN(new_n685));
  XNOR2_X1  g484(.A(KEYINPUT43), .B(G22gat), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n685), .B(new_n686), .Z(G1327gat));
  NOR2_X1   g486(.A1(new_n297), .A2(new_n298), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n689), .A2(new_n358), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n634), .B1(new_n622), .B2(new_n623), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(KEYINPUT38), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n625), .B1(new_n632), .B2(new_n620), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n663), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT85), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n607), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n694), .B1(new_n697), .B2(new_n654), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n698), .A2(new_n664), .A3(new_n659), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n252), .B1(new_n699), .B2(new_n615), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n690), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(G29gat), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n701), .A2(new_n702), .A3(new_n669), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT45), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n705), .B1(new_n666), .B2(new_n251), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT108), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(KEYINPUT108), .B1(new_n700), .B2(new_n705), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n664), .A2(KEYINPUT109), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT109), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n592), .A2(new_n711), .A3(new_n663), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n713), .A2(new_n698), .A3(new_n659), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n615), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n715), .A2(new_n705), .A3(new_n251), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n708), .A2(new_n709), .A3(new_n716), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n717), .A2(new_n690), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n718), .A2(new_n669), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n704), .B1(new_n719), .B2(new_n702), .ZN(G1328gat));
  INV_X1    g519(.A(G36gat), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n701), .A2(new_n721), .A3(new_n637), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT46), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n721), .B1(new_n718), .B2(new_n637), .ZN(new_n724));
  OR2_X1    g523(.A1(new_n723), .A2(new_n724), .ZN(G1329gat));
  INV_X1    g524(.A(new_n659), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n718), .A2(G43gat), .A3(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n701), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n204), .B1(new_n728), .B2(new_n679), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g530(.A(new_n716), .B1(new_n706), .B2(new_n707), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n700), .A2(KEYINPUT108), .A3(new_n705), .ZN(new_n733));
  OAI211_X1 g532(.A(new_n663), .B(new_n690), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(KEYINPUT112), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT112), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n717), .A2(new_n736), .A3(new_n663), .A4(new_n690), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n202), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n419), .A2(G50gat), .ZN(new_n739));
  XOR2_X1   g538(.A(new_n739), .B(KEYINPUT111), .Z(new_n740));
  NOR2_X1   g539(.A1(new_n728), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(KEYINPUT48), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT113), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n734), .A2(G50gat), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n741), .A2(KEYINPUT48), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n734), .A2(KEYINPUT110), .A3(G50gat), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  AND3_X1   g548(.A1(new_n742), .A2(new_n743), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n743), .B1(new_n742), .B2(new_n749), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n750), .A2(new_n751), .ZN(G1331gat));
  NOR3_X1   g551(.A1(new_n303), .A2(new_n333), .A3(new_n357), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n753), .A2(new_n715), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n669), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g555(.A(new_n607), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT114), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n759), .B(new_n760), .Z(G1333gat));
  NAND3_X1  g560(.A1(new_n754), .A2(new_n258), .A3(new_n599), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n754), .A2(new_n726), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n762), .B1(new_n763), .B2(new_n258), .ZN(new_n764));
  XOR2_X1   g563(.A(KEYINPUT115), .B(KEYINPUT50), .Z(new_n765));
  XNOR2_X1  g564(.A(new_n764), .B(new_n765), .ZN(G1334gat));
  NAND2_X1  g565(.A1(new_n754), .A2(new_n663), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g567(.A1(new_n689), .A2(new_n333), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n252), .B1(new_n714), .B2(new_n615), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n356), .A2(new_n227), .A3(new_n669), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT118), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n689), .A2(new_n333), .A3(new_n357), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(KEYINPUT116), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n717), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT117), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n778), .A2(KEYINPUT117), .A3(new_n717), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n782), .A2(new_n563), .A3(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n776), .B1(new_n785), .B2(new_n227), .ZN(G1336gat));
  NAND4_X1  g585(.A1(new_n773), .A2(new_n228), .A3(new_n637), .A4(new_n356), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n778), .A2(new_n637), .A3(new_n717), .ZN(new_n788));
  AOI21_X1  g587(.A(KEYINPUT52), .B1(new_n788), .B2(G92gat), .ZN(new_n789));
  AND2_X1   g588(.A1(KEYINPUT119), .A2(KEYINPUT52), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n787), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n787), .A2(KEYINPUT119), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n781), .A2(new_n637), .A3(new_n783), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n792), .B1(new_n793), .B2(G92gat), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n791), .B1(new_n794), .B2(new_n795), .ZN(G1337gat));
  NAND2_X1  g595(.A1(new_n726), .A2(G99gat), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n782), .A2(new_n784), .A3(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(G99gat), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n773), .A2(new_n599), .A3(new_n356), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(G1338gat));
  XNOR2_X1  g600(.A(KEYINPUT120), .B(G106gat), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n802), .B1(new_n779), .B2(new_n419), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n773), .A2(new_n356), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n419), .A2(G106gat), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n803), .B(new_n804), .C1(new_n805), .C2(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n805), .A2(new_n807), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n781), .A2(new_n663), .A3(new_n783), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n809), .B1(new_n810), .B2(new_n802), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n808), .B1(new_n811), .B2(new_n804), .ZN(G1339gat));
  NAND2_X1  g611(.A1(new_n607), .A2(new_n669), .ZN(new_n813));
  INV_X1    g612(.A(new_n333), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n301), .A2(new_n302), .A3(new_n814), .A4(new_n357), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n350), .B1(new_n353), .B2(KEYINPUT54), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n817));
  INV_X1    g616(.A(new_n339), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n817), .B1(new_n818), .B2(new_n344), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n816), .B1(new_n342), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n352), .B1(new_n820), .B2(KEYINPUT55), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n821), .B1(KEYINPUT55), .B2(new_n820), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n333), .A2(new_n822), .ZN(new_n823));
  OAI22_X1  g622(.A1(new_n315), .A2(new_n316), .B1(new_n318), .B2(new_n319), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n308), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n332), .A2(new_n356), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n251), .B1(new_n823), .B2(new_n826), .ZN(new_n827));
  AOI22_X1  g626(.A1(new_n330), .A2(new_n331), .B1(new_n308), .B2(new_n824), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n822), .A2(new_n251), .A3(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n688), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n813), .B1(new_n815), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n531), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(G113gat), .B1(new_n835), .B2(new_n333), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n832), .A2(new_n419), .A3(new_n599), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n837), .A2(new_n431), .A3(new_n814), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n836), .A2(new_n838), .ZN(G1340gat));
  AOI21_X1  g638(.A(G120gat), .B1(new_n835), .B2(new_n356), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n837), .A2(new_n432), .A3(new_n357), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n840), .A2(new_n841), .ZN(G1341gat));
  OAI21_X1  g641(.A(G127gat), .B1(new_n837), .B2(new_n688), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n689), .A2(new_n422), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n843), .B1(new_n834), .B2(new_n844), .ZN(G1342gat));
  NAND4_X1  g644(.A1(new_n832), .A2(new_n424), .A3(new_n833), .A4(new_n251), .ZN(new_n846));
  XOR2_X1   g645(.A(new_n846), .B(KEYINPUT56), .Z(new_n847));
  OAI21_X1  g646(.A(G134gat), .B1(new_n837), .B2(new_n252), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(G1343gat));
  NOR2_X1   g648(.A1(new_n726), .A2(new_n813), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(KEYINPUT121), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n419), .B1(new_n815), .B2(new_n831), .ZN(new_n852));
  XNOR2_X1  g651(.A(KEYINPUT122), .B(KEYINPUT57), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT123), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n826), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n828), .A2(KEYINPUT123), .A3(new_n356), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n251), .B1(new_n860), .B2(new_n823), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n688), .B1(new_n861), .B2(new_n830), .ZN(new_n862));
  AOI211_X1 g661(.A(new_n856), .B(new_n419), .C1(new_n815), .C2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n851), .B1(new_n855), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(G141gat), .B1(new_n864), .B2(new_n814), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n852), .A2(new_n850), .ZN(new_n866));
  OR3_X1    g665(.A1(new_n866), .A2(G141gat), .A3(new_n814), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(KEYINPUT58), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT58), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n865), .A2(new_n870), .A3(new_n867), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n871), .ZN(G1344gat));
  INV_X1    g671(.A(new_n866), .ZN(new_n873));
  INV_X1    g672(.A(G148gat), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n873), .A2(new_n874), .A3(new_n356), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n876));
  OAI21_X1  g675(.A(KEYINPUT124), .B1(new_n861), .B2(new_n830), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT124), .ZN(new_n878));
  AOI22_X1  g677(.A1(new_n858), .A2(new_n859), .B1(new_n333), .B2(new_n822), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n878), .B(new_n829), .C1(new_n879), .C2(new_n251), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n689), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n815), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n663), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n883), .A2(new_n856), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n852), .A2(new_n854), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n356), .B(new_n851), .C1(new_n884), .C2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n876), .B1(new_n887), .B2(G148gat), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n864), .A2(new_n357), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n889), .A2(KEYINPUT59), .A3(new_n874), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n875), .B1(new_n888), .B2(new_n890), .ZN(G1345gat));
  OAI21_X1  g690(.A(G155gat), .B1(new_n864), .B2(new_n688), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n873), .A2(new_n364), .A3(new_n689), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(G1346gat));
  OAI21_X1  g693(.A(G162gat), .B1(new_n864), .B2(new_n252), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n873), .A2(new_n365), .A3(new_n251), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(G1347gat));
  NAND2_X1  g696(.A1(new_n815), .A2(new_n831), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n607), .A2(new_n669), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n900), .A2(new_n531), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(G169gat), .B1(new_n903), .B2(new_n333), .ZN(new_n904));
  AOI211_X1 g703(.A(new_n600), .B(new_n900), .C1(new_n815), .C2(new_n831), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n333), .A2(G169gat), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(G1348gat));
  INV_X1    g706(.A(G176gat), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n903), .A2(new_n908), .A3(new_n356), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n905), .A2(new_n356), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n910), .B2(new_n908), .ZN(G1349gat));
  AOI211_X1 g710(.A(new_n688), .B(new_n902), .C1(new_n492), .C2(new_n491), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n466), .B1(new_n905), .B2(new_n689), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  XOR2_X1   g713(.A(KEYINPUT125), .B(KEYINPUT60), .Z(new_n915));
  XNOR2_X1  g714(.A(new_n914), .B(new_n915), .ZN(G1350gat));
  AOI21_X1  g715(.A(new_n457), .B1(new_n905), .B2(new_n251), .ZN(new_n917));
  XOR2_X1   g716(.A(new_n917), .B(KEYINPUT61), .Z(new_n918));
  NAND3_X1  g717(.A1(new_n903), .A2(new_n457), .A3(new_n251), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(G1351gat));
  AOI22_X1  g719(.A1(new_n883), .A2(new_n856), .B1(new_n852), .B2(new_n854), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n726), .A2(new_n900), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n333), .A2(G197gat), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n921), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n927));
  INV_X1    g726(.A(new_n852), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n928), .A2(new_n923), .ZN(new_n929));
  AOI21_X1  g728(.A(G197gat), .B1(new_n929), .B2(new_n333), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n926), .A2(new_n927), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(KEYINPUT126), .B1(new_n925), .B2(new_n930), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1352gat));
  NOR4_X1   g733(.A1(new_n928), .A2(G204gat), .A3(new_n357), .A4(new_n923), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT62), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n921), .A2(new_n357), .A3(new_n923), .ZN(new_n937));
  INV_X1    g736(.A(G204gat), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(G1353gat));
  NAND3_X1  g738(.A1(new_n929), .A2(new_n380), .A3(new_n689), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT63), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n883), .A2(new_n856), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n923), .B1(new_n942), .B2(new_n885), .ZN(new_n943));
  AOI211_X1 g742(.A(new_n941), .B(new_n380), .C1(new_n943), .C2(new_n689), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n689), .B(new_n922), .C1(new_n884), .C2(new_n886), .ZN(new_n945));
  AOI21_X1  g744(.A(KEYINPUT63), .B1(new_n945), .B2(G211gat), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n940), .B1(new_n944), .B2(new_n946), .ZN(G1354gat));
  AOI21_X1  g746(.A(G218gat), .B1(new_n929), .B2(new_n251), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT127), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n943), .B(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n252), .B1(new_n381), .B2(new_n382), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(G1355gat));
endmodule


