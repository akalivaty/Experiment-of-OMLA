//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 0 1 1 1 1 1 0 1 0 1 0 1 0 1 0 0 1 1 1 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308;
  OR3_X1    g0000(.A1(KEYINPUT64), .A2(G58), .A3(G68), .ZN(new_n201));
  OAI21_X1  g0001(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n202));
  AOI211_X1 g0002(.A(G50), .B(G77), .C1(new_n201), .C2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n206));
  INV_X1    g0006(.A(G68), .ZN(new_n207));
  INV_X1    g0007(.A(G238), .ZN(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n206), .B1(new_n207), .B2(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n205), .B1(new_n211), .B2(new_n214), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n215), .A2(KEYINPUT1), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n201), .A2(new_n202), .ZN(new_n217));
  INV_X1    g0017(.A(G50), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n205), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT0), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n216), .A2(new_n223), .A3(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n215), .ZN(G361));
  XOR2_X1   g0028(.A(G250), .B(G257), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT65), .ZN(new_n230));
  XOR2_X1   g0030(.A(G264), .B(G270), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n232), .B(new_n236), .Z(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XOR2_X1   g0038(.A(G107), .B(G116), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  INV_X1    g0044(.A(G1), .ZN(new_n245));
  INV_X1    g0045(.A(G41), .ZN(new_n246));
  OAI211_X1 g0046(.A(new_n245), .B(G45), .C1(new_n246), .C2(KEYINPUT5), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT78), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G45), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n250), .A2(G1), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT5), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G41), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n251), .A2(KEYINPUT78), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n246), .A2(KEYINPUT5), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n249), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G1), .A3(G13), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n256), .A2(G270), .A3(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  OAI211_X1 g0061(.A(G264), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G1698), .ZN(new_n263));
  OAI211_X1 g0063(.A(G257), .B(new_n263), .C1(new_n260), .C2(new_n261), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT3), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(G303), .A3(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n262), .A2(new_n264), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n220), .B1(G33), .B2(G41), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n247), .A2(new_n248), .B1(KEYINPUT5), .B2(new_n246), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n258), .A2(G274), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n273), .A2(new_n274), .A3(new_n254), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n259), .A2(new_n272), .A3(G179), .A4(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G283), .ZN(new_n278));
  INV_X1    g0078(.A(G97), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n278), .B(new_n221), .C1(G33), .C2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n220), .ZN(new_n282));
  INV_X1    g0082(.A(G116), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G20), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n280), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT20), .ZN(new_n286));
  XNOR2_X1  g0086(.A(new_n285), .B(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n245), .A2(G13), .A3(G20), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n245), .A2(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NOR3_X1   g0090(.A1(new_n290), .A2(new_n283), .A3(new_n282), .ZN(new_n291));
  INV_X1    g0091(.A(new_n288), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n291), .B1(new_n283), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n287), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n277), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G169), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n296), .B1(new_n287), .B2(new_n293), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n259), .A2(new_n272), .A3(new_n275), .ZN(new_n298));
  AOI21_X1  g0098(.A(KEYINPUT80), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT21), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n295), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n298), .A2(G200), .ZN(new_n302));
  INV_X1    g0102(.A(G190), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  NOR3_X1   g0104(.A1(new_n302), .A2(new_n304), .A3(new_n294), .ZN(new_n305));
  AOI211_X1 g0105(.A(KEYINPUT80), .B(KEYINPUT21), .C1(new_n297), .C2(new_n298), .ZN(new_n306));
  NOR3_X1   g0106(.A1(new_n301), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT70), .ZN(new_n308));
  AOI21_X1  g0108(.A(G1698), .B1(new_n267), .B2(new_n268), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G222), .ZN(new_n310));
  INV_X1    g0110(.A(G77), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT3), .B(G33), .ZN(new_n312));
  INV_X1    g0112(.A(G223), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(G1698), .ZN(new_n314));
  OAI221_X1 g0114(.A(new_n310), .B1(new_n311), .B2(new_n312), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n271), .ZN(new_n316));
  OR2_X1    g0116(.A1(KEYINPUT66), .A2(G45), .ZN(new_n317));
  NAND2_X1  g0117(.A1(KEYINPUT66), .A2(G45), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n317), .A2(new_n246), .A3(new_n318), .ZN(new_n319));
  AND3_X1   g0119(.A1(new_n274), .A2(new_n245), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(G1), .B1(new_n246), .B2(new_n250), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n271), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n320), .B1(G226), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n316), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n308), .B1(new_n324), .B2(new_n303), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n316), .A2(new_n323), .A3(KEYINPUT70), .A4(G190), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n325), .A2(new_n326), .B1(G200), .B2(new_n324), .ZN(new_n327));
  INV_X1    g0127(.A(new_n282), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n221), .B1(new_n217), .B2(new_n218), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n329), .B(KEYINPUT68), .ZN(new_n330));
  NOR2_X1   g0130(.A1(KEYINPUT8), .A2(G58), .ZN(new_n331));
  XNOR2_X1  g0131(.A(KEYINPUT67), .B(G58), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n331), .B1(new_n333), .B2(KEYINPUT8), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n221), .A2(G33), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(G20), .A2(G33), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n334), .A2(new_n336), .B1(G150), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n328), .B1(new_n330), .B2(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n288), .A2(G50), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n282), .B1(new_n245), .B2(G20), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n340), .B1(new_n341), .B2(G50), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT9), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NOR3_X1   g0146(.A1(new_n339), .A2(KEYINPUT9), .A3(new_n343), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n327), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n348), .B(KEYINPUT10), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n274), .A2(new_n245), .A3(new_n319), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n322), .A2(G238), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n309), .A2(G226), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G33), .A2(G97), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n312), .A2(G232), .A3(G1698), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n271), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT13), .ZN(new_n358));
  AND3_X1   g0158(.A1(new_n352), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n358), .B1(new_n352), .B2(new_n357), .ZN(new_n360));
  OAI21_X1  g0160(.A(G169), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT14), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT14), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n363), .B(G169), .C1(new_n359), .C2(new_n360), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT71), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n352), .A2(new_n357), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n365), .B1(new_n366), .B2(KEYINPUT13), .ZN(new_n367));
  INV_X1    g0167(.A(new_n360), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n352), .A2(new_n357), .A3(KEYINPUT71), .A4(new_n358), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n367), .A2(new_n368), .A3(G179), .A4(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n362), .A2(new_n364), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n341), .A2(G68), .ZN(new_n372));
  XNOR2_X1  g0172(.A(new_n372), .B(KEYINPUT72), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n337), .A2(G50), .B1(G20), .B2(new_n207), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n311), .B2(new_n335), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n375), .A2(new_n282), .ZN(new_n376));
  OR2_X1    g0176(.A1(new_n376), .A2(KEYINPUT11), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n292), .A2(new_n207), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n378), .B(KEYINPUT12), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n376), .A2(KEYINPUT11), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n373), .A2(new_n377), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n371), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n367), .A2(new_n368), .A3(G190), .A4(new_n369), .ZN(new_n384));
  OAI21_X1  g0184(.A(G200), .B1(new_n359), .B2(new_n360), .ZN(new_n385));
  INV_X1    g0185(.A(new_n381), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n383), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n324), .A2(new_n296), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(G179), .B2(new_n324), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n391), .A2(new_n344), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n320), .B1(G244), .B2(new_n322), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n312), .A2(G232), .A3(new_n263), .ZN(new_n395));
  INV_X1    g0195(.A(G107), .ZN(new_n396));
  OAI221_X1 g0196(.A(new_n395), .B1(new_n396), .B2(new_n312), .C1(new_n314), .C2(new_n208), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n271), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G200), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n292), .A2(new_n311), .ZN(new_n401));
  INV_X1    g0201(.A(new_n341), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n401), .B1(new_n402), .B2(new_n311), .ZN(new_n403));
  XOR2_X1   g0203(.A(KEYINPUT8), .B(G58), .Z(new_n404));
  AOI22_X1  g0204(.A1(new_n404), .A2(new_n337), .B1(G20), .B2(G77), .ZN(new_n405));
  XNOR2_X1  g0205(.A(KEYINPUT15), .B(G87), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n407), .A2(KEYINPUT69), .A3(new_n336), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT69), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n406), .B2(new_n335), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n405), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n403), .B1(new_n282), .B2(new_n411), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n400), .B(new_n412), .C1(new_n303), .C2(new_n399), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n412), .B1(new_n399), .B2(new_n296), .ZN(new_n414));
  INV_X1    g0214(.A(G179), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n394), .A2(new_n415), .A3(new_n398), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n349), .A2(new_n389), .A3(new_n393), .A4(new_n418), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n334), .A2(new_n292), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n420), .B1(new_n334), .B2(new_n402), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n201), .B(new_n202), .C1(new_n332), .C2(new_n207), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n422), .A2(G20), .B1(G159), .B2(new_n337), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n260), .A2(new_n261), .ZN(new_n424));
  AOI21_X1  g0224(.A(KEYINPUT7), .B1(new_n424), .B2(new_n221), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n267), .A2(KEYINPUT7), .A3(new_n221), .A4(new_n268), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(G68), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n423), .A2(KEYINPUT16), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n282), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n267), .A2(new_n221), .A3(new_n268), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT7), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT73), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n433), .A2(new_n434), .A3(new_n426), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n427), .A2(KEYINPUT73), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(G68), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n423), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT16), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT74), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n430), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(KEYINPUT16), .B1(new_n437), .B2(new_n423), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(KEYINPUT74), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n421), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n322), .A2(G232), .ZN(new_n446));
  MUX2_X1   g0246(.A(G223), .B(G226), .S(G1698), .Z(new_n447));
  AOI22_X1  g0247(.A1(new_n447), .A2(new_n312), .B1(G33), .B2(G87), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n350), .B(new_n446), .C1(new_n448), .C2(new_n258), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(G169), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(new_n415), .B2(new_n449), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(KEYINPUT18), .B1(new_n445), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n421), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n448), .A2(new_n258), .ZN(new_n455));
  INV_X1    g0255(.A(new_n446), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n457), .A2(KEYINPUT75), .A3(new_n303), .A4(new_n350), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT75), .ZN(new_n459));
  INV_X1    g0259(.A(G200), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n459), .B1(new_n449), .B2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n449), .A2(G190), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n458), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n444), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n282), .B(new_n429), .C1(new_n443), .C2(KEYINPUT74), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n454), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT17), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n454), .B1(new_n464), .B2(new_n465), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT18), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n469), .A2(new_n470), .A3(new_n451), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n442), .A2(new_n444), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n472), .A2(KEYINPUT17), .A3(new_n454), .A4(new_n463), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n453), .A2(new_n468), .A3(new_n471), .A4(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n419), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n271), .B1(new_n273), .B2(new_n254), .ZN(new_n476));
  OAI211_X1 g0276(.A(G257), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n477));
  OAI211_X1 g0277(.A(G250), .B(new_n263), .C1(new_n260), .C2(new_n261), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G33), .A2(G294), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n476), .A2(G264), .B1(new_n271), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n275), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n296), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n481), .A2(new_n415), .A3(new_n275), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT23), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n486), .B1(new_n221), .B2(G107), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n396), .A2(KEYINPUT23), .A3(G20), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n266), .A2(new_n283), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n487), .A2(new_n488), .B1(new_n489), .B2(new_n221), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n221), .B(G87), .C1(new_n260), .C2(new_n261), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(KEYINPUT82), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT82), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n312), .A2(new_n493), .A3(new_n221), .A4(G87), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT81), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(KEYINPUT22), .ZN(new_n496));
  AND3_X1   g0296(.A1(new_n492), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n496), .B1(new_n492), .B2(new_n494), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n490), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT24), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT24), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n501), .B(new_n490), .C1(new_n497), .C2(new_n498), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n282), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n328), .A2(KEYINPUT77), .A3(new_n288), .A4(new_n289), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT77), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n506), .B1(new_n290), .B2(new_n282), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n505), .A2(new_n507), .A3(G107), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n288), .A2(G107), .ZN(new_n509));
  XNOR2_X1  g0309(.A(new_n509), .B(KEYINPUT25), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n485), .B1(new_n504), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n328), .B1(new_n500), .B2(new_n502), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n256), .A2(G264), .A3(new_n258), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n480), .A2(new_n271), .ZN(new_n516));
  AND4_X1   g0316(.A1(new_n303), .A2(new_n515), .A3(new_n275), .A4(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n517), .B1(new_n460), .B2(new_n482), .ZN(new_n518));
  NOR3_X1   g0318(.A1(new_n514), .A2(new_n518), .A3(new_n511), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n513), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(G250), .B1(new_n250), .B2(G1), .ZN(new_n521));
  OAI21_X1  g0321(.A(KEYINPUT79), .B1(new_n271), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n210), .B1(new_n245), .B2(G45), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT79), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(new_n258), .A3(new_n524), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n522), .A2(new_n525), .B1(new_n274), .B2(new_n251), .ZN(new_n526));
  OAI211_X1 g0326(.A(G244), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n527));
  OAI211_X1 g0327(.A(G238), .B(new_n263), .C1(new_n260), .C2(new_n261), .ZN(new_n528));
  INV_X1    g0328(.A(new_n489), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n271), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(G200), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT19), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n221), .B1(new_n354), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(G97), .A2(G107), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n209), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n221), .B(G68), .C1(new_n260), .C2(new_n261), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n534), .B1(new_n335), .B2(new_n279), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n541), .A2(new_n282), .B1(new_n292), .B2(new_n406), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n505), .A2(new_n507), .A3(G87), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n526), .A2(new_n531), .A3(G190), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n533), .A2(new_n542), .A3(new_n543), .A4(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n532), .A2(new_n296), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n505), .A2(new_n507), .A3(new_n407), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n526), .A2(new_n531), .A3(new_n415), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n546), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n435), .A2(G107), .A3(new_n436), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT76), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT6), .ZN(new_n555));
  AND2_X1   g0355(.A1(G97), .A2(G107), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n555), .B1(new_n556), .B2(new_n536), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n396), .A2(KEYINPUT6), .A3(G97), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n221), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n337), .A2(G77), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n554), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n558), .ZN(new_n563));
  XNOR2_X1  g0363(.A(G97), .B(G107), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n563), .B1(new_n555), .B2(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(KEYINPUT76), .B(new_n560), .C1(new_n565), .C2(new_n221), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n553), .A2(new_n562), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n282), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n505), .A2(new_n507), .A3(G97), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n292), .A2(new_n279), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n249), .A2(new_n254), .A3(new_n255), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n476), .A2(G257), .B1(new_n574), .B2(new_n274), .ZN(new_n575));
  OAI211_X1 g0375(.A(G244), .B(new_n263), .C1(new_n260), .C2(new_n261), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT4), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n312), .A2(KEYINPUT4), .A3(G244), .A4(new_n263), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n312), .A2(G250), .A3(G1698), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n578), .A2(new_n579), .A3(new_n278), .A4(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n271), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n575), .A2(new_n415), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(G169), .B1(new_n575), .B2(new_n582), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n573), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n571), .B1(new_n567), .B2(new_n282), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n476), .A2(G257), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n582), .A2(new_n275), .A3(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n589), .A2(G190), .ZN(new_n590));
  AOI21_X1  g0390(.A(G200), .B1(new_n575), .B2(new_n582), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n587), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AND3_X1   g0392(.A1(new_n552), .A2(new_n586), .A3(new_n592), .ZN(new_n593));
  AND4_X1   g0393(.A1(new_n307), .A2(new_n475), .A3(new_n520), .A4(new_n593), .ZN(G372));
  INV_X1    g0394(.A(new_n550), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n542), .A2(KEYINPUT83), .A3(new_n543), .ZN(new_n596));
  AOI21_X1  g0396(.A(KEYINPUT83), .B1(new_n542), .B2(new_n543), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n533), .B(new_n544), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n586), .A2(new_n592), .A3(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n599), .A2(new_n519), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n484), .B(new_n483), .C1(new_n514), .C2(new_n511), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n299), .A2(new_n300), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n294), .A2(new_n298), .A3(G169), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT80), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(KEYINPUT21), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n601), .A2(new_n602), .A3(new_n295), .A4(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n595), .B1(new_n600), .B2(new_n607), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n581), .A2(new_n271), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n256), .A2(new_n258), .ZN(new_n610));
  INV_X1    g0410(.A(G257), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n275), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NOR3_X1   g0412(.A1(new_n609), .A2(new_n612), .A3(G179), .ZN(new_n613));
  NOR3_X1   g0413(.A1(new_n587), .A2(new_n613), .A3(new_n584), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT84), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n614), .A2(new_n552), .A3(new_n615), .A4(KEYINPUT26), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n613), .A2(new_n584), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n617), .A2(new_n573), .A3(new_n598), .A4(new_n550), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT26), .ZN(new_n619));
  AOI21_X1  g0419(.A(KEYINPUT84), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NOR3_X1   g0420(.A1(new_n586), .A2(new_n551), .A3(new_n619), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n616), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n608), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n475), .A2(new_n623), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n445), .A2(KEYINPUT18), .A3(new_n452), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n470), .B1(new_n469), .B2(new_n451), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n417), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n383), .B1(new_n387), .B2(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n468), .A2(new_n473), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n627), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n392), .B1(new_n632), .B2(new_n349), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n624), .A2(new_n633), .ZN(G369));
  NAND3_X1  g0434(.A1(new_n606), .A2(new_n602), .A3(new_n295), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n245), .A2(new_n221), .A3(G13), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n636), .A2(KEYINPUT27), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(KEYINPUT27), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(G213), .A3(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(G343), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n635), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n520), .ZN(new_n644));
  XOR2_X1   g0444(.A(new_n641), .B(KEYINPUT85), .Z(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n644), .B1(new_n601), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT86), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n647), .B(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n641), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n294), .ZN(new_n651));
  MUX2_X1   g0451(.A(new_n635), .B(new_n307), .S(new_n651), .Z(new_n652));
  AND2_X1   g0452(.A1(new_n652), .A2(G330), .ZN(new_n653));
  INV_X1    g0453(.A(new_n520), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n641), .B1(new_n504), .B2(new_n512), .ZN(new_n655));
  OAI22_X1  g0455(.A1(new_n654), .A2(new_n655), .B1(new_n601), .B2(new_n641), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n649), .A2(new_n657), .ZN(G399));
  INV_X1    g0458(.A(new_n224), .ZN(new_n659));
  OR3_X1    g0459(.A1(new_n659), .A2(KEYINPUT87), .A3(G41), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT87), .B1(new_n659), .B2(G41), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n537), .A2(G116), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(G1), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n219), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n664), .B(KEYINPUT88), .C1(new_n665), .C2(new_n662), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(KEYINPUT88), .B2(new_n664), .ZN(new_n667));
  XOR2_X1   g0467(.A(new_n667), .B(KEYINPUT28), .Z(new_n668));
  AND2_X1   g0468(.A1(new_n598), .A2(new_n550), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n669), .A2(KEYINPUT26), .A3(new_n614), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n619), .B1(new_n586), .B2(new_n551), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(KEYINPUT90), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(KEYINPUT90), .B2(new_n670), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n586), .A2(new_n592), .ZN(new_n674));
  OR3_X1    g0474(.A1(new_n514), .A2(new_n518), .A3(new_n511), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(new_n675), .A3(new_n598), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n513), .A2(new_n635), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n550), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  OAI211_X1 g0478(.A(KEYINPUT29), .B(new_n641), .C1(new_n673), .C2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n646), .B1(new_n608), .B2(new_n622), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n679), .B1(KEYINPUT29), .B2(new_n680), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n520), .A2(new_n307), .A3(new_n593), .A4(new_n645), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n489), .B1(new_n309), .B2(G238), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n258), .B1(new_n683), .B2(new_n527), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n258), .A2(G274), .A3(new_n251), .ZN(new_n685));
  INV_X1    g0485(.A(new_n525), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n524), .B1(new_n523), .B2(new_n258), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n685), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n689), .A2(new_n575), .A3(new_n481), .A4(new_n582), .ZN(new_n690));
  OAI21_X1  g0490(.A(KEYINPUT30), .B1(new_n690), .B2(new_n276), .ZN(new_n691));
  INV_X1    g0491(.A(new_n589), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT30), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n515), .A2(new_n526), .A3(new_n516), .A4(new_n531), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n692), .A2(new_n277), .A3(new_n693), .A4(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n691), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT89), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n684), .B2(new_n688), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n526), .A2(new_n531), .A3(KEYINPUT89), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(G179), .B1(new_n481), .B2(new_n275), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n701), .A2(new_n298), .A3(new_n589), .A4(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n641), .B1(new_n697), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n298), .B1(new_n609), .B2(new_n612), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n699), .A2(new_n700), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AOI22_X1  g0507(.A1(new_n691), .A2(new_n696), .B1(new_n707), .B2(new_n702), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n646), .A2(KEYINPUT31), .ZN(new_n709));
  OAI221_X1 g0509(.A(new_n682), .B1(KEYINPUT31), .B2(new_n704), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G330), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n681), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n668), .B1(new_n713), .B2(G1), .ZN(G364));
  INV_X1    g0514(.A(new_n662), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n221), .A2(G13), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT91), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n245), .B1(new_n717), .B2(G45), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n653), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(G330), .B2(new_n652), .ZN(new_n722));
  INV_X1    g0522(.A(new_n720), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n296), .A2(KEYINPUT95), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n221), .B1(KEYINPUT95), .B2(new_n296), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n220), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(G179), .A2(G200), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(G20), .A3(new_n303), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  OR2_X1    g0531(.A1(new_n731), .A2(KEYINPUT97), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(KEYINPUT97), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(G159), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g0536(.A(new_n736), .B(KEYINPUT32), .ZN(new_n737));
  NOR4_X1   g0537(.A1(new_n221), .A2(new_n460), .A3(G179), .A4(G190), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n396), .ZN(new_n740));
  NAND2_X1  g0540(.A1(G20), .A2(G179), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G200), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n303), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n221), .B1(new_n729), .B2(G190), .ZN(new_n746));
  OAI22_X1  g0546(.A1(new_n745), .A2(new_n218), .B1(new_n746), .B2(new_n279), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n743), .A2(G190), .ZN(new_n748));
  AOI211_X1 g0548(.A(new_n740), .B(new_n747), .C1(G68), .C2(new_n748), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n741), .A2(new_n303), .A3(G200), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n312), .B1(new_n751), .B2(new_n332), .ZN(new_n752));
  NOR4_X1   g0552(.A1(new_n221), .A2(new_n303), .A3(new_n460), .A4(G179), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n209), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G190), .A2(G200), .ZN(new_n756));
  AND3_X1   g0556(.A1(new_n742), .A2(KEYINPUT96), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(KEYINPUT96), .B1(new_n742), .B2(new_n756), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI211_X1 g0560(.A(new_n752), .B(new_n755), .C1(G77), .C2(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n737), .A2(new_n749), .A3(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G326), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n745), .A2(new_n763), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n312), .B(new_n764), .C1(G322), .C2(new_n750), .ZN(new_n765));
  INV_X1    g0565(.A(new_n748), .ZN(new_n766));
  XOR2_X1   g0566(.A(KEYINPUT33), .B(G317), .Z(new_n767));
  INV_X1    g0567(.A(G283), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n766), .A2(new_n767), .B1(new_n768), .B2(new_n739), .ZN(new_n769));
  INV_X1    g0569(.A(G303), .ZN(new_n770));
  INV_X1    g0570(.A(G294), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n754), .A2(new_n770), .B1(new_n771), .B2(new_n746), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n760), .A2(G311), .ZN(new_n774));
  INV_X1    g0574(.A(new_n734), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G329), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n765), .A2(new_n773), .A3(new_n774), .A4(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n728), .B1(new_n762), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G13), .A2(G33), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n727), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n424), .A2(new_n224), .ZN(new_n783));
  XOR2_X1   g0583(.A(new_n783), .B(KEYINPUT94), .Z(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n317), .A2(new_n318), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n785), .B1(new_n219), .B2(new_n787), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n243), .A2(new_n250), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n659), .A2(new_n424), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT92), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G355), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(G116), .B2(new_n224), .ZN(new_n793));
  INV_X1    g0593(.A(KEYINPUT93), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n788), .A2(new_n789), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n723), .B(new_n778), .C1(new_n782), .C2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n781), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n798), .B1(new_n652), .B2(new_n799), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n722), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(G396));
  NAND2_X1  g0602(.A1(new_n728), .A2(new_n780), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n720), .B1(G77), .B2(new_n803), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n768), .A2(new_n766), .B1(new_n745), .B2(new_n770), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(new_n760), .B2(G116), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT98), .Z(new_n807));
  OAI21_X1  g0607(.A(new_n424), .B1(new_n751), .B2(new_n771), .ZN(new_n808));
  INV_X1    g0608(.A(new_n746), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n808), .B1(G97), .B2(new_n809), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n753), .A2(G107), .B1(new_n738), .B2(G87), .ZN(new_n811));
  INV_X1    g0611(.A(G311), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n810), .B(new_n811), .C1(new_n812), .C2(new_n734), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n744), .A2(G137), .B1(G143), .B2(new_n750), .ZN(new_n814));
  INV_X1    g0614(.A(G150), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n814), .B1(new_n815), .B2(new_n766), .C1(new_n735), .C2(new_n759), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(KEYINPUT34), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n312), .B1(new_n746), .B2(new_n332), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n754), .A2(new_n218), .B1(new_n739), .B2(new_n207), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n819), .B(new_n820), .C1(new_n775), .C2(G132), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT34), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n821), .B1(new_n822), .B2(new_n816), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n807), .A2(new_n813), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n804), .B1(new_n824), .B2(new_n727), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n413), .B1(new_n412), .B2(new_n641), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n417), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n628), .A2(new_n641), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n825), .B1(new_n830), .B2(new_n780), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n680), .A2(new_n830), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n680), .A2(new_n830), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n711), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n723), .ZN(new_n836));
  NOR3_X1   g0636(.A1(new_n833), .A2(new_n711), .A3(new_n834), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n831), .B1(new_n836), .B2(new_n837), .ZN(G384));
  NOR2_X1   g0638(.A1(new_n717), .A2(new_n245), .ZN(new_n839));
  INV_X1    g0639(.A(G330), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT31), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n641), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(KEYINPUT101), .B1(new_n708), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n589), .A2(new_n694), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n693), .B1(new_n845), .B2(new_n277), .ZN(new_n846));
  NOR4_X1   g0646(.A1(new_n589), .A2(new_n694), .A3(new_n276), .A4(KEYINPUT30), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n703), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT101), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n848), .A2(new_n849), .A3(new_n842), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n844), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(KEYINPUT100), .B1(new_n704), .B2(KEYINPUT31), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT100), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n853), .B(new_n841), .C1(new_n708), .C2(new_n641), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n682), .A2(new_n851), .A3(new_n852), .A4(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n381), .A2(new_n650), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n382), .A2(new_n387), .A3(new_n856), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n381), .B(new_n650), .C1(new_n388), .C2(new_n371), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n829), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(KEYINPUT102), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT16), .B1(new_n423), .B2(new_n428), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n430), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n863), .A2(new_n421), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n864), .A2(new_n639), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n474), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n469), .A2(new_n451), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n469), .A2(new_n640), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT37), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n867), .A2(new_n868), .A3(new_n869), .A4(new_n466), .ZN(new_n870));
  OAI22_X1  g0670(.A1(new_n863), .A2(new_n421), .B1(new_n451), .B2(new_n640), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n466), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(KEYINPUT37), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n866), .A2(KEYINPUT38), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n466), .B1(new_n445), .B2(new_n452), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n445), .A2(new_n639), .ZN(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT37), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n870), .A2(new_n878), .B1(new_n474), .B2(new_n877), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n875), .B1(new_n879), .B2(KEYINPUT38), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT102), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n855), .A2(new_n859), .A3(new_n881), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n861), .A2(new_n880), .A3(KEYINPUT40), .A4(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(KEYINPUT103), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n855), .A2(new_n881), .A3(new_n859), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n881), .B1(new_n855), .B2(new_n859), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT40), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT38), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n878), .A2(new_n870), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n868), .B1(new_n627), .B2(new_n630), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n888), .B1(new_n892), .B2(new_n875), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT103), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n887), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n866), .A2(KEYINPUT38), .A3(new_n874), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT38), .B1(new_n866), .B2(new_n874), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n859), .B(new_n855), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n884), .A2(new_n895), .B1(new_n888), .B2(new_n898), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n475), .A2(new_n855), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n840), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n899), .B2(new_n900), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n627), .A2(new_n640), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n857), .A2(new_n858), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n832), .B2(new_n828), .ZN(new_n906));
  INV_X1    g0706(.A(new_n897), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n875), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n903), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT39), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n880), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n907), .A2(KEYINPUT39), .A3(new_n875), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n382), .A2(new_n650), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n909), .A2(new_n914), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n475), .B(new_n679), .C1(KEYINPUT29), .C2(new_n680), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n916), .A2(new_n633), .ZN(new_n917));
  XOR2_X1   g0717(.A(new_n915), .B(new_n917), .Z(new_n918));
  AOI21_X1  g0718(.A(new_n839), .B1(new_n902), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n918), .B2(new_n902), .ZN(new_n920));
  INV_X1    g0720(.A(new_n565), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n921), .A2(KEYINPUT35), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(KEYINPUT35), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n922), .A2(G116), .A3(new_n222), .A4(new_n923), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n924), .B(KEYINPUT36), .Z(new_n925));
  AOI211_X1 g0725(.A(new_n311), .B(new_n665), .C1(G68), .C2(new_n333), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT99), .ZN(new_n927));
  AOI22_X1  g0727(.A1(new_n926), .A2(new_n927), .B1(new_n218), .B2(G68), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n927), .B2(new_n926), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n245), .A2(G13), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n925), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n920), .A2(new_n931), .ZN(G367));
  NOR2_X1   g0732(.A1(new_n232), .A2(new_n785), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n782), .B1(new_n224), .B2(new_n406), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n720), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n424), .B1(new_n751), .B2(new_n770), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(G97), .B2(new_n738), .ZN(new_n937));
  INV_X1    g0737(.A(G317), .ZN(new_n938));
  OAI221_X1 g0738(.A(new_n937), .B1(new_n768), .B2(new_n759), .C1(new_n938), .C2(new_n734), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n753), .A2(G116), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT46), .ZN(new_n941));
  XOR2_X1   g0741(.A(KEYINPUT107), .B(G311), .Z(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n744), .A2(new_n943), .B1(new_n809), .B2(G107), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n941), .B(new_n944), .C1(new_n771), .C2(new_n766), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n312), .B1(new_n751), .B2(new_n815), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(G68), .B2(new_n809), .ZN(new_n947));
  INV_X1    g0747(.A(G137), .ZN(new_n948));
  OAI221_X1 g0748(.A(new_n947), .B1(new_n218), .B2(new_n759), .C1(new_n948), .C2(new_n734), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n744), .A2(G143), .B1(G77), .B2(new_n738), .ZN(new_n950));
  OAI221_X1 g0750(.A(new_n950), .B1(new_n735), .B2(new_n766), .C1(new_n332), .C2(new_n754), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n939), .A2(new_n945), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT47), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n935), .B1(new_n953), .B2(new_n727), .ZN(new_n954));
  OR3_X1    g0754(.A1(new_n596), .A2(new_n597), .A3(new_n641), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n955), .A2(new_n550), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(new_n669), .B2(new_n955), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n781), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n662), .B(KEYINPUT41), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT106), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT44), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n674), .B1(new_n587), .B2(new_n645), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n586), .B2(new_n645), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT105), .Z(new_n965));
  OAI21_X1  g0765(.A(new_n962), .B1(new_n649), .B2(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n647), .B(KEYINPUT86), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n964), .B(KEYINPUT105), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n967), .A2(KEYINPUT44), .A3(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT45), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n967), .B2(new_n968), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n649), .A2(KEYINPUT45), .A3(new_n965), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n966), .A2(new_n969), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n961), .B1(new_n973), .B2(new_n657), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n966), .A2(new_n969), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n971), .A2(new_n972), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n657), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n977), .A2(KEYINPUT106), .A3(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n644), .B1(new_n656), .B2(new_n643), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(new_n653), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n713), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n975), .A2(new_n976), .A3(new_n657), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n974), .A2(new_n979), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n960), .B1(new_n985), .B2(new_n713), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n986), .A2(new_n719), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n586), .B1(new_n968), .B2(new_n601), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n645), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n968), .A2(new_n644), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT42), .ZN(new_n991));
  XOR2_X1   g0791(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n992));
  AND4_X1   g0792(.A1(new_n989), .A2(new_n991), .A3(new_n957), .A4(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n965), .A2(new_n978), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n957), .A2(new_n992), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT43), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n995), .B1(new_n996), .B2(new_n957), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(new_n991), .B2(new_n989), .ZN(new_n998));
  OR3_X1    g0798(.A1(new_n993), .A2(new_n994), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n994), .B1(new_n993), .B2(new_n998), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n959), .B1(new_n987), .B2(new_n1001), .ZN(G387));
  NOR2_X1   g0802(.A1(new_n656), .A2(new_n799), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n663), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n791), .A2(new_n1004), .B1(new_n396), .B2(new_n659), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n236), .A2(new_n786), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT108), .Z(new_n1007));
  OR2_X1    g0807(.A1(new_n1004), .A2(KEYINPUT109), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1004), .A2(KEYINPUT109), .ZN(new_n1009));
  AOI21_X1  g0809(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1011), .A2(KEYINPUT110), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(KEYINPUT110), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n404), .A2(new_n218), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT50), .Z(new_n1015));
  NAND3_X1  g0815(.A1(new_n1012), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n784), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1005), .B1(new_n1007), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n723), .B1(new_n1018), .B2(new_n782), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT111), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n312), .B1(new_n751), .B2(new_n218), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n754), .A2(new_n311), .B1(new_n406), .B2(new_n746), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n1021), .B(new_n1022), .C1(G97), .C2(new_n738), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n744), .A2(KEYINPUT112), .A3(G159), .ZN(new_n1024));
  AOI21_X1  g0824(.A(KEYINPUT112), .B1(new_n744), .B2(G159), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n334), .B2(new_n748), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n775), .A2(G150), .B1(G68), .B2(new_n760), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1023), .A2(new_n1024), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n744), .A2(G322), .B1(G317), .B2(new_n750), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n766), .B2(new_n942), .C1(new_n770), .C2(new_n759), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT48), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n753), .A2(G294), .B1(new_n809), .B2(G283), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT49), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(KEYINPUT113), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n312), .B1(new_n738), .B2(G116), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1037), .B(new_n1038), .C1(new_n763), .C2(new_n734), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1036), .A2(KEYINPUT113), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1028), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n1003), .B(new_n1020), .C1(new_n727), .C2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n719), .B2(new_n981), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n982), .A2(new_n715), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n713), .A2(new_n981), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(G393));
  XNOR2_X1  g0846(.A(new_n973), .B(new_n978), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n985), .B(new_n715), .C1(new_n983), .C2(new_n1047), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n312), .B(new_n740), .C1(new_n775), .C2(G322), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n766), .A2(new_n770), .B1(new_n754), .B2(new_n768), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(G116), .B2(new_n809), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1049), .B(new_n1051), .C1(new_n771), .C2(new_n759), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n744), .A2(G317), .B1(G311), .B2(new_n750), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT52), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n744), .A2(G150), .B1(G159), .B2(new_n750), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT51), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n746), .A2(new_n311), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n754), .A2(new_n207), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n1057), .B(new_n1058), .C1(G50), .C2(new_n748), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n775), .A2(G143), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n760), .A2(new_n404), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n424), .B1(new_n738), .B2(G87), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n1052), .A2(new_n1054), .B1(new_n1056), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n727), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n784), .A2(new_n240), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1066), .B(new_n782), .C1(new_n279), .C2(new_n224), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1065), .A2(new_n720), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n968), .B2(new_n781), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n1047), .B2(new_n719), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1048), .A2(new_n1070), .ZN(G390));
  NAND2_X1  g0871(.A1(new_n911), .A2(new_n912), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n913), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n828), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n680), .B2(new_n830), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1073), .B1(new_n1075), .B2(new_n905), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n641), .B(new_n827), .C1(new_n673), .C2(new_n678), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n828), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n904), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n913), .B1(new_n892), .B2(new_n875), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n1072), .A2(new_n1076), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT114), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n710), .A2(G330), .A3(new_n830), .A4(new_n904), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(KEYINPUT39), .B1(new_n892), .B2(new_n875), .ZN(new_n1085));
  NOR3_X1   g0885(.A1(new_n896), .A2(new_n897), .A3(new_n910), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1076), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1087), .A2(new_n1088), .A3(new_n1083), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(KEYINPUT114), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n855), .A2(new_n859), .A3(G330), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1084), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n719), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1072), .A2(new_n779), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n720), .B1(new_n334), .B2(new_n803), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n396), .A2(new_n766), .B1(new_n745), .B2(new_n768), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n1057), .B(new_n1097), .C1(G68), .C2(new_n738), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n760), .A2(G97), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n775), .A2(G294), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n312), .B(new_n755), .C1(G116), .C2(new_n750), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .A4(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n753), .A2(G150), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n775), .A2(G125), .B1(KEYINPUT53), .B2(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(KEYINPUT54), .B(G143), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n759), .A2(new_n1105), .B1(new_n766), .B2(new_n948), .ZN(new_n1106));
  OR2_X1    g0906(.A1(new_n1106), .A2(KEYINPUT116), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(KEYINPUT116), .ZN(new_n1108));
  OR2_X1    g0908(.A1(new_n1103), .A2(KEYINPUT53), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1104), .A2(new_n1107), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n424), .B1(new_n738), .B2(G50), .ZN(new_n1111));
  OR2_X1    g0911(.A1(new_n1111), .A2(KEYINPUT117), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(KEYINPUT117), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n744), .A2(G128), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n809), .A2(G159), .B1(new_n750), .B2(G132), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1102), .B1(new_n1110), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1096), .B1(new_n1117), .B2(new_n727), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1095), .A2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT118), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n1077), .A2(new_n828), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n855), .A2(G330), .A3(new_n830), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n905), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1121), .A2(new_n1083), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT115), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1121), .A2(new_n1123), .A3(KEYINPUT115), .A4(new_n1083), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1075), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n905), .B1(new_n711), .B2(new_n829), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n1091), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n1126), .A2(new_n1127), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n475), .A2(G330), .A3(new_n855), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n917), .A2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n715), .B1(new_n1093), .B2(new_n1134), .ZN(new_n1135));
  AND4_X1   g0935(.A1(new_n1082), .A2(new_n1087), .A3(new_n1088), .A4(new_n1083), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1082), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1092), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1136), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1131), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1133), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1094), .B(new_n1120), .C1(new_n1135), .C2(new_n1143), .ZN(G378));
  NAND2_X1  g0944(.A1(new_n884), .A2(new_n895), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n840), .B1(new_n898), .B2(new_n888), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n1145), .A2(new_n915), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n915), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n349), .A2(new_n393), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n344), .A2(new_n639), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1150), .B(KEYINPUT55), .ZN(new_n1151));
  OR2_X1    g0951(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  XOR2_X1   g0952(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n1153));
  NAND2_X1  g0953(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1153), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NOR3_X1   g0958(.A1(new_n1147), .A2(new_n1148), .A3(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n883), .A2(KEYINPUT103), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n894), .B1(new_n887), .B2(new_n893), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1146), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n915), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1145), .A2(new_n915), .A3(new_n1146), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1157), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1159), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1141), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1168));
  AOI21_X1  g0968(.A(KEYINPUT57), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1158), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1164), .A2(new_n1165), .A3(new_n1157), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1170), .A2(KEYINPUT57), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1133), .B1(new_n1093), .B2(new_n1134), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n715), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1169), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1170), .A2(new_n719), .A3(new_n1171), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n720), .B1(G50), .B2(new_n803), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n312), .A2(G41), .ZN(new_n1178));
  AOI211_X1 g0978(.A(G50), .B(new_n1178), .C1(new_n266), .C2(new_n246), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n739), .A2(new_n332), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n766), .A2(new_n279), .B1(new_n754), .B2(new_n311), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1180), .B(new_n1181), .C1(G116), .C2(new_n744), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1178), .B1(new_n207), .B2(new_n746), .C1(new_n396), .C2(new_n751), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n775), .B2(G283), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1182), .B(new_n1184), .C1(new_n406), .C2(new_n759), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT58), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1179), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  AOI211_X1 g0987(.A(G33), .B(G41), .C1(new_n738), .C2(G159), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(KEYINPUT120), .B(G124), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n748), .A2(G132), .B1(G128), .B2(new_n750), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n754), .B2(new_n1105), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n744), .A2(G125), .B1(new_n809), .B2(G150), .ZN(new_n1192));
  XOR2_X1   g0992(.A(new_n1192), .B(KEYINPUT119), .Z(new_n1193));
  AOI211_X1 g0993(.A(new_n1191), .B(new_n1193), .C1(G137), .C2(new_n760), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT59), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1188), .B1(new_n734), .B2(new_n1189), .C1(new_n1194), .C2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1194), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1197), .A2(KEYINPUT59), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1187), .B1(new_n1186), .B2(new_n1185), .C1(new_n1196), .C2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1177), .B1(new_n1199), .B2(new_n727), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n1157), .B2(new_n780), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1176), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1175), .A2(new_n1203), .ZN(G375));
  NAND2_X1  g1004(.A1(new_n905), .A2(new_n779), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n720), .B1(G68), .B2(new_n803), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n759), .A2(new_n396), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n751), .A2(new_n768), .B1(new_n746), .B2(new_n406), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1207), .B(new_n1208), .C1(new_n775), .C2(G303), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n748), .A2(G116), .B1(new_n753), .B2(G97), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1209), .B(new_n1210), .C1(new_n771), .C2(new_n745), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n312), .B1(new_n738), .B2(G77), .ZN(new_n1212));
  XOR2_X1   g1012(.A(new_n1212), .B(KEYINPUT122), .Z(new_n1213));
  NOR2_X1   g1013(.A1(new_n1211), .A2(new_n1213), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n1214), .A2(KEYINPUT123), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(KEYINPUT123), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n754), .A2(new_n735), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n766), .A2(new_n1105), .B1(new_n218), .B2(new_n746), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1217), .B(new_n1218), .C1(G132), .C2(new_n744), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n760), .A2(G150), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n775), .A2(G128), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n424), .B(new_n1180), .C1(G137), .C2(new_n750), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .A4(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1215), .A2(new_n1216), .A3(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1206), .B1(new_n1224), .B2(new_n727), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1205), .A2(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n1131), .B2(new_n718), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1134), .A2(new_n960), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1228), .B1(new_n1229), .B2(new_n1231), .ZN(G381));
  OR3_X1    g1032(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1233));
  NOR4_X1   g1033(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1094), .A2(new_n1120), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1143), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n662), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1235), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1234), .A2(new_n1238), .A3(new_n1175), .A4(new_n1203), .ZN(G407));
  INV_X1    g1039(.A(G343), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(G213), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1238), .A2(new_n1242), .ZN(new_n1243));
  OAI211_X1 g1043(.A(G407), .B(G213), .C1(G375), .C2(new_n1243), .ZN(G409));
  INV_X1    g1044(.A(G390), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(G387), .A2(new_n1245), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n959), .B(G390), .C1(new_n987), .C2(new_n1001), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(G393), .B(new_n801), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1246), .A2(new_n1247), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(KEYINPUT126), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT126), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1246), .A2(new_n1247), .A3(new_n1252), .A4(new_n1249), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1251), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT125), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1246), .A2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(G387), .A2(KEYINPUT125), .A3(new_n1245), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1256), .A2(new_n1257), .A3(new_n1247), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1248), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1254), .A2(new_n1259), .ZN(new_n1260));
  OAI211_X1 g1060(.A(G378), .B(new_n1203), .C1(new_n1169), .C2(new_n1174), .ZN(new_n1261));
  NOR4_X1   g1061(.A1(new_n1173), .A2(new_n1159), .A3(new_n1166), .A4(new_n960), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1238), .B1(new_n1262), .B2(new_n1202), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1261), .A2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(KEYINPUT60), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n662), .B1(new_n1265), .B2(new_n1230), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1131), .A2(KEYINPUT60), .A3(new_n1133), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(G384), .B(KEYINPUT124), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1268), .A2(new_n1228), .A3(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(G384), .A2(KEYINPUT124), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(new_n1268), .B2(new_n1228), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1270), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1264), .A2(new_n1241), .A3(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT63), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1242), .B1(new_n1261), .B2(new_n1263), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1278), .A2(KEYINPUT63), .A3(new_n1274), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1264), .A2(new_n1241), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1242), .A2(G2897), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1282), .B1(new_n1270), .B2(new_n1273), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1227), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1269), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1285), .B(new_n1281), .C1(new_n1284), .C2(new_n1272), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1283), .A2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT61), .B1(new_n1280), .B2(new_n1287), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1260), .A2(new_n1277), .A3(new_n1279), .A4(new_n1288), .ZN(new_n1289));
  AOI22_X1  g1089(.A1(new_n1251), .A2(new_n1253), .B1(new_n1258), .B2(new_n1248), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT61), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1283), .A2(new_n1286), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1291), .B1(new_n1278), .B2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT62), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1275), .A2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1278), .A2(KEYINPUT62), .A3(new_n1274), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1293), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1290), .B1(new_n1297), .B2(KEYINPUT127), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1296), .ZN(new_n1299));
  AOI21_X1  g1099(.A(KEYINPUT62), .B1(new_n1278), .B2(new_n1274), .ZN(new_n1300));
  OAI211_X1 g1100(.A(KEYINPUT127), .B(new_n1288), .C1(new_n1299), .C2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1289), .B1(new_n1298), .B2(new_n1302), .ZN(G405));
  AOI21_X1  g1103(.A(G378), .B1(new_n1175), .B2(new_n1203), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1261), .ZN(new_n1305));
  OR3_X1    g1105(.A1(new_n1304), .A2(new_n1305), .A3(new_n1274), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1274), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  XNOR2_X1  g1108(.A(new_n1290), .B(new_n1308), .ZN(G402));
endmodule


