//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 1 1 0 1 0 0 0 1 0 0 0 1 0 1 1 1 0 0 0 1 0 0 0 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 1 0 0 0 0 0 0 0 1 0 1 1 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1272, new_n1273,
    new_n1274, new_n1275, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  INV_X1    g0009(.A(new_n202), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G50), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n206), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n209), .B(new_n216), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT65), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n232), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G58), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  INV_X1    g0040(.A(G107), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(G97), .ZN(new_n242));
  INV_X1    g0042(.A(G97), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G107), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n240), .B(new_n247), .ZN(G351));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(new_n213), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(KEYINPUT67), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT67), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n249), .A2(new_n252), .A3(new_n213), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n214), .A2(G68), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G20), .A2(G33), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n256), .B1(G50), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G77), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(G20), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n258), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(KEYINPUT11), .B1(new_n255), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n251), .A2(new_n253), .B1(new_n265), .B2(G20), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n264), .B1(G68), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n255), .A2(new_n263), .A3(KEYINPUT11), .ZN(new_n268));
  INV_X1    g0068(.A(G13), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(G1), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n256), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n271), .B1(KEYINPUT73), .B2(KEYINPUT12), .ZN(new_n272));
  NOR2_X1   g0072(.A1(KEYINPUT73), .A2(KEYINPUT12), .ZN(new_n273));
  XNOR2_X1  g0073(.A(new_n272), .B(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n267), .A2(new_n268), .A3(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT66), .B(G45), .ZN(new_n276));
  INV_X1    g0076(.A(G41), .ZN(new_n277));
  AND2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G274), .ZN(new_n279));
  AND2_X1   g0079(.A1(G1), .A2(G13), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n265), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n278), .A2(new_n283), .ZN(new_n284));
  AND2_X1   g0084(.A1(G33), .A2(G41), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(new_n213), .ZN(new_n286));
  INV_X1    g0086(.A(G45), .ZN(new_n287));
  AOI21_X1  g0087(.A(G1), .B1(new_n277), .B2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n284), .B1(G238), .B2(new_n289), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT3), .B(G33), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(G232), .A3(G1698), .ZN(new_n292));
  INV_X1    g0092(.A(G1698), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n291), .A2(G226), .A3(new_n293), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n292), .B(new_n294), .C1(new_n260), .C2(new_n243), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n286), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n290), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT13), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT13), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n290), .A2(new_n299), .A3(new_n296), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n298), .A2(G179), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n300), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n299), .B1(new_n290), .B2(new_n296), .ZN(new_n303));
  OAI21_X1  g0103(.A(G169), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n301), .B1(new_n304), .B2(KEYINPUT14), .ZN(new_n305));
  INV_X1    g0105(.A(G169), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n306), .B1(new_n298), .B2(new_n300), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT14), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n275), .B1(new_n305), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(G200), .B1(new_n302), .B2(new_n303), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n298), .A2(G190), .A3(new_n300), .ZN(new_n312));
  INV_X1    g0112(.A(new_n275), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT74), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT74), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n310), .A2(new_n317), .A3(new_n314), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n265), .A2(G13), .A3(G20), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G50), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n253), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n252), .B1(new_n249), .B2(new_n213), .ZN(new_n325));
  OAI22_X1  g0125(.A1(new_n324), .A2(new_n325), .B1(G1), .B2(new_n214), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n323), .B1(new_n326), .B2(new_n322), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT69), .ZN(new_n328));
  INV_X1    g0128(.A(G58), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT8), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT8), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G58), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n330), .A2(new_n332), .A3(KEYINPUT68), .ZN(new_n333));
  OR3_X1    g0133(.A1(new_n331), .A2(KEYINPUT68), .A3(G58), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n328), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n333), .A2(new_n334), .A3(new_n328), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n261), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n257), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n327), .B1(new_n341), .B2(new_n255), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT9), .ZN(new_n343));
  XNOR2_X1  g0143(.A(new_n342), .B(new_n343), .ZN(new_n344));
  AND2_X1   g0144(.A1(new_n289), .A2(G226), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n291), .A2(G222), .A3(new_n293), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n291), .A2(G1698), .ZN(new_n347));
  INV_X1    g0147(.A(G223), .ZN(new_n348));
  OAI221_X1 g0148(.A(new_n346), .B1(new_n259), .B2(new_n291), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  AOI211_X1 g0149(.A(new_n345), .B(new_n284), .C1(new_n349), .C2(new_n286), .ZN(new_n350));
  XOR2_X1   g0150(.A(KEYINPUT71), .B(G200), .Z(new_n351));
  NOR2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n352), .B1(G190), .B2(new_n350), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT72), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT10), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n344), .A2(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n354), .A2(new_n355), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n344), .A2(new_n353), .A3(KEYINPUT72), .A4(KEYINPUT10), .ZN(new_n360));
  INV_X1    g0160(.A(G179), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n350), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(G169), .B2(new_n350), .ZN(new_n363));
  OR2_X1    g0163(.A1(new_n363), .A2(new_n342), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n359), .A2(new_n360), .A3(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n291), .A2(G223), .A3(new_n293), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n291), .A2(G226), .A3(G1698), .ZN(new_n367));
  NAND2_X1  g0167(.A1(G33), .A2(G87), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n286), .ZN(new_n370));
  OAI21_X1  g0170(.A(G274), .B1(new_n285), .B2(new_n213), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n371), .A2(G1), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n276), .A2(new_n277), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n372), .A2(new_n373), .B1(new_n289), .B2(G232), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n370), .A2(G179), .A3(new_n374), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n370), .A2(new_n374), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n375), .B1(new_n376), .B2(new_n306), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT16), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT3), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n260), .ZN(new_n380));
  NAND2_X1  g0180(.A1(KEYINPUT3), .A2(G33), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(new_n214), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT7), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n380), .A2(KEYINPUT7), .A3(new_n214), .A4(new_n381), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n218), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n329), .A2(new_n218), .ZN(new_n387));
  OAI21_X1  g0187(.A(G20), .B1(new_n387), .B2(new_n202), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n257), .A2(G159), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n378), .B1(new_n386), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT75), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n384), .A2(new_n385), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n390), .B1(new_n393), .B2(G68), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n254), .B1(new_n394), .B2(KEYINPUT16), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT75), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n396), .B(new_n378), .C1(new_n386), .C2(new_n390), .ZN(new_n397));
  AND3_X1   g0197(.A1(new_n392), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n266), .B1(new_n336), .B2(new_n337), .ZN(new_n399));
  INV_X1    g0199(.A(new_n337), .ZN(new_n400));
  NOR3_X1   g0200(.A1(new_n400), .A2(new_n321), .A3(new_n335), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT76), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n326), .B1(new_n400), .B2(new_n335), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n336), .A2(new_n337), .A3(new_n320), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT76), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n377), .B1(new_n398), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT18), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT18), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n410), .B(new_n377), .C1(new_n398), .C2(new_n407), .ZN(new_n411));
  AND3_X1   g0211(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n405), .B1(new_n403), .B2(new_n404), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(G200), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n415), .B1(new_n370), .B2(new_n374), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n416), .B1(G190), .B2(new_n376), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n392), .A2(new_n395), .A3(new_n397), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n414), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT17), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n414), .A2(new_n417), .A3(KEYINPUT17), .A4(new_n418), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n409), .A2(new_n411), .A3(new_n421), .A4(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n284), .B1(G244), .B2(new_n289), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n291), .A2(G232), .A3(new_n293), .ZN(new_n425));
  OAI221_X1 g0225(.A(new_n425), .B1(new_n241), .B2(new_n291), .C1(new_n347), .C2(new_n219), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n286), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(G190), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n266), .A2(G77), .ZN(new_n431));
  XNOR2_X1  g0231(.A(KEYINPUT15), .B(G87), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT70), .ZN(new_n433));
  OR3_X1    g0233(.A1(new_n432), .A2(new_n262), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n330), .A2(new_n332), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n435), .A2(new_n257), .B1(G20), .B2(G77), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n433), .B1(new_n432), .B2(new_n262), .ZN(new_n437));
  AND3_X1   g0237(.A1(new_n434), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  OAI221_X1 g0238(.A(new_n431), .B1(G77), .B2(new_n320), .C1(new_n438), .C2(new_n254), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n351), .B1(new_n424), .B2(new_n427), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n430), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n428), .A2(new_n306), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n424), .A2(new_n427), .A3(new_n361), .ZN(new_n443));
  AND3_X1   g0243(.A1(new_n439), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  OR3_X1    g0244(.A1(new_n423), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  NOR3_X1   g0245(.A1(new_n319), .A2(new_n365), .A3(new_n445), .ZN(new_n446));
  XNOR2_X1  g0246(.A(KEYINPUT5), .B(G41), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n287), .A2(G1), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n447), .A2(new_n448), .B1(new_n280), .B2(new_n281), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(KEYINPUT80), .A3(G257), .ZN(new_n450));
  NAND2_X1  g0250(.A1(KEYINPUT5), .A2(G41), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(KEYINPUT5), .A2(G41), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n448), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n280), .A2(new_n281), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n454), .A2(G257), .A3(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT80), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT79), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n459), .B1(new_n454), .B2(new_n371), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n265), .A2(G45), .ZN(new_n461));
  OR2_X1    g0261(.A1(KEYINPUT5), .A2(G41), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n461), .B1(new_n462), .B2(new_n451), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n463), .A2(KEYINPUT79), .A3(new_n282), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n450), .A2(new_n458), .B1(new_n460), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT4), .ZN(new_n466));
  AND2_X1   g0266(.A1(KEYINPUT3), .A2(G33), .ZN(new_n467));
  NOR2_X1   g0267(.A1(KEYINPUT3), .A2(G33), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n293), .A2(G244), .ZN(new_n470));
  OAI211_X1 g0270(.A(KEYINPUT78), .B(new_n466), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n380), .A2(KEYINPUT78), .A3(new_n381), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(KEYINPUT78), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n472), .A2(KEYINPUT4), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G283), .ZN(new_n475));
  OAI211_X1 g0275(.A(G250), .B(G1698), .C1(new_n467), .C2(new_n468), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n471), .A2(new_n474), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n286), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n465), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n306), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n465), .A2(new_n361), .A3(new_n478), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n257), .A2(G77), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT77), .ZN(new_n483));
  XNOR2_X1  g0283(.A(new_n482), .B(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT6), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n242), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g0286(.A(G97), .B(G107), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n486), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n484), .B1(new_n488), .B2(new_n214), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n241), .B1(new_n384), .B2(new_n385), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n255), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n320), .A2(G97), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n320), .B1(G1), .B2(new_n260), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n493), .B1(new_n251), .B2(new_n253), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n492), .B1(new_n494), .B2(G97), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n480), .A2(new_n481), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n450), .A2(new_n458), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n460), .A2(new_n464), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(KEYINPUT4), .B1(new_n472), .B2(new_n473), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n476), .A2(new_n475), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n455), .B1(new_n503), .B2(new_n474), .ZN(new_n504));
  OAI21_X1  g0304(.A(G200), .B1(new_n500), .B2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n495), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n487), .A2(new_n485), .ZN(new_n507));
  INV_X1    g0307(.A(new_n486), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n214), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g0309(.A(new_n482), .B(KEYINPUT77), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n490), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n506), .B1(new_n513), .B2(new_n255), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n465), .A2(G190), .A3(new_n478), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n505), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n262), .A2(new_n243), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n214), .A2(G68), .ZN(new_n518));
  OAI22_X1  g0318(.A1(new_n517), .A2(KEYINPUT19), .B1(new_n469), .B2(new_n518), .ZN(new_n519));
  XNOR2_X1  g0319(.A(KEYINPUT83), .B(G87), .ZN(new_n520));
  NOR2_X1   g0320(.A1(G97), .A2(G107), .ZN(new_n521));
  NAND3_X1  g0321(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n520), .A2(new_n521), .B1(new_n214), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n255), .B1(new_n519), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n432), .A2(new_n321), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n494), .A2(G87), .ZN(new_n526));
  AND3_X1   g0326(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  OAI211_X1 g0327(.A(G244), .B(G1698), .C1(new_n467), .C2(new_n468), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT82), .ZN(new_n529));
  XNOR2_X1  g0329(.A(new_n528), .B(new_n529), .ZN(new_n530));
  OAI211_X1 g0330(.A(G238), .B(new_n293), .C1(new_n467), .C2(new_n468), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(KEYINPUT81), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT81), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n291), .A2(new_n533), .A3(G238), .A4(new_n293), .ZN(new_n534));
  NAND2_X1  g0334(.A1(G33), .A2(G116), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n532), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n286), .B1(new_n530), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n448), .A2(new_n221), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n455), .A2(new_n538), .B1(new_n282), .B2(new_n448), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(G190), .A3(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n539), .ZN(new_n541));
  XNOR2_X1  g0341(.A(new_n528), .B(KEYINPUT82), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n531), .A2(KEYINPUT81), .B1(G33), .B2(G116), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n542), .A2(new_n534), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n541), .B1(new_n544), .B2(new_n286), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n527), .B(new_n540), .C1(new_n545), .C2(new_n351), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n537), .A2(new_n361), .A3(new_n539), .ZN(new_n547));
  XOR2_X1   g0347(.A(new_n432), .B(KEYINPUT84), .Z(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n494), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n524), .A2(new_n549), .A3(new_n525), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n547), .B(new_n550), .C1(new_n545), .C2(G169), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n497), .A2(new_n516), .A3(new_n546), .A4(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(G257), .B(G1698), .C1(new_n467), .C2(new_n468), .ZN(new_n553));
  OAI211_X1 g0353(.A(G250), .B(new_n293), .C1(new_n467), .C2(new_n468), .ZN(new_n554));
  INV_X1    g0354(.A(G294), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n553), .B(new_n554), .C1(new_n260), .C2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n286), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT90), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n558), .B1(new_n449), .B2(G264), .ZN(new_n559));
  AND4_X1   g0359(.A1(new_n558), .A2(new_n454), .A3(G264), .A4(new_n455), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n557), .B(new_n499), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n415), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n449), .A2(G264), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n557), .A2(new_n499), .A3(new_n429), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT25), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n320), .B2(G107), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n321), .A2(KEYINPUT25), .A3(new_n241), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n494), .A2(G107), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n535), .A2(G20), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT23), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(new_n214), .B2(G107), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n241), .A2(KEYINPUT23), .A3(G20), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n570), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(KEYINPUT87), .A2(G20), .ZN(new_n575));
  OAI211_X1 g0375(.A(G87), .B(new_n575), .C1(new_n467), .C2(new_n468), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT22), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT88), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT88), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(KEYINPUT22), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  NOR3_X1   g0382(.A1(new_n220), .A2(KEYINPUT87), .A3(G20), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n291), .A2(new_n583), .B1(new_n578), .B2(new_n580), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n574), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT24), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n575), .A2(G87), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n581), .B1(new_n469), .B2(new_n587), .ZN(new_n588));
  XNOR2_X1  g0388(.A(KEYINPUT88), .B(KEYINPUT22), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n291), .A2(new_n589), .A3(new_n583), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT24), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(new_n592), .A3(new_n574), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n586), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT89), .B1(new_n594), .B2(new_n255), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT89), .ZN(new_n596));
  AOI211_X1 g0396(.A(new_n596), .B(new_n254), .C1(new_n586), .C2(new_n593), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n565), .B(new_n569), .C1(new_n595), .C2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT91), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n591), .A2(new_n592), .A3(new_n574), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n592), .B1(new_n591), .B2(new_n574), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n255), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n596), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n594), .A2(KEYINPUT89), .A3(new_n255), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n606), .A2(KEYINPUT91), .A3(new_n565), .A4(new_n569), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n552), .B1(new_n600), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT86), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n609), .A2(KEYINPUT21), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n449), .A2(G270), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n499), .A2(new_n611), .ZN(new_n612));
  OAI211_X1 g0412(.A(G264), .B(G1698), .C1(new_n467), .C2(new_n468), .ZN(new_n613));
  OAI211_X1 g0413(.A(G257), .B(new_n293), .C1(new_n467), .C2(new_n468), .ZN(new_n614));
  INV_X1    g0414(.A(G303), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n613), .B(new_n614), .C1(new_n615), .C2(new_n291), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n616), .A2(new_n286), .ZN(new_n617));
  OAI21_X1  g0417(.A(G169), .B1(new_n612), .B2(new_n617), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n270), .A2(G20), .B1(new_n265), .B2(G33), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n619), .B(G116), .C1(new_n324), .C2(new_n325), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n320), .A2(G116), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(G116), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n249), .A2(new_n213), .B1(G20), .B2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(G20), .B1(G33), .B2(G283), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n260), .A2(G97), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT85), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n628), .B1(new_n626), .B2(new_n627), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n625), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT20), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI211_X1 g0433(.A(KEYINPUT20), .B(new_n625), .C1(new_n629), .C2(new_n630), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n623), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n610), .B1(new_n618), .B2(new_n635), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n460), .A2(new_n464), .B1(new_n449), .B2(G270), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n616), .A2(new_n286), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(G190), .A3(new_n638), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n638), .A2(new_n499), .A3(new_n611), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n635), .B(new_n639), .C1(new_n640), .C2(new_n415), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n621), .B1(new_n494), .B2(G116), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n626), .A2(new_n627), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(KEYINPUT85), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(KEYINPUT20), .B1(new_n646), .B2(new_n625), .ZN(new_n647));
  INV_X1    g0447(.A(new_n634), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n642), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n640), .A2(new_n649), .A3(G179), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n637), .A2(new_n638), .ZN(new_n651));
  INV_X1    g0451(.A(new_n610), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n649), .A2(new_n651), .A3(G169), .A4(new_n652), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n636), .A2(new_n641), .A3(new_n650), .A4(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n606), .A2(new_n569), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n563), .A2(KEYINPUT90), .ZN(new_n656));
  INV_X1    g0456(.A(new_n560), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n656), .A2(new_n657), .B1(new_n286), .B2(new_n556), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n658), .A2(G179), .A3(new_n499), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n557), .A2(new_n499), .A3(new_n563), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(G169), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n654), .B1(new_n655), .B2(new_n662), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n446), .A2(new_n608), .A3(new_n663), .ZN(G372));
  INV_X1    g0464(.A(new_n364), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n314), .A2(new_n444), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n310), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n667), .A2(new_n421), .A3(new_n422), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n668), .A2(new_n409), .A3(new_n411), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n359), .A2(new_n360), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n665), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n446), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n480), .A2(new_n481), .A3(new_n496), .ZN(new_n673));
  XOR2_X1   g0473(.A(KEYINPUT93), .B(KEYINPUT26), .Z(new_n674));
  NAND4_X1  g0474(.A1(new_n673), .A2(new_n551), .A3(new_n546), .A4(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n551), .B1(new_n675), .B2(KEYINPUT94), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n546), .A2(new_n551), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n673), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT26), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n675), .A2(KEYINPUT94), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n676), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n653), .A2(new_n650), .ZN(new_n683));
  INV_X1    g0483(.A(new_n569), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n684), .B1(new_n604), .B2(new_n605), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n659), .A2(new_n661), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n636), .B(new_n683), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  AND4_X1   g0487(.A1(new_n497), .A2(new_n516), .A3(new_n546), .A4(new_n551), .ZN(new_n688));
  INV_X1    g0488(.A(new_n607), .ZN(new_n689));
  AOI21_X1  g0489(.A(KEYINPUT91), .B1(new_n685), .B2(new_n565), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n687), .B(new_n688), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT92), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(KEYINPUT92), .B1(new_n608), .B2(new_n687), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n682), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n671), .B1(new_n672), .B2(new_n696), .ZN(G369));
  NOR2_X1   g0497(.A1(new_n685), .A2(new_n686), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n270), .A2(new_n214), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(KEYINPUT27), .ZN(new_n700));
  XOR2_X1   g0500(.A(new_n700), .B(KEYINPUT95), .Z(new_n701));
  INV_X1    g0501(.A(G213), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n702), .B1(new_n699), .B2(KEYINPUT27), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(G343), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n698), .A2(new_n706), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n707), .A2(KEYINPUT97), .ZN(new_n708));
  INV_X1    g0508(.A(new_n706), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n685), .B1(new_n686), .B2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n710), .B1(new_n600), .B2(new_n607), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n707), .A2(KEYINPUT97), .ZN(new_n712));
  OR3_X1    g0512(.A1(new_n708), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n709), .A2(new_n635), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT96), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n715), .B1(new_n654), .B2(new_n716), .ZN(new_n717));
  OR2_X1    g0517(.A1(new_n654), .A2(new_n716), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n683), .A2(new_n636), .ZN(new_n719));
  AOI22_X1  g0519(.A1(new_n717), .A2(new_n718), .B1(new_n719), .B2(new_n715), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G330), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n714), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n698), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n706), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n719), .A2(new_n706), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n725), .B1(new_n713), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n723), .A2(new_n727), .ZN(G399));
  INV_X1    g0528(.A(new_n207), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G41), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n520), .A2(new_n624), .A3(new_n521), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n730), .A2(new_n731), .A3(new_n265), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT98), .ZN(new_n733));
  AOI22_X1  g0533(.A1(new_n732), .A2(new_n733), .B1(new_n212), .B2(new_n730), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(new_n733), .B2(new_n732), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT28), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT29), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n678), .A2(new_n674), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n677), .A2(new_n679), .A3(new_n673), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n691), .A2(new_n551), .A3(new_n738), .A4(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n737), .B1(new_n740), .B2(new_n709), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n691), .A2(new_n692), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n608), .A2(KEYINPUT92), .A3(new_n687), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n706), .B1(new_n744), .B2(new_n682), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n741), .B1(new_n745), .B2(new_n737), .ZN(new_n746));
  INV_X1    g0546(.A(G330), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n600), .A2(new_n607), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n748), .A2(new_n688), .A3(new_n663), .A4(new_n709), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT101), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n608), .A2(KEYINPUT101), .A3(new_n663), .A4(new_n709), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n479), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n651), .A2(new_n361), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n754), .A2(new_n545), .A3(new_n755), .A4(new_n658), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT30), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AND3_X1   g0558(.A1(new_n658), .A2(new_n478), .A3(new_n465), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n759), .A2(KEYINPUT30), .A3(new_n545), .A4(new_n755), .ZN(new_n760));
  AOI21_X1  g0560(.A(G179), .B1(new_n637), .B2(new_n638), .ZN(new_n761));
  AND3_X1   g0561(.A1(new_n479), .A2(new_n561), .A3(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n545), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n758), .A2(new_n760), .A3(new_n764), .ZN(new_n765));
  XNOR2_X1  g0565(.A(KEYINPUT99), .B(KEYINPUT31), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AND4_X1   g0567(.A1(KEYINPUT100), .A2(new_n765), .A3(new_n706), .A4(new_n767), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n756), .A2(new_n757), .B1(new_n762), .B2(new_n763), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n709), .B1(new_n769), .B2(new_n760), .ZN(new_n770));
  OAI21_X1  g0570(.A(KEYINPUT100), .B1(new_n770), .B2(KEYINPUT31), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n767), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n768), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n747), .B1(new_n753), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n746), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n736), .B1(new_n777), .B2(G1), .ZN(G364));
  NOR2_X1   g0578(.A1(new_n720), .A2(G330), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT102), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n269), .A2(G20), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n265), .B1(new_n781), .B2(G45), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n730), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n780), .A2(new_n721), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n213), .B1(G20), .B2(new_n306), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n214), .A2(new_n361), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n789), .A2(G190), .A3(new_n415), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n214), .A2(G179), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G190), .A2(G200), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n791), .A2(G322), .B1(new_n795), .B2(G329), .ZN(new_n796));
  INV_X1    g0596(.A(G311), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n789), .A2(new_n793), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n796), .B(new_n469), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n351), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n800), .A2(new_n429), .A3(new_n792), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n799), .B1(G283), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n789), .A2(G200), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(G190), .ZN(new_n805));
  NOR2_X1   g0605(.A1(KEYINPUT33), .A2(G317), .ZN(new_n806));
  AND2_X1   g0606(.A1(KEYINPUT33), .A2(G317), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n804), .A2(new_n429), .ZN(new_n809));
  XOR2_X1   g0609(.A(KEYINPUT105), .B(G326), .Z(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n361), .A2(new_n415), .A3(G190), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G20), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n809), .A2(new_n811), .B1(G294), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n803), .A2(new_n808), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n800), .A2(G190), .A3(new_n792), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  OR2_X1    g0617(.A1(new_n817), .A2(KEYINPUT104), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(KEYINPUT104), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n820), .A2(new_n615), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n820), .A2(new_n520), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n291), .B1(new_n798), .B2(new_n259), .C1(new_n329), .C2(new_n790), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT32), .ZN(new_n824));
  INV_X1    g0624(.A(G159), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n824), .B1(new_n794), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n795), .A2(KEYINPUT32), .A3(G159), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n823), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n809), .A2(G50), .ZN(new_n829));
  INV_X1    g0629(.A(new_n813), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n830), .A2(new_n243), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(G68), .B2(new_n805), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n802), .A2(G107), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n828), .A2(new_n829), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n815), .A2(new_n821), .B1(new_n822), .B2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT106), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n788), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n836), .B2(new_n835), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n729), .A2(new_n469), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n839), .A2(G355), .B1(new_n624), .B2(new_n729), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n240), .A2(new_n287), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n729), .A2(new_n291), .ZN(new_n842));
  INV_X1    g0642(.A(new_n276), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n842), .B1(new_n211), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n840), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n269), .A2(new_n260), .A3(KEYINPUT103), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT103), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(G13), .B2(G33), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n850), .A2(G20), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n851), .A2(new_n787), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n785), .B1(new_n845), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n851), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n838), .B(new_n853), .C1(new_n720), .C2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n786), .A2(new_n855), .ZN(G396));
  NAND2_X1  g0656(.A1(new_n695), .A2(new_n709), .ZN(new_n857));
  AND2_X1   g0657(.A1(new_n706), .A2(new_n439), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n441), .A2(new_n858), .ZN(new_n859));
  OR2_X1    g0659(.A1(new_n859), .A2(new_n444), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n444), .A2(new_n709), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n862), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n695), .A2(new_n709), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n785), .B1(new_n866), .B2(new_n775), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n867), .A2(KEYINPUT109), .B1(new_n775), .B2(new_n866), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(KEYINPUT109), .B2(new_n867), .ZN(new_n869));
  XOR2_X1   g0669(.A(KEYINPUT108), .B(G143), .Z(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n798), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n791), .A2(new_n871), .B1(new_n872), .B2(G159), .ZN(new_n873));
  INV_X1    g0673(.A(new_n805), .ZN(new_n874));
  INV_X1    g0674(.A(G150), .ZN(new_n875));
  INV_X1    g0675(.A(G137), .ZN(new_n876));
  INV_X1    g0676(.A(new_n809), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n873), .B1(new_n874), .B2(new_n875), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  XOR2_X1   g0678(.A(new_n878), .B(KEYINPUT34), .Z(new_n879));
  NAND2_X1  g0679(.A1(new_n802), .A2(G68), .ZN(new_n880));
  INV_X1    g0680(.A(G132), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n291), .B1(new_n794), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(G58), .B2(new_n813), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n880), .B(new_n883), .C1(new_n820), .C2(new_n322), .ZN(new_n884));
  XNOR2_X1  g0684(.A(KEYINPUT107), .B(G283), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n874), .A2(new_n885), .ZN(new_n886));
  AOI211_X1 g0686(.A(new_n831), .B(new_n886), .C1(G303), .C2(new_n809), .ZN(new_n887));
  OAI22_X1  g0687(.A1(new_n798), .A2(new_n624), .B1(new_n794), .B2(new_n797), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n291), .B(new_n888), .C1(G294), .C2(new_n791), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n887), .B(new_n889), .C1(new_n220), .C2(new_n801), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n820), .A2(new_n241), .ZN(new_n891));
  OAI22_X1  g0691(.A1(new_n879), .A2(new_n884), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n787), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n849), .A2(new_n787), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n785), .B1(new_n259), .B2(new_n894), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n893), .B(new_n895), .C1(new_n864), .C2(new_n850), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n869), .A2(new_n896), .ZN(G384));
  OR3_X1    g0697(.A1(new_n211), .A2(new_n259), .A3(new_n387), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n201), .A2(G68), .ZN(new_n899));
  AOI211_X1 g0699(.A(new_n265), .B(G13), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT111), .ZN(new_n901));
  INV_X1    g0701(.A(new_n488), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n902), .A2(KEYINPUT35), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(KEYINPUT35), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n903), .A2(G116), .A3(new_n215), .A4(new_n904), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n905), .B(KEYINPUT36), .Z(new_n906));
  INV_X1    g0706(.A(KEYINPUT110), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n901), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(new_n907), .B2(new_n906), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n395), .A2(new_n391), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n399), .A2(new_n401), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n912), .A2(new_n704), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n423), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n704), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n398), .B2(new_n407), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT37), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n408), .A2(new_n916), .A3(new_n917), .A4(new_n419), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n910), .A2(new_n911), .B1(new_n377), .B2(new_n915), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n919), .A2(new_n419), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n918), .B1(new_n920), .B2(new_n917), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n914), .A2(KEYINPUT38), .A3(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT39), .ZN(new_n923));
  INV_X1    g0723(.A(new_n916), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n408), .A2(new_n916), .A3(new_n419), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(KEYINPUT37), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n423), .A2(new_n924), .B1(new_n926), .B2(new_n918), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n922), .B(new_n923), .C1(new_n927), .C2(KEYINPUT38), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n914), .A2(new_n921), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT38), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n923), .B1(new_n932), .B2(new_n922), .ZN(new_n933));
  OAI21_X1  g0733(.A(KEYINPUT112), .B1(new_n929), .B2(new_n933), .ZN(new_n934));
  AND3_X1   g0734(.A1(new_n914), .A2(KEYINPUT38), .A3(new_n921), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT38), .B1(new_n914), .B2(new_n921), .ZN(new_n936));
  OAI21_X1  g0736(.A(KEYINPUT39), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT112), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n937), .A2(new_n938), .A3(new_n928), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n304), .A2(KEYINPUT14), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n307), .A2(new_n308), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n940), .A2(new_n941), .A3(new_n301), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n942), .A2(new_n275), .A3(new_n709), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n934), .A2(new_n939), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n865), .A2(new_n861), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n932), .A2(new_n922), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n275), .A2(new_n706), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n310), .A2(new_n314), .A3(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n314), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n275), .B(new_n706), .C1(new_n942), .C2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n946), .A2(new_n947), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n409), .A2(new_n411), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n704), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n945), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n671), .ZN(new_n957));
  INV_X1    g0757(.A(new_n741), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n857), .B2(KEYINPUT29), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n957), .B1(new_n959), .B2(new_n446), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n956), .B(new_n960), .Z(new_n961));
  NAND3_X1  g0761(.A1(new_n765), .A2(KEYINPUT31), .A3(new_n706), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n770), .B2(new_n767), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n753), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n862), .B1(new_n949), .B2(new_n951), .ZN(new_n966));
  OR2_X1    g0766(.A1(KEYINPUT113), .A2(KEYINPUT40), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT113), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n963), .B1(new_n751), .B2(new_n752), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n864), .A2(new_n952), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n968), .A2(new_n947), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n922), .B1(new_n927), .B2(KEYINPUT38), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n965), .A2(new_n974), .A3(new_n966), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(KEYINPUT40), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n672), .A2(new_n970), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n747), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n978), .B2(new_n977), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n961), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n265), .B2(new_n781), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n961), .A2(new_n980), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n909), .B1(new_n982), .B2(new_n983), .ZN(G367));
  OAI211_X1 g0784(.A(new_n497), .B(new_n516), .C1(new_n709), .C2(new_n514), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n497), .B2(new_n709), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n713), .A2(new_n726), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n497), .B1(new_n724), .B2(new_n985), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n987), .A2(KEYINPUT42), .B1(new_n709), .B2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT42), .ZN(new_n990));
  INV_X1    g0790(.A(new_n987), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n989), .A2(KEYINPUT114), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n988), .A2(new_n709), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n991), .B2(new_n990), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT114), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n709), .A2(new_n527), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n997), .A2(new_n551), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n677), .A2(new_n997), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n992), .A2(new_n996), .B1(KEYINPUT43), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1000), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT43), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n722), .A2(new_n986), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n992), .A2(new_n996), .A3(new_n1003), .A4(new_n1002), .ZN(new_n1008));
  AND3_X1   g0808(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1007), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n730), .B(KEYINPUT41), .Z(new_n1012));
  INV_X1    g0812(.A(KEYINPUT45), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT115), .ZN(new_n1014));
  AND3_X1   g0814(.A1(new_n727), .A2(new_n1014), .A3(new_n986), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1014), .B1(new_n727), .B2(new_n986), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1013), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n727), .A2(new_n986), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(KEYINPUT115), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n727), .A2(new_n1014), .A3(new_n986), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1019), .A2(KEYINPUT45), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT44), .ZN(new_n1022));
  OR3_X1    g0822(.A1(new_n727), .A2(new_n1022), .A3(new_n986), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1022), .B1(new_n727), .B2(new_n986), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1017), .A2(new_n1021), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n722), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n726), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n713), .B(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(new_n721), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1017), .A2(new_n1021), .A3(new_n1025), .A4(new_n723), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1027), .A2(new_n777), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1012), .B1(new_n1032), .B2(new_n777), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1011), .B1(new_n1033), .B2(new_n783), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n842), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n236), .A2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n852), .B1(new_n207), .B2(new_n432), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n784), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT46), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n820), .B2(new_n624), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n874), .A2(new_n555), .B1(new_n877), .B2(new_n797), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(G107), .B2(new_n813), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n802), .A2(G97), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n469), .B1(new_n790), .B2(new_n615), .ZN(new_n1044));
  INV_X1    g0844(.A(G317), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n798), .A2(new_n885), .B1(new_n794), .B2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1040), .A2(new_n1042), .A3(new_n1043), .A4(new_n1047), .ZN(new_n1048));
  NOR3_X1   g0848(.A1(new_n820), .A2(new_n1039), .A3(new_n624), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n820), .A2(new_n329), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n790), .A2(new_n875), .B1(new_n794), .B2(new_n876), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n201), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n469), .B(new_n1051), .C1(new_n1052), .C2(new_n872), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n809), .A2(new_n871), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n830), .A2(new_n218), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(G159), .B2(new_n805), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n802), .A2(G77), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1053), .A2(new_n1054), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n1048), .A2(new_n1049), .B1(new_n1050), .B2(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT47), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1038), .B1(new_n1060), .B2(new_n787), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n854), .B2(new_n1000), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1034), .A2(new_n1062), .ZN(G387));
  OR2_X1    g0863(.A1(new_n1030), .A2(new_n777), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1030), .A2(new_n777), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1064), .A2(new_n730), .A3(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n469), .B1(new_n810), .B2(new_n794), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n791), .A2(G317), .B1(new_n872), .B2(G303), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n809), .A2(G322), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1068), .B(new_n1069), .C1(new_n797), .C2(new_n874), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT48), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1071), .B1(new_n555), .B2(new_n820), .C1(new_n830), .C2(new_n885), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT49), .Z(new_n1073));
  AOI211_X1 g0873(.A(new_n1067), .B(new_n1073), .C1(G116), .C2(new_n802), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n790), .A2(new_n322), .B1(new_n794), .B2(new_n875), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n469), .B(new_n1075), .C1(G68), .C2(new_n872), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n809), .A2(G159), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n548), .A2(new_n813), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1076), .A2(new_n1043), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n820), .A2(new_n259), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n1079), .B(new_n1080), .C1(new_n338), .C2(new_n805), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n787), .B1(new_n1074), .B2(new_n1081), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n232), .A2(new_n276), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n1083), .A2(new_n842), .B1(new_n731), .B2(new_n839), .ZN(new_n1084));
  AOI211_X1 g0884(.A(G45), .B(new_n731), .C1(G68), .C2(G77), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT50), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n435), .A2(new_n322), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT116), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1085), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n1084), .A2(new_n1090), .B1(G107), .B2(new_n207), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n785), .B1(new_n1091), .B2(new_n852), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1082), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n714), .B2(new_n851), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(new_n1030), .B2(new_n783), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1066), .A2(new_n1095), .ZN(G393));
  NAND2_X1  g0896(.A1(new_n1027), .A2(new_n1031), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n1065), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1098), .A2(new_n730), .A3(new_n1032), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1027), .A2(new_n783), .A3(new_n1031), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n852), .B1(new_n243), .B2(new_n207), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n247), .A2(new_n1035), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n784), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  OR2_X1    g0903(.A1(new_n820), .A2(new_n885), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n877), .A2(new_n1045), .B1(new_n797), .B2(new_n790), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT52), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n469), .B1(new_n798), .B2(new_n555), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n874), .A2(new_n615), .B1(new_n624), .B2(new_n830), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1107), .B(new_n1108), .C1(G322), .C2(new_n795), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1104), .A2(new_n833), .A3(new_n1106), .A4(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n820), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n1111), .A2(G68), .B1(new_n795), .B2(new_n871), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1113), .A2(KEYINPUT117), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(G150), .A2(new_n809), .B1(new_n791), .B2(G159), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT51), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n801), .A2(new_n220), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n830), .A2(new_n259), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n469), .B1(new_n872), .B2(new_n435), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n874), .B2(new_n201), .ZN(new_n1120));
  NOR4_X1   g0920(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .A4(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT117), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1121), .B1(new_n1112), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1110), .B1(new_n1114), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1103), .B1(new_n1124), .B2(new_n787), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n986), .B2(new_n854), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1100), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1099), .A2(new_n1127), .ZN(G390));
  NOR2_X1   g0928(.A1(new_n970), .A2(new_n747), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n446), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1130), .B(new_n671), .C1(new_n746), .C2(new_n672), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n952), .B1(new_n774), .B2(new_n864), .ZN(new_n1132));
  NOR3_X1   g0932(.A1(new_n970), .A2(new_n971), .A3(new_n747), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n946), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n774), .A2(new_n864), .A3(new_n952), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n740), .A2(new_n709), .A3(new_n860), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n861), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  NOR3_X1   g0938(.A1(new_n970), .A2(new_n747), .A3(new_n862), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1135), .B(new_n1138), .C1(new_n952), .C2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1131), .B1(new_n1134), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n974), .A2(new_n943), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(new_n1137), .B2(new_n952), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n937), .A2(new_n938), .A3(new_n928), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n938), .B1(new_n937), .B2(new_n928), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n944), .B1(new_n946), .B2(new_n952), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1144), .B(new_n1135), .C1(new_n1147), .C2(new_n1148), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n745), .A2(new_n860), .B1(new_n444), .B2(new_n709), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n952), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n943), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n934), .A2(new_n939), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1143), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1133), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1141), .B(new_n1149), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1149), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1141), .ZN(new_n1158));
  AND3_X1   g0958(.A1(new_n1157), .A2(KEYINPUT118), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT118), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n730), .B(new_n1156), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1161));
  OR2_X1    g0961(.A1(new_n1157), .A2(new_n782), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n894), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n784), .B1(new_n338), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1111), .A2(G87), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n874), .A2(new_n241), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1118), .B(new_n1166), .C1(G283), .C2(new_n809), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n798), .A2(new_n243), .B1(new_n794), .B2(new_n555), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n291), .B(new_n1168), .C1(G116), .C2(new_n791), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1165), .A2(new_n880), .A3(new_n1167), .A4(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1111), .A2(G150), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT53), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n291), .B1(new_n801), .B2(new_n201), .ZN(new_n1173));
  OR2_X1    g0973(.A1(new_n1173), .A2(KEYINPUT119), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n874), .A2(new_n876), .B1(new_n825), .B2(new_n830), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(G128), .B2(new_n809), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1173), .A2(KEYINPUT119), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(KEYINPUT54), .B(G143), .ZN(new_n1178));
  INV_X1    g0978(.A(G125), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n798), .A2(new_n1178), .B1(new_n794), .B2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(G132), .B2(new_n791), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1174), .A2(new_n1176), .A3(new_n1177), .A4(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1170), .B1(new_n1172), .B2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1164), .B1(new_n1183), .B2(new_n787), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n1147), .B2(new_n850), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1161), .A2(new_n1162), .A3(new_n1185), .ZN(G378));
  INV_X1    g0986(.A(G128), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n790), .A2(new_n1187), .B1(new_n798), .B2(new_n876), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(G132), .B2(new_n805), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n809), .A2(G125), .B1(G150), .B2(new_n813), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1189), .B(new_n1190), .C1(new_n820), .C2(new_n1178), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n1191), .A2(KEYINPUT59), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(KEYINPUT59), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n802), .A2(G159), .ZN(new_n1194));
  AOI211_X1 g0994(.A(G33), .B(G41), .C1(new_n795), .C2(G124), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n548), .A2(new_n872), .B1(G97), .B2(new_n805), .ZN(new_n1197));
  XOR2_X1   g0997(.A(new_n1197), .B(KEYINPUT120), .Z(new_n1198));
  NAND2_X1  g0998(.A1(new_n802), .A2(G58), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1055), .B1(G116), .B2(new_n809), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n791), .A2(G107), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n469), .A2(new_n277), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G283), .B2(new_n795), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .A4(new_n1203), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(new_n1198), .A2(new_n1080), .A3(new_n1204), .ZN(new_n1205));
  OR2_X1    g1005(.A1(new_n1205), .A2(KEYINPUT58), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(KEYINPUT58), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1202), .B(new_n322), .C1(G33), .C2(G41), .ZN(new_n1208));
  AND4_X1   g1008(.A1(new_n1196), .A2(new_n1206), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n784), .B1(new_n1052), .B2(new_n1163), .C1(new_n1209), .C2(new_n788), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n342), .A2(new_n704), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n365), .B(new_n1211), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1212), .B(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1210), .B1(new_n1214), .B2(new_n849), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n977), .A2(G330), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1216), .A2(new_n953), .A3(new_n945), .A4(new_n955), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n747), .B1(new_n973), .B2(new_n976), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n956), .A2(new_n1218), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1217), .A2(new_n1214), .A3(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1214), .B1(new_n1217), .B2(new_n1219), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1215), .B1(new_n1222), .B2(new_n783), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1131), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1156), .A2(new_n1224), .ZN(new_n1225));
  OAI211_X1 g1025(.A(KEYINPUT57), .B(new_n1225), .C1(new_n1220), .C2(new_n1221), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1226), .A2(KEYINPUT121), .A3(new_n730), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1225), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT57), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1227), .A2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT121), .B1(new_n1226), .B2(new_n730), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1223), .B1(new_n1231), .B2(new_n1232), .ZN(G375));
  OAI21_X1  g1033(.A(new_n784), .B1(G68), .B2(new_n1163), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n881), .A2(new_n877), .B1(new_n874), .B2(new_n1178), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G50), .B2(new_n813), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n291), .B1(new_n794), .B2(new_n1187), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n790), .A2(new_n876), .B1(new_n798), .B2(new_n875), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n1237), .B(new_n1238), .C1(new_n802), .C2(G58), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1236), .B(new_n1239), .C1(new_n820), .C2(new_n825), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n820), .A2(new_n243), .B1(new_n615), .B2(new_n794), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1241), .B(KEYINPUT124), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1057), .A2(new_n469), .ZN(new_n1243));
  XOR2_X1   g1043(.A(new_n1243), .B(KEYINPUT123), .Z(new_n1244));
  INV_X1    g1044(.A(G283), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n790), .A2(new_n1245), .B1(new_n798), .B2(new_n241), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n877), .A2(new_n555), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n1246), .B(new_n1247), .C1(G116), .C2(new_n805), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1244), .A2(new_n1248), .A3(new_n1078), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1240), .B1(new_n1242), .B2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1234), .B1(new_n1250), .B2(new_n787), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n952), .B2(new_n850), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1134), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1140), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1252), .B1(new_n1255), .B2(new_n782), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT125), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1256), .B(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1255), .A2(new_n1131), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1012), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1260), .A2(new_n1261), .A3(new_n1158), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1259), .B1(KEYINPUT122), .B2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(KEYINPUT122), .B2(new_n1263), .ZN(G381));
  INV_X1    g1065(.A(G390), .ZN(new_n1266));
  INV_X1    g1066(.A(G384), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(G393), .A2(G396), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1266), .A2(new_n1267), .A3(new_n1268), .ZN(new_n1269));
  OR2_X1    g1069(.A1(new_n1269), .A2(G387), .ZN(new_n1270));
  OR4_X1    g1070(.A1(G378), .A2(new_n1270), .A3(G375), .A4(G381), .ZN(G407));
  INV_X1    g1071(.A(G378), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n705), .A2(G213), .ZN(new_n1273));
  XOR2_X1   g1073(.A(new_n1273), .B(KEYINPUT126), .Z(new_n1274));
  NAND2_X1  g1074(.A1(new_n1272), .A2(new_n1274), .ZN(new_n1275));
  OAI211_X1 g1075(.A(G407), .B(G213), .C1(G375), .C2(new_n1275), .ZN(G409));
  OAI211_X1 g1076(.A(G378), .B(new_n1223), .C1(new_n1231), .C2(new_n1232), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1223), .B1(new_n1012), .B2(new_n1228), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n1272), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1277), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1274), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(KEYINPUT127), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT60), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1260), .B1(new_n1284), .B2(new_n1141), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1255), .A2(KEYINPUT60), .A3(new_n1131), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1285), .A2(new_n730), .A3(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1258), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n1267), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1258), .A2(new_n1287), .A3(G384), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(new_n1289), .A2(new_n1290), .B1(G2897), .B2(new_n1274), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1258), .A2(G384), .A3(new_n1287), .ZN(new_n1292));
  AOI21_X1  g1092(.A(G384), .B1(new_n1258), .B2(new_n1287), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1274), .A2(G2897), .ZN(new_n1294));
  NOR3_X1   g1094(.A1(new_n1292), .A2(new_n1293), .A3(new_n1294), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1291), .A2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1274), .B1(new_n1277), .B2(new_n1279), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT127), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1296), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1283), .A2(new_n1299), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1297), .A2(KEYINPUT63), .A3(new_n1301), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1034), .A2(new_n1062), .A3(G390), .ZN(new_n1303));
  AOI21_X1  g1103(.A(G390), .B1(new_n1034), .B2(new_n1062), .ZN(new_n1304));
  AND2_X1   g1104(.A1(G393), .A2(G396), .ZN(new_n1305));
  OAI22_X1  g1105(.A1(new_n1303), .A2(new_n1304), .B1(new_n1268), .B2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(G387), .A2(new_n1266), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1305), .A2(new_n1268), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1034), .A2(new_n1062), .A3(G390), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1307), .A2(new_n1308), .A3(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT61), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1306), .A2(new_n1310), .A3(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1280), .A2(new_n1281), .A3(new_n1301), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT63), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1312), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1300), .A2(new_n1302), .A3(new_n1315), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1313), .A2(KEYINPUT62), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1311), .B1(new_n1297), .B2(new_n1296), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT62), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1319), .B1(new_n1297), .B2(new_n1301), .ZN(new_n1320));
  NOR3_X1   g1120(.A1(new_n1317), .A2(new_n1318), .A3(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1306), .A2(new_n1310), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1316), .B1(new_n1321), .B2(new_n1323), .ZN(G405));
  NAND2_X1  g1124(.A1(G375), .A2(new_n1272), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(new_n1277), .ZN(new_n1326));
  AND2_X1   g1126(.A1(new_n1326), .A2(new_n1301), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1326), .A2(new_n1301), .ZN(new_n1328));
  OR3_X1    g1128(.A1(new_n1327), .A2(new_n1328), .A3(new_n1322), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1322), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(G402));
endmodule


