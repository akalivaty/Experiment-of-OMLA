

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U553 ( .A(KEYINPUT1), .B(n538), .Z(n668) );
  OR2_X1 U554 ( .A1(n797), .A2(n796), .ZN(n821) );
  OR2_X1 U555 ( .A1(n810), .A2(n809), .ZN(n819) );
  XOR2_X1 U556 ( .A(KEYINPUT32), .B(n782), .Z(n809) );
  NOR2_X1 U557 ( .A1(G164), .A2(G1384), .ZN(n726) );
  NOR2_X1 U558 ( .A1(n527), .A2(G2105), .ZN(n621) );
  NOR2_X1 U559 ( .A1(n821), .A2(n820), .ZN(n520) );
  OR2_X1 U560 ( .A1(n520), .A2(n521), .ZN(n837) );
  OR2_X1 U561 ( .A1(n522), .A2(n822), .ZN(n521) );
  INV_X1 U562 ( .A(n844), .ZN(n522) );
  NAND2_X1 U563 ( .A1(n910), .A2(G138), .ZN(n525) );
  NOR2_X1 U564 ( .A1(n732), .A2(n997), .ZN(n734) );
  NOR2_X1 U565 ( .A1(n717), .A2(n716), .ZN(n724) );
  XNOR2_X1 U566 ( .A(n532), .B(KEYINPUT91), .ZN(G164) );
  OR2_X1 U567 ( .A1(n531), .A2(n530), .ZN(n532) );
  AND2_X1 U568 ( .A1(n724), .A2(G1996), .ZN(n725) );
  AND2_X1 U569 ( .A1(n726), .A2(n725), .ZN(n728) );
  INV_X1 U570 ( .A(KEYINPUT27), .ZN(n744) );
  XNOR2_X1 U571 ( .A(n744), .B(KEYINPUT101), .ZN(n745) );
  XNOR2_X1 U572 ( .A(n746), .B(n745), .ZN(n749) );
  NOR2_X1 U573 ( .A1(n787), .A2(n764), .ZN(n765) );
  NOR2_X1 U574 ( .A1(n769), .A2(n768), .ZN(n770) );
  OR2_X1 U575 ( .A1(n808), .A2(n817), .ZN(n810) );
  INV_X1 U576 ( .A(KEYINPUT17), .ZN(n523) );
  NOR2_X2 U577 ( .A1(G651), .A2(G543), .ZN(n660) );
  INV_X1 U578 ( .A(KEYINPUT109), .ZN(n836) );
  XNOR2_X1 U579 ( .A(n837), .B(n836), .ZN(n852) );
  XOR2_X1 U580 ( .A(G2104), .B(KEYINPUT66), .Z(n527) );
  AND2_X1 U581 ( .A1(G2105), .A2(n527), .ZN(n914) );
  NAND2_X1 U582 ( .A1(G126), .A2(n914), .ZN(n526) );
  NOR2_X1 U583 ( .A1(G2105), .A2(G2104), .ZN(n524) );
  XNOR2_X2 U584 ( .A(n524), .B(n523), .ZN(n910) );
  NAND2_X1 U585 ( .A1(n526), .A2(n525), .ZN(n531) );
  AND2_X1 U586 ( .A1(G2105), .A2(G2104), .ZN(n915) );
  NAND2_X1 U587 ( .A1(G114), .A2(n915), .ZN(n529) );
  NAND2_X1 U588 ( .A1(G102), .A2(n621), .ZN(n528) );
  NAND2_X1 U589 ( .A1(n529), .A2(n528), .ZN(n530) );
  NAND2_X1 U590 ( .A1(G90), .A2(n660), .ZN(n534) );
  XOR2_X1 U591 ( .A(G543), .B(KEYINPUT0), .Z(n643) );
  INV_X1 U592 ( .A(G651), .ZN(n537) );
  NOR2_X1 U593 ( .A1(n643), .A2(n537), .ZN(n664) );
  NAND2_X1 U594 ( .A1(G77), .A2(n664), .ZN(n533) );
  NAND2_X1 U595 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U596 ( .A(KEYINPUT9), .B(n535), .ZN(n542) );
  NOR2_X1 U597 ( .A1(G651), .A2(n643), .ZN(n536) );
  XOR2_X1 U598 ( .A(KEYINPUT65), .B(n536), .Z(n661) );
  NAND2_X1 U599 ( .A1(G52), .A2(n661), .ZN(n540) );
  NOR2_X1 U600 ( .A1(G543), .A2(n537), .ZN(n538) );
  NAND2_X1 U601 ( .A1(G64), .A2(n668), .ZN(n539) );
  AND2_X1 U602 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U603 ( .A1(n542), .A2(n541), .ZN(G301) );
  INV_X1 U604 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U605 ( .A(G2435), .B(G2443), .ZN(n552) );
  XOR2_X1 U606 ( .A(G2454), .B(G2430), .Z(n544) );
  XNOR2_X1 U607 ( .A(G2446), .B(KEYINPUT113), .ZN(n543) );
  XNOR2_X1 U608 ( .A(n544), .B(n543), .ZN(n548) );
  XOR2_X1 U609 ( .A(G2451), .B(G2427), .Z(n546) );
  XNOR2_X1 U610 ( .A(G1341), .B(G1348), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U612 ( .A(n548), .B(n547), .Z(n550) );
  XNOR2_X1 U613 ( .A(KEYINPUT112), .B(G2438), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U615 ( .A(n552), .B(n551), .ZN(n553) );
  AND2_X1 U616 ( .A1(n553), .A2(G14), .ZN(G401) );
  AND2_X1 U617 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U618 ( .A(G860), .ZN(n628) );
  NAND2_X1 U619 ( .A1(G81), .A2(n660), .ZN(n554) );
  XOR2_X1 U620 ( .A(KEYINPUT12), .B(n554), .Z(n555) );
  XNOR2_X1 U621 ( .A(n555), .B(KEYINPUT69), .ZN(n557) );
  NAND2_X1 U622 ( .A1(G68), .A2(n664), .ZN(n556) );
  NAND2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(KEYINPUT13), .ZN(n560) );
  NAND2_X1 U625 ( .A1(G43), .A2(n661), .ZN(n559) );
  NAND2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n563) );
  NAND2_X1 U627 ( .A1(n668), .A2(G56), .ZN(n561) );
  XOR2_X1 U628 ( .A(KEYINPUT14), .B(n561), .Z(n562) );
  NOR2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X2 U630 ( .A(KEYINPUT70), .B(n564), .Z(n997) );
  OR2_X1 U631 ( .A1(n628), .A2(n997), .ZN(G153) );
  NAND2_X1 U632 ( .A1(G53), .A2(n661), .ZN(n566) );
  NAND2_X1 U633 ( .A1(G65), .A2(n668), .ZN(n565) );
  NAND2_X1 U634 ( .A1(n566), .A2(n565), .ZN(n570) );
  NAND2_X1 U635 ( .A1(G91), .A2(n660), .ZN(n568) );
  NAND2_X1 U636 ( .A1(G78), .A2(n664), .ZN(n567) );
  NAND2_X1 U637 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X1 U638 ( .A1(n570), .A2(n569), .ZN(n753) );
  INV_X1 U639 ( .A(n753), .ZN(G299) );
  INV_X1 U640 ( .A(G57), .ZN(G237) );
  INV_X1 U641 ( .A(G132), .ZN(G219) );
  INV_X1 U642 ( .A(G82), .ZN(G220) );
  NAND2_X1 U643 ( .A1(G101), .A2(n621), .ZN(n571) );
  XNOR2_X1 U644 ( .A(n571), .B(KEYINPUT23), .ZN(n572) );
  XNOR2_X1 U645 ( .A(n572), .B(KEYINPUT67), .ZN(n575) );
  NAND2_X1 U646 ( .A1(G137), .A2(n910), .ZN(n573) );
  XNOR2_X1 U647 ( .A(n573), .B(KEYINPUT68), .ZN(n574) );
  NAND2_X1 U648 ( .A1(n575), .A2(n574), .ZN(n717) );
  NAND2_X1 U649 ( .A1(G125), .A2(n914), .ZN(n577) );
  NAND2_X1 U650 ( .A1(G113), .A2(n915), .ZN(n576) );
  NAND2_X1 U651 ( .A1(n577), .A2(n576), .ZN(n714) );
  NOR2_X1 U652 ( .A1(n717), .A2(n714), .ZN(G160) );
  NAND2_X1 U653 ( .A1(n668), .A2(G63), .ZN(n578) );
  XNOR2_X1 U654 ( .A(n578), .B(KEYINPUT76), .ZN(n580) );
  NAND2_X1 U655 ( .A1(G51), .A2(n661), .ZN(n579) );
  NAND2_X1 U656 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U657 ( .A(KEYINPUT6), .B(n581), .ZN(n589) );
  NAND2_X1 U658 ( .A1(G89), .A2(n660), .ZN(n582) );
  XNOR2_X1 U659 ( .A(n582), .B(KEYINPUT4), .ZN(n583) );
  XNOR2_X1 U660 ( .A(n583), .B(KEYINPUT74), .ZN(n585) );
  NAND2_X1 U661 ( .A1(G76), .A2(n664), .ZN(n584) );
  NAND2_X1 U662 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U663 ( .A(KEYINPUT5), .B(n586), .ZN(n587) );
  XNOR2_X1 U664 ( .A(KEYINPUT75), .B(n587), .ZN(n588) );
  NOR2_X1 U665 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U666 ( .A(n590), .B(KEYINPUT7), .ZN(n591) );
  XNOR2_X1 U667 ( .A(n591), .B(KEYINPUT77), .ZN(G168) );
  XOR2_X1 U668 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U669 ( .A1(G7), .A2(G661), .ZN(n592) );
  XNOR2_X1 U670 ( .A(n592), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U671 ( .A(G223), .ZN(n854) );
  NAND2_X1 U672 ( .A1(n854), .A2(G567), .ZN(n593) );
  XOR2_X1 U673 ( .A(KEYINPUT11), .B(n593), .Z(G234) );
  NAND2_X1 U674 ( .A1(G92), .A2(n660), .ZN(n595) );
  NAND2_X1 U675 ( .A1(G79), .A2(n664), .ZN(n594) );
  NAND2_X1 U676 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U677 ( .A1(G54), .A2(n661), .ZN(n597) );
  NAND2_X1 U678 ( .A1(G66), .A2(n668), .ZN(n596) );
  NAND2_X1 U679 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U680 ( .A1(n599), .A2(n598), .ZN(n601) );
  XNOR2_X1 U681 ( .A(KEYINPUT15), .B(KEYINPUT72), .ZN(n600) );
  XNOR2_X1 U682 ( .A(n601), .B(n600), .ZN(n602) );
  XNOR2_X1 U683 ( .A(KEYINPUT71), .B(n602), .ZN(n992) );
  NOR2_X1 U684 ( .A1(G868), .A2(n992), .ZN(n604) );
  INV_X1 U685 ( .A(G868), .ZN(n606) );
  NOR2_X1 U686 ( .A1(G171), .A2(n606), .ZN(n603) );
  NOR2_X1 U687 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U688 ( .A(KEYINPUT73), .B(n605), .ZN(G284) );
  NOR2_X1 U689 ( .A1(G286), .A2(n606), .ZN(n608) );
  NOR2_X1 U690 ( .A1(G868), .A2(G299), .ZN(n607) );
  NOR2_X1 U691 ( .A1(n608), .A2(n607), .ZN(G297) );
  NAND2_X1 U692 ( .A1(n628), .A2(G559), .ZN(n609) );
  NAND2_X1 U693 ( .A1(n609), .A2(n992), .ZN(n610) );
  XNOR2_X1 U694 ( .A(n610), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U695 ( .A1(n997), .A2(G868), .ZN(n613) );
  NAND2_X1 U696 ( .A1(n992), .A2(G868), .ZN(n611) );
  NOR2_X1 U697 ( .A1(G559), .A2(n611), .ZN(n612) );
  NOR2_X1 U698 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U699 ( .A(KEYINPUT78), .B(n614), .ZN(G282) );
  NAND2_X1 U700 ( .A1(n914), .A2(G123), .ZN(n615) );
  XNOR2_X1 U701 ( .A(n615), .B(KEYINPUT18), .ZN(n617) );
  NAND2_X1 U702 ( .A1(G135), .A2(n910), .ZN(n616) );
  NAND2_X1 U703 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U704 ( .A(n618), .B(KEYINPUT79), .ZN(n620) );
  NAND2_X1 U705 ( .A1(G111), .A2(n915), .ZN(n619) );
  NAND2_X1 U706 ( .A1(n620), .A2(n619), .ZN(n624) );
  BUF_X1 U707 ( .A(n621), .Z(n911) );
  NAND2_X1 U708 ( .A1(n911), .A2(G99), .ZN(n622) );
  XOR2_X1 U709 ( .A(KEYINPUT80), .B(n622), .Z(n623) );
  NOR2_X1 U710 ( .A1(n624), .A2(n623), .ZN(n938) );
  XNOR2_X1 U711 ( .A(G2096), .B(n938), .ZN(n626) );
  INV_X1 U712 ( .A(G2100), .ZN(n625) );
  NAND2_X1 U713 ( .A1(n626), .A2(n625), .ZN(G156) );
  NAND2_X1 U714 ( .A1(n992), .A2(G559), .ZN(n627) );
  XOR2_X1 U715 ( .A(n997), .B(n627), .Z(n679) );
  NAND2_X1 U716 ( .A1(n628), .A2(n679), .ZN(n636) );
  NAND2_X1 U717 ( .A1(G93), .A2(n660), .ZN(n630) );
  NAND2_X1 U718 ( .A1(G80), .A2(n664), .ZN(n629) );
  NAND2_X1 U719 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U720 ( .A1(G55), .A2(n661), .ZN(n631) );
  XNOR2_X1 U721 ( .A(KEYINPUT81), .B(n631), .ZN(n632) );
  NOR2_X1 U722 ( .A1(n633), .A2(n632), .ZN(n635) );
  NAND2_X1 U723 ( .A1(n668), .A2(G67), .ZN(n634) );
  AND2_X1 U724 ( .A1(n635), .A2(n634), .ZN(n673) );
  XOR2_X1 U725 ( .A(n636), .B(n673), .Z(G145) );
  NAND2_X1 U726 ( .A1(G651), .A2(G74), .ZN(n637) );
  XNOR2_X1 U727 ( .A(KEYINPUT83), .B(n637), .ZN(n640) );
  NAND2_X1 U728 ( .A1(n661), .A2(G49), .ZN(n638) );
  XOR2_X1 U729 ( .A(KEYINPUT82), .B(n638), .Z(n639) );
  NOR2_X1 U730 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U731 ( .A(KEYINPUT84), .B(n641), .Z(n642) );
  NOR2_X1 U732 ( .A1(n668), .A2(n642), .ZN(n645) );
  NAND2_X1 U733 ( .A1(n643), .A2(G87), .ZN(n644) );
  NAND2_X1 U734 ( .A1(n645), .A2(n644), .ZN(G288) );
  NAND2_X1 U735 ( .A1(G50), .A2(n661), .ZN(n647) );
  NAND2_X1 U736 ( .A1(G62), .A2(n668), .ZN(n646) );
  NAND2_X1 U737 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U738 ( .A(KEYINPUT85), .B(n648), .ZN(n653) );
  NAND2_X1 U739 ( .A1(G88), .A2(n660), .ZN(n650) );
  NAND2_X1 U740 ( .A1(G75), .A2(n664), .ZN(n649) );
  NAND2_X1 U741 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U742 ( .A(KEYINPUT86), .B(n651), .Z(n652) );
  NAND2_X1 U743 ( .A1(n653), .A2(n652), .ZN(G303) );
  INV_X1 U744 ( .A(G303), .ZN(G166) );
  AND2_X1 U745 ( .A1(n661), .A2(G47), .ZN(n657) );
  NAND2_X1 U746 ( .A1(G85), .A2(n660), .ZN(n655) );
  NAND2_X1 U747 ( .A1(G72), .A2(n664), .ZN(n654) );
  NAND2_X1 U748 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U749 ( .A1(n657), .A2(n656), .ZN(n659) );
  NAND2_X1 U750 ( .A1(n668), .A2(G60), .ZN(n658) );
  NAND2_X1 U751 ( .A1(n659), .A2(n658), .ZN(G290) );
  NAND2_X1 U752 ( .A1(G86), .A2(n660), .ZN(n663) );
  NAND2_X1 U753 ( .A1(G48), .A2(n661), .ZN(n662) );
  NAND2_X1 U754 ( .A1(n663), .A2(n662), .ZN(n667) );
  NAND2_X1 U755 ( .A1(n664), .A2(G73), .ZN(n665) );
  XOR2_X1 U756 ( .A(KEYINPUT2), .B(n665), .Z(n666) );
  NOR2_X1 U757 ( .A1(n667), .A2(n666), .ZN(n670) );
  NAND2_X1 U758 ( .A1(n668), .A2(G61), .ZN(n669) );
  NAND2_X1 U759 ( .A1(n670), .A2(n669), .ZN(G305) );
  NOR2_X1 U760 ( .A1(n673), .A2(G868), .ZN(n671) );
  XNOR2_X1 U761 ( .A(KEYINPUT89), .B(n671), .ZN(n683) );
  XOR2_X1 U762 ( .A(KEYINPUT87), .B(KEYINPUT19), .Z(n672) );
  XOR2_X1 U763 ( .A(n673), .B(n672), .Z(n674) );
  XNOR2_X1 U764 ( .A(G288), .B(n674), .ZN(n676) );
  XNOR2_X1 U765 ( .A(n753), .B(G166), .ZN(n675) );
  XNOR2_X1 U766 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U767 ( .A(n677), .B(G290), .ZN(n678) );
  XNOR2_X1 U768 ( .A(n678), .B(G305), .ZN(n860) );
  XNOR2_X1 U769 ( .A(n860), .B(n679), .ZN(n680) );
  NAND2_X1 U770 ( .A1(n680), .A2(G868), .ZN(n681) );
  XNOR2_X1 U771 ( .A(KEYINPUT88), .B(n681), .ZN(n682) );
  NAND2_X1 U772 ( .A1(n683), .A2(n682), .ZN(G295) );
  NAND2_X1 U773 ( .A1(G2084), .A2(G2078), .ZN(n684) );
  XOR2_X1 U774 ( .A(KEYINPUT20), .B(n684), .Z(n685) );
  NAND2_X1 U775 ( .A1(G2090), .A2(n685), .ZN(n686) );
  XNOR2_X1 U776 ( .A(KEYINPUT21), .B(n686), .ZN(n687) );
  NAND2_X1 U777 ( .A1(n687), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U778 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U779 ( .A1(G661), .A2(G483), .ZN(n695) );
  NOR2_X1 U780 ( .A1(G220), .A2(G219), .ZN(n688) );
  XOR2_X1 U781 ( .A(KEYINPUT22), .B(n688), .Z(n689) );
  NOR2_X1 U782 ( .A1(G218), .A2(n689), .ZN(n690) );
  NAND2_X1 U783 ( .A1(G96), .A2(n690), .ZN(n858) );
  NAND2_X1 U784 ( .A1(n858), .A2(G2106), .ZN(n694) );
  NAND2_X1 U785 ( .A1(G69), .A2(G120), .ZN(n691) );
  NOR2_X1 U786 ( .A1(G237), .A2(n691), .ZN(n692) );
  NAND2_X1 U787 ( .A1(G108), .A2(n692), .ZN(n859) );
  NAND2_X1 U788 ( .A1(n859), .A2(G567), .ZN(n693) );
  NAND2_X1 U789 ( .A1(n694), .A2(n693), .ZN(n934) );
  NOR2_X1 U790 ( .A1(n695), .A2(n934), .ZN(n696) );
  XNOR2_X1 U791 ( .A(n696), .B(KEYINPUT90), .ZN(n857) );
  NAND2_X1 U792 ( .A1(G36), .A2(n857), .ZN(G176) );
  NAND2_X1 U793 ( .A1(G107), .A2(n915), .ZN(n698) );
  NAND2_X1 U794 ( .A1(G95), .A2(n911), .ZN(n697) );
  NAND2_X1 U795 ( .A1(n698), .A2(n697), .ZN(n702) );
  NAND2_X1 U796 ( .A1(G119), .A2(n914), .ZN(n700) );
  NAND2_X1 U797 ( .A1(G131), .A2(n910), .ZN(n699) );
  NAND2_X1 U798 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U799 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U800 ( .A(n703), .B(KEYINPUT96), .Z(n892) );
  AND2_X1 U801 ( .A1(G1991), .A2(n892), .ZN(n713) );
  NAND2_X1 U802 ( .A1(G105), .A2(n911), .ZN(n704) );
  XOR2_X1 U803 ( .A(KEYINPUT38), .B(n704), .Z(n709) );
  NAND2_X1 U804 ( .A1(G129), .A2(n914), .ZN(n706) );
  NAND2_X1 U805 ( .A1(G117), .A2(n915), .ZN(n705) );
  NAND2_X1 U806 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U807 ( .A(KEYINPUT97), .B(n707), .Z(n708) );
  NOR2_X1 U808 ( .A1(n709), .A2(n708), .ZN(n711) );
  NAND2_X1 U809 ( .A1(n910), .A2(G141), .ZN(n710) );
  NAND2_X1 U810 ( .A1(n711), .A2(n710), .ZN(n893) );
  AND2_X1 U811 ( .A1(n893), .A2(G1996), .ZN(n712) );
  NOR2_X1 U812 ( .A1(n713), .A2(n712), .ZN(n946) );
  INV_X1 U813 ( .A(G40), .ZN(n715) );
  OR2_X1 U814 ( .A1(n715), .A2(n714), .ZN(n716) );
  INV_X1 U815 ( .A(n724), .ZN(n718) );
  NOR2_X1 U816 ( .A1(n726), .A2(n718), .ZN(n849) );
  XOR2_X1 U817 ( .A(n849), .B(KEYINPUT98), .Z(n719) );
  NOR2_X1 U818 ( .A1(n946), .A2(n719), .ZN(n840) );
  INV_X1 U819 ( .A(n840), .ZN(n721) );
  XNOR2_X1 U820 ( .A(G1986), .B(G290), .ZN(n994) );
  NAND2_X1 U821 ( .A1(n849), .A2(n994), .ZN(n720) );
  NAND2_X1 U822 ( .A1(n721), .A2(n720), .ZN(n822) );
  XOR2_X1 U823 ( .A(KEYINPUT25), .B(G2078), .Z(n961) );
  NAND2_X1 U824 ( .A1(n726), .A2(n724), .ZN(n772) );
  NOR2_X1 U825 ( .A1(n961), .A2(n772), .ZN(n723) );
  INV_X1 U826 ( .A(n772), .ZN(n747) );
  NOR2_X1 U827 ( .A1(n747), .A2(G1961), .ZN(n722) );
  NOR2_X1 U828 ( .A1(n723), .A2(n722), .ZN(n767) );
  NOR2_X1 U829 ( .A1(n767), .A2(G301), .ZN(n760) );
  INV_X1 U830 ( .A(G1996), .ZN(n960) );
  XOR2_X1 U831 ( .A(KEYINPUT26), .B(KEYINPUT102), .Z(n727) );
  XNOR2_X1 U832 ( .A(n728), .B(n727), .ZN(n730) );
  NAND2_X1 U833 ( .A1(n772), .A2(G1341), .ZN(n729) );
  NAND2_X1 U834 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U835 ( .A(KEYINPUT103), .B(n731), .Z(n732) );
  INV_X1 U836 ( .A(KEYINPUT64), .ZN(n733) );
  XNOR2_X1 U837 ( .A(n734), .B(n733), .ZN(n741) );
  INV_X1 U838 ( .A(n992), .ZN(n861) );
  OR2_X1 U839 ( .A1(n741), .A2(n861), .ZN(n740) );
  NAND2_X1 U840 ( .A1(G2067), .A2(n747), .ZN(n735) );
  XNOR2_X1 U841 ( .A(n735), .B(KEYINPUT104), .ZN(n737) );
  NAND2_X1 U842 ( .A1(G1348), .A2(n772), .ZN(n736) );
  NAND2_X1 U843 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U844 ( .A(KEYINPUT105), .B(n738), .Z(n739) );
  NAND2_X1 U845 ( .A1(n740), .A2(n739), .ZN(n743) );
  NAND2_X1 U846 ( .A1(n861), .A2(n741), .ZN(n742) );
  NAND2_X1 U847 ( .A1(n743), .A2(n742), .ZN(n751) );
  NAND2_X1 U848 ( .A1(G2072), .A2(n747), .ZN(n746) );
  INV_X1 U849 ( .A(G1956), .ZN(n1010) );
  NOR2_X1 U850 ( .A1(n747), .A2(n1010), .ZN(n748) );
  NOR2_X1 U851 ( .A1(n749), .A2(n748), .ZN(n752) );
  NAND2_X1 U852 ( .A1(n753), .A2(n752), .ZN(n750) );
  NAND2_X1 U853 ( .A1(n751), .A2(n750), .ZN(n756) );
  NOR2_X1 U854 ( .A1(n753), .A2(n752), .ZN(n754) );
  XOR2_X1 U855 ( .A(n754), .B(KEYINPUT28), .Z(n755) );
  NAND2_X1 U856 ( .A1(n756), .A2(n755), .ZN(n758) );
  XNOR2_X1 U857 ( .A(KEYINPUT29), .B(KEYINPUT106), .ZN(n757) );
  XNOR2_X1 U858 ( .A(n758), .B(n757), .ZN(n759) );
  NOR2_X1 U859 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U860 ( .A(n761), .B(KEYINPUT107), .ZN(n784) );
  NAND2_X1 U861 ( .A1(n772), .A2(G8), .ZN(n762) );
  XOR2_X1 U862 ( .A(KEYINPUT99), .B(n762), .Z(n792) );
  NOR2_X1 U863 ( .A1(G1966), .A2(n792), .ZN(n787) );
  NOR2_X1 U864 ( .A1(G2084), .A2(n772), .ZN(n763) );
  XOR2_X1 U865 ( .A(KEYINPUT100), .B(n763), .Z(n785) );
  NAND2_X1 U866 ( .A1(G8), .A2(n785), .ZN(n764) );
  XOR2_X1 U867 ( .A(KEYINPUT30), .B(n765), .Z(n766) );
  NOR2_X1 U868 ( .A1(G168), .A2(n766), .ZN(n769) );
  AND2_X1 U869 ( .A1(G301), .A2(n767), .ZN(n768) );
  XOR2_X1 U870 ( .A(n770), .B(KEYINPUT31), .Z(n771) );
  XNOR2_X1 U871 ( .A(n771), .B(KEYINPUT108), .ZN(n783) );
  NOR2_X1 U872 ( .A1(G1971), .A2(n792), .ZN(n774) );
  NOR2_X1 U873 ( .A1(G2090), .A2(n772), .ZN(n773) );
  NOR2_X1 U874 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U875 ( .A1(n775), .A2(G303), .ZN(n777) );
  AND2_X1 U876 ( .A1(n783), .A2(n777), .ZN(n776) );
  NAND2_X1 U877 ( .A1(n784), .A2(n776), .ZN(n781) );
  INV_X1 U878 ( .A(n777), .ZN(n778) );
  OR2_X1 U879 ( .A1(n778), .A2(G286), .ZN(n779) );
  AND2_X1 U880 ( .A1(G8), .A2(n779), .ZN(n780) );
  NAND2_X1 U881 ( .A1(n781), .A2(n780), .ZN(n782) );
  AND2_X1 U882 ( .A1(n784), .A2(n783), .ZN(n791) );
  INV_X1 U883 ( .A(n785), .ZN(n786) );
  NAND2_X1 U884 ( .A1(G8), .A2(n786), .ZN(n789) );
  INV_X1 U885 ( .A(n787), .ZN(n788) );
  NAND2_X1 U886 ( .A1(n789), .A2(n788), .ZN(n790) );
  NOR2_X1 U887 ( .A1(n791), .A2(n790), .ZN(n808) );
  INV_X1 U888 ( .A(n792), .ZN(n801) );
  OR2_X1 U889 ( .A1(n808), .A2(n801), .ZN(n793) );
  NOR2_X1 U890 ( .A1(n809), .A2(n793), .ZN(n797) );
  NAND2_X1 U891 ( .A1(G166), .A2(G8), .ZN(n794) );
  NOR2_X1 U892 ( .A1(G2090), .A2(n794), .ZN(n795) );
  AND2_X1 U893 ( .A1(n792), .A2(n795), .ZN(n796) );
  NOR2_X1 U894 ( .A1(G1981), .A2(G305), .ZN(n798) );
  XNOR2_X1 U895 ( .A(n798), .B(KEYINPUT24), .ZN(n799) );
  NAND2_X1 U896 ( .A1(n799), .A2(n801), .ZN(n814) );
  INV_X1 U897 ( .A(n814), .ZN(n807) );
  NAND2_X1 U898 ( .A1(G1976), .A2(G288), .ZN(n989) );
  AND2_X1 U899 ( .A1(n801), .A2(n989), .ZN(n800) );
  NOR2_X1 U900 ( .A1(KEYINPUT33), .A2(n800), .ZN(n805) );
  NOR2_X1 U901 ( .A1(G1976), .A2(G288), .ZN(n988) );
  AND2_X1 U902 ( .A1(n988), .A2(KEYINPUT33), .ZN(n802) );
  AND2_X1 U903 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U904 ( .A(G1981), .B(G305), .ZN(n986) );
  OR2_X1 U905 ( .A1(n803), .A2(n986), .ZN(n804) );
  NOR2_X1 U906 ( .A1(n805), .A2(n804), .ZN(n806) );
  NOR2_X1 U907 ( .A1(n807), .A2(n806), .ZN(n817) );
  NOR2_X1 U908 ( .A1(G1971), .A2(G303), .ZN(n811) );
  NOR2_X1 U909 ( .A1(n988), .A2(n811), .ZN(n813) );
  INV_X1 U910 ( .A(KEYINPUT33), .ZN(n812) );
  AND2_X1 U911 ( .A1(n813), .A2(n812), .ZN(n815) );
  AND2_X1 U912 ( .A1(n815), .A2(n814), .ZN(n816) );
  OR2_X1 U913 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U914 ( .A1(n819), .A2(n818), .ZN(n820) );
  XOR2_X1 U915 ( .A(G2067), .B(KEYINPUT37), .Z(n846) );
  NAND2_X1 U916 ( .A1(n910), .A2(G140), .ZN(n823) );
  XNOR2_X1 U917 ( .A(KEYINPUT93), .B(n823), .ZN(n826) );
  NAND2_X1 U918 ( .A1(n911), .A2(G104), .ZN(n824) );
  XOR2_X1 U919 ( .A(n824), .B(KEYINPUT92), .Z(n825) );
  NOR2_X1 U920 ( .A1(n826), .A2(n825), .ZN(n827) );
  XOR2_X1 U921 ( .A(KEYINPUT95), .B(n827), .Z(n829) );
  XOR2_X1 U922 ( .A(KEYINPUT34), .B(KEYINPUT94), .Z(n828) );
  XNOR2_X1 U923 ( .A(n829), .B(n828), .ZN(n834) );
  NAND2_X1 U924 ( .A1(G128), .A2(n914), .ZN(n831) );
  NAND2_X1 U925 ( .A1(G116), .A2(n915), .ZN(n830) );
  NAND2_X1 U926 ( .A1(n831), .A2(n830), .ZN(n832) );
  XOR2_X1 U927 ( .A(KEYINPUT35), .B(n832), .Z(n833) );
  NOR2_X1 U928 ( .A1(n834), .A2(n833), .ZN(n835) );
  XOR2_X1 U929 ( .A(KEYINPUT36), .B(n835), .Z(n894) );
  AND2_X1 U930 ( .A1(n846), .A2(n894), .ZN(n944) );
  NAND2_X1 U931 ( .A1(n849), .A2(n944), .ZN(n844) );
  NOR2_X1 U932 ( .A1(G1996), .A2(n893), .ZN(n936) );
  NOR2_X1 U933 ( .A1(G1986), .A2(G290), .ZN(n838) );
  NOR2_X1 U934 ( .A1(G1991), .A2(n892), .ZN(n939) );
  NOR2_X1 U935 ( .A1(n838), .A2(n939), .ZN(n839) );
  NOR2_X1 U936 ( .A1(n840), .A2(n839), .ZN(n841) );
  XNOR2_X1 U937 ( .A(n841), .B(KEYINPUT110), .ZN(n842) );
  NOR2_X1 U938 ( .A1(n936), .A2(n842), .ZN(n843) );
  XNOR2_X1 U939 ( .A(n843), .B(KEYINPUT39), .ZN(n845) );
  NAND2_X1 U940 ( .A1(n845), .A2(n844), .ZN(n848) );
  NOR2_X1 U941 ( .A1(n894), .A2(n846), .ZN(n847) );
  XNOR2_X1 U942 ( .A(n847), .B(KEYINPUT111), .ZN(n953) );
  NAND2_X1 U943 ( .A1(n848), .A2(n953), .ZN(n850) );
  NAND2_X1 U944 ( .A1(n850), .A2(n849), .ZN(n851) );
  NAND2_X1 U945 ( .A1(n852), .A2(n851), .ZN(n853) );
  XNOR2_X1 U946 ( .A(n853), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U947 ( .A1(G2106), .A2(n854), .ZN(G217) );
  AND2_X1 U948 ( .A1(G15), .A2(G2), .ZN(n855) );
  NAND2_X1 U949 ( .A1(G661), .A2(n855), .ZN(G259) );
  NAND2_X1 U950 ( .A1(G3), .A2(G1), .ZN(n856) );
  NAND2_X1 U951 ( .A1(n857), .A2(n856), .ZN(G188) );
  INV_X1 U953 ( .A(G120), .ZN(G236) );
  INV_X1 U954 ( .A(G96), .ZN(G221) );
  INV_X1 U955 ( .A(G69), .ZN(G235) );
  NOR2_X1 U956 ( .A1(n859), .A2(n858), .ZN(G325) );
  INV_X1 U957 ( .A(G325), .ZN(G261) );
  XOR2_X1 U958 ( .A(n860), .B(G286), .Z(n863) );
  XNOR2_X1 U959 ( .A(G171), .B(n861), .ZN(n862) );
  XNOR2_X1 U960 ( .A(n863), .B(n862), .ZN(n864) );
  XNOR2_X1 U961 ( .A(n997), .B(n864), .ZN(n865) );
  NOR2_X1 U962 ( .A1(G37), .A2(n865), .ZN(G397) );
  XOR2_X1 U963 ( .A(G2096), .B(KEYINPUT43), .Z(n867) );
  XNOR2_X1 U964 ( .A(G2090), .B(KEYINPUT114), .ZN(n866) );
  XNOR2_X1 U965 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U966 ( .A(n868), .B(G2678), .Z(n870) );
  XNOR2_X1 U967 ( .A(G2067), .B(G2072), .ZN(n869) );
  XNOR2_X1 U968 ( .A(n870), .B(n869), .ZN(n874) );
  XOR2_X1 U969 ( .A(KEYINPUT42), .B(G2100), .Z(n872) );
  XNOR2_X1 U970 ( .A(G2084), .B(G2078), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n872), .B(n871), .ZN(n873) );
  XNOR2_X1 U972 ( .A(n874), .B(n873), .ZN(G227) );
  XOR2_X1 U973 ( .A(G1976), .B(G1971), .Z(n876) );
  XNOR2_X1 U974 ( .A(G1961), .B(G1956), .ZN(n875) );
  XNOR2_X1 U975 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U976 ( .A(n877), .B(G2474), .Z(n879) );
  XNOR2_X1 U977 ( .A(G1996), .B(G1991), .ZN(n878) );
  XNOR2_X1 U978 ( .A(n879), .B(n878), .ZN(n883) );
  XOR2_X1 U979 ( .A(KEYINPUT41), .B(G1981), .Z(n881) );
  XNOR2_X1 U980 ( .A(G1986), .B(G1966), .ZN(n880) );
  XNOR2_X1 U981 ( .A(n881), .B(n880), .ZN(n882) );
  XNOR2_X1 U982 ( .A(n883), .B(n882), .ZN(G229) );
  NAND2_X1 U983 ( .A1(G112), .A2(n915), .ZN(n885) );
  NAND2_X1 U984 ( .A1(G100), .A2(n911), .ZN(n884) );
  NAND2_X1 U985 ( .A1(n885), .A2(n884), .ZN(n891) );
  NAND2_X1 U986 ( .A1(G124), .A2(n914), .ZN(n886) );
  XNOR2_X1 U987 ( .A(n886), .B(KEYINPUT44), .ZN(n889) );
  NAND2_X1 U988 ( .A1(G136), .A2(n910), .ZN(n887) );
  XOR2_X1 U989 ( .A(KEYINPUT115), .B(n887), .Z(n888) );
  NAND2_X1 U990 ( .A1(n889), .A2(n888), .ZN(n890) );
  NOR2_X1 U991 ( .A1(n891), .A2(n890), .ZN(G162) );
  XOR2_X1 U992 ( .A(n938), .B(n892), .Z(n896) );
  XOR2_X1 U993 ( .A(n894), .B(n893), .Z(n895) );
  XNOR2_X1 U994 ( .A(n896), .B(n895), .ZN(n900) );
  XOR2_X1 U995 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n898) );
  XNOR2_X1 U996 ( .A(G160), .B(G162), .ZN(n897) );
  XNOR2_X1 U997 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U998 ( .A(n900), .B(n899), .Z(n926) );
  NAND2_X1 U999 ( .A1(n915), .A2(G118), .ZN(n901) );
  XNOR2_X1 U1000 ( .A(n901), .B(KEYINPUT116), .ZN(n903) );
  NAND2_X1 U1001 ( .A1(G130), .A2(n914), .ZN(n902) );
  NAND2_X1 U1002 ( .A1(n903), .A2(n902), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n904), .B(KEYINPUT117), .ZN(n909) );
  NAND2_X1 U1004 ( .A1(G142), .A2(n910), .ZN(n906) );
  NAND2_X1 U1005 ( .A1(G106), .A2(n911), .ZN(n905) );
  NAND2_X1 U1006 ( .A1(n906), .A2(n905), .ZN(n907) );
  XNOR2_X1 U1007 ( .A(KEYINPUT45), .B(n907), .ZN(n908) );
  NAND2_X1 U1008 ( .A1(n909), .A2(n908), .ZN(n923) );
  NAND2_X1 U1009 ( .A1(G139), .A2(n910), .ZN(n913) );
  NAND2_X1 U1010 ( .A1(G103), .A2(n911), .ZN(n912) );
  NAND2_X1 U1011 ( .A1(n913), .A2(n912), .ZN(n921) );
  NAND2_X1 U1012 ( .A1(G127), .A2(n914), .ZN(n917) );
  NAND2_X1 U1013 ( .A1(G115), .A2(n915), .ZN(n916) );
  NAND2_X1 U1014 ( .A1(n917), .A2(n916), .ZN(n918) );
  XOR2_X1 U1015 ( .A(KEYINPUT118), .B(n918), .Z(n919) );
  XNOR2_X1 U1016 ( .A(KEYINPUT47), .B(n919), .ZN(n920) );
  NOR2_X1 U1017 ( .A1(n921), .A2(n920), .ZN(n922) );
  XOR2_X1 U1018 ( .A(KEYINPUT119), .B(n922), .Z(n947) );
  XNOR2_X1 U1019 ( .A(n923), .B(n947), .ZN(n924) );
  XNOR2_X1 U1020 ( .A(G164), .B(n924), .ZN(n925) );
  XNOR2_X1 U1021 ( .A(n926), .B(n925), .ZN(n927) );
  NOR2_X1 U1022 ( .A1(G37), .A2(n927), .ZN(G395) );
  NOR2_X1 U1023 ( .A1(G227), .A2(G229), .ZN(n928) );
  XNOR2_X1 U1024 ( .A(KEYINPUT49), .B(n928), .ZN(n929) );
  NOR2_X1 U1025 ( .A1(G397), .A2(n929), .ZN(n933) );
  NOR2_X1 U1026 ( .A1(n934), .A2(G401), .ZN(n930) );
  XOR2_X1 U1027 ( .A(KEYINPUT120), .B(n930), .Z(n931) );
  NOR2_X1 U1028 ( .A1(G395), .A2(n931), .ZN(n932) );
  NAND2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(G225) );
  INV_X1 U1030 ( .A(G225), .ZN(G308) );
  INV_X1 U1031 ( .A(n934), .ZN(G319) );
  INV_X1 U1032 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1033 ( .A(G2090), .B(G162), .Z(n935) );
  NOR2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1035 ( .A(KEYINPUT51), .B(n937), .Z(n942) );
  NOR2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1037 ( .A(KEYINPUT121), .B(n940), .Z(n941) );
  NAND2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n956) );
  XOR2_X1 U1039 ( .A(G160), .B(G2084), .Z(n943) );
  NOR2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n952) );
  XOR2_X1 U1042 ( .A(G2072), .B(n947), .Z(n949) );
  XOR2_X1 U1043 ( .A(G164), .B(G2078), .Z(n948) );
  NOR2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1045 ( .A(KEYINPUT50), .B(n950), .Z(n951) );
  NOR2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n954) );
  NAND2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1048 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1049 ( .A(KEYINPUT52), .B(n957), .ZN(n958) );
  XOR2_X1 U1050 ( .A(KEYINPUT55), .B(KEYINPUT122), .Z(n981) );
  NAND2_X1 U1051 ( .A1(n958), .A2(n981), .ZN(n959) );
  NAND2_X1 U1052 ( .A1(n959), .A2(G29), .ZN(n1039) );
  XOR2_X1 U1053 ( .A(KEYINPUT125), .B(KEYINPUT53), .Z(n974) );
  XNOR2_X1 U1054 ( .A(G32), .B(n960), .ZN(n965) );
  XNOR2_X1 U1055 ( .A(n961), .B(G27), .ZN(n963) );
  XNOR2_X1 U1056 ( .A(G2072), .B(G33), .ZN(n962) );
  NOR2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n968) );
  XOR2_X1 U1059 ( .A(KEYINPUT123), .B(G2067), .Z(n966) );
  XNOR2_X1 U1060 ( .A(G26), .B(n966), .ZN(n967) );
  NOR2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1062 ( .A(KEYINPUT124), .B(n969), .Z(n971) );
  XNOR2_X1 U1063 ( .A(G1991), .B(G25), .ZN(n970) );
  NOR2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1065 ( .A1(n972), .A2(G28), .ZN(n973) );
  XNOR2_X1 U1066 ( .A(n974), .B(n973), .ZN(n979) );
  XNOR2_X1 U1067 ( .A(G2084), .B(G34), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(n975), .B(KEYINPUT54), .ZN(n977) );
  XNOR2_X1 U1069 ( .A(G35), .B(G2090), .ZN(n976) );
  NOR2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1072 ( .A(n981), .B(n980), .ZN(n983) );
  INV_X1 U1073 ( .A(G29), .ZN(n982) );
  NAND2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1075 ( .A1(G11), .A2(n984), .ZN(n1037) );
  XNOR2_X1 U1076 ( .A(G16), .B(KEYINPUT56), .ZN(n1009) );
  XOR2_X1 U1077 ( .A(G168), .B(G1966), .Z(n985) );
  NOR2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1079 ( .A(KEYINPUT57), .B(n987), .Z(n1007) );
  INV_X1 U1080 ( .A(n988), .ZN(n990) );
  NAND2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n1005) );
  XNOR2_X1 U1082 ( .A(G1971), .B(G166), .ZN(n991) );
  XNOR2_X1 U1083 ( .A(n991), .B(KEYINPUT126), .ZN(n1003) );
  XNOR2_X1 U1084 ( .A(G1348), .B(n992), .ZN(n996) );
  XNOR2_X1 U1085 ( .A(G1956), .B(G299), .ZN(n993) );
  NOR2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n1001) );
  XOR2_X1 U1088 ( .A(n997), .B(G1341), .Z(n999) );
  XNOR2_X1 U1089 ( .A(G171), .B(G1961), .ZN(n998) );
  NAND2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NOR2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1035) );
  INV_X1 U1096 ( .A(G16), .ZN(n1033) );
  XNOR2_X1 U1097 ( .A(G20), .B(n1010), .ZN(n1014) );
  XNOR2_X1 U1098 ( .A(G1341), .B(G19), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(G6), .B(G1981), .ZN(n1011) );
  NOR2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1017) );
  XOR2_X1 U1102 ( .A(KEYINPUT59), .B(G1348), .Z(n1015) );
  XNOR2_X1 U1103 ( .A(G4), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1019) );
  XOR2_X1 U1105 ( .A(KEYINPUT127), .B(KEYINPUT60), .Z(n1018) );
  XNOR2_X1 U1106 ( .A(n1019), .B(n1018), .ZN(n1023) );
  XNOR2_X1 U1107 ( .A(G1966), .B(G21), .ZN(n1021) );
  XNOR2_X1 U1108 ( .A(G1961), .B(G5), .ZN(n1020) );
  NOR2_X1 U1109 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1030) );
  XNOR2_X1 U1111 ( .A(G1986), .B(G24), .ZN(n1025) );
  XNOR2_X1 U1112 ( .A(G1971), .B(G22), .ZN(n1024) );
  NOR2_X1 U1113 ( .A1(n1025), .A2(n1024), .ZN(n1027) );
  XOR2_X1 U1114 ( .A(G1976), .B(G23), .Z(n1026) );
  NAND2_X1 U1115 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1116 ( .A(KEYINPUT58), .B(n1028), .ZN(n1029) );
  NOR2_X1 U1117 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1118 ( .A(KEYINPUT61), .B(n1031), .ZN(n1032) );
  NAND2_X1 U1119 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1120 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NOR2_X1 U1121 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NAND2_X1 U1122 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  XOR2_X1 U1123 ( .A(KEYINPUT62), .B(n1040), .Z(G311) );
  INV_X1 U1124 ( .A(G311), .ZN(G150) );
endmodule

