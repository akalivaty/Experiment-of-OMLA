//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 1 0 1 1 0 0 1 0 0 0 1 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 0 0 1 1 1 0 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n603,
    new_n604, new_n605, new_n606, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n648, new_n649, new_n650, new_n653,
    new_n655, new_n656, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1217, new_n1218, new_n1219;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT65), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  XOR2_X1   g030(.A(G325), .B(KEYINPUT66), .Z(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  NAND2_X1  g032(.A1(G113), .A2(G2104), .ZN(new_n458));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G125), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n458), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(new_n466), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n465), .A2(new_n472), .ZN(G160));
  OAI21_X1  g048(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(G112), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n474), .B1(new_n475), .B2(G2105), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n461), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(KEYINPUT67), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n470), .A2(new_n479), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n461), .A2(new_n466), .ZN(new_n483));
  AOI211_X1 g058(.A(new_n476), .B(new_n482), .C1(G124), .C2(new_n483), .ZN(G162));
  OAI211_X1 g059(.A(G138), .B(new_n466), .C1(new_n459), .C2(new_n460), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT4), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n487), .A2(new_n466), .A3(G138), .ZN(new_n488));
  NOR3_X1   g063(.A1(new_n461), .A2(KEYINPUT69), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT69), .ZN(new_n490));
  AND3_X1   g065(.A1(new_n487), .A2(new_n466), .A3(G138), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(new_n469), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n486), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n494), .B1(new_n495), .B2(G2105), .ZN(new_n496));
  AND2_X1   g071(.A1(G126), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(new_n459), .B2(new_n460), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT68), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g075(.A(KEYINPUT68), .B(new_n497), .C1(new_n459), .C2(new_n460), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n496), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n493), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  NAND2_X1  g079(.A1(G75), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n506), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n509), .B1(new_n506), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  NOR3_X1   g086(.A1(new_n511), .A2(KEYINPUT70), .A3(KEYINPUT5), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n508), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G62), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n505), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n517), .A2(new_n511), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n515), .A2(G651), .B1(G50), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g094(.A(KEYINPUT71), .B1(new_n513), .B2(new_n517), .ZN(new_n520));
  OAI21_X1  g095(.A(KEYINPUT70), .B1(new_n511), .B2(KEYINPUT5), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n509), .A2(new_n506), .A3(G543), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n507), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT71), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(new_n524), .A3(new_n516), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT72), .B(G88), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n520), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n519), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(G166));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT75), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n523), .A2(G63), .A3(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n520), .A2(new_n525), .ZN(new_n534));
  INV_X1    g109(.A(G89), .ZN(new_n535));
  OAI211_X1 g110(.A(new_n532), .B(new_n533), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT74), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT73), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n511), .B1(new_n516), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(KEYINPUT6), .A2(G651), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(KEYINPUT6), .A2(G651), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n541), .A2(KEYINPUT73), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n537), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n542), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n538), .B1(new_n545), .B2(new_n540), .ZN(new_n546));
  AND4_X1   g121(.A1(new_n537), .A2(new_n543), .A3(new_n546), .A4(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(G51), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n536), .A2(new_n550), .ZN(G168));
  NAND2_X1  g126(.A1(new_n521), .A2(new_n522), .ZN(new_n552));
  AND4_X1   g127(.A1(new_n524), .A2(new_n552), .A3(new_n508), .A4(new_n516), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n524), .B1(new_n523), .B2(new_n516), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G90), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G651), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  XOR2_X1   g135(.A(KEYINPUT76), .B(G52), .Z(new_n561));
  OAI21_X1  g136(.A(new_n561), .B1(new_n544), .B2(new_n547), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n560), .A2(new_n563), .ZN(G171));
  INV_X1    g139(.A(KEYINPUT78), .ZN(new_n565));
  OAI21_X1  g140(.A(G43), .B1(new_n544), .B2(new_n547), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n520), .A2(G81), .A3(new_n525), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT77), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n523), .A2(G56), .ZN(new_n570));
  NAND2_X1  g145(.A1(G68), .A2(G543), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n571), .ZN(new_n573));
  AOI211_X1 g148(.A(KEYINPUT77), .B(new_n573), .C1(new_n523), .C2(G56), .ZN(new_n574));
  NOR3_X1   g149(.A1(new_n572), .A2(new_n574), .A3(new_n558), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n565), .B1(new_n568), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n570), .A2(new_n571), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(KEYINPUT77), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n570), .A2(new_n569), .A3(new_n571), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n578), .A2(G651), .A3(new_n579), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n580), .A2(KEYINPUT78), .A3(new_n566), .A4(new_n567), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(G860), .ZN(G153));
  NAND4_X1  g159(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g160(.A(KEYINPUT79), .B(KEYINPUT8), .Z(new_n586));
  NAND2_X1  g161(.A1(G1), .A2(G3), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n586), .B(new_n587), .ZN(new_n588));
  NAND4_X1  g163(.A1(G319), .A2(G483), .A3(G661), .A4(new_n588), .ZN(G188));
  NAND4_X1  g164(.A1(new_n543), .A2(new_n546), .A3(G53), .A4(G543), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(KEYINPUT9), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT9), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n539), .A2(new_n592), .A3(G53), .A4(new_n543), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n520), .A2(G91), .A3(new_n525), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n523), .A2(G65), .ZN(new_n596));
  NAND2_X1  g171(.A1(G78), .A2(G543), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G651), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n594), .A2(new_n595), .A3(new_n599), .ZN(G299));
  INV_X1    g175(.A(G171), .ZN(G301));
  INV_X1    g176(.A(G168), .ZN(G286));
  INV_X1    g177(.A(KEYINPUT80), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n519), .A2(new_n603), .A3(new_n527), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n603), .B1(new_n519), .B2(new_n527), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n605), .A2(new_n606), .ZN(G303));
  AND2_X1   g182(.A1(new_n555), .A2(G87), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n539), .A2(G49), .A3(new_n543), .ZN(new_n609));
  OAI21_X1  g184(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(G288));
  NAND2_X1  g188(.A1(G73), .A2(G543), .ZN(new_n614));
  INV_X1    g189(.A(G61), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n513), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n616), .A2(KEYINPUT81), .A3(G651), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT81), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n523), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n558), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n520), .A2(G86), .A3(new_n525), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n516), .A2(G48), .A3(G543), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT82), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND4_X1  g199(.A1(new_n617), .A2(new_n620), .A3(new_n621), .A4(new_n624), .ZN(G305));
  INV_X1    g200(.A(new_n548), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G47), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n555), .A2(G85), .ZN(new_n628));
  AOI22_X1  g203(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n629), .A2(new_n558), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n627), .A2(new_n628), .A3(new_n630), .ZN(G290));
  INV_X1    g206(.A(G868), .ZN(new_n632));
  NOR2_X1   g207(.A1(G171), .A2(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(KEYINPUT83), .ZN(new_n634));
  NAND2_X1  g209(.A1(G79), .A2(G543), .ZN(new_n635));
  INV_X1    g210(.A(G66), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n513), .B2(new_n636), .ZN(new_n637));
  AOI22_X1  g212(.A1(new_n626), .A2(G54), .B1(G651), .B2(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(KEYINPUT10), .ZN(new_n639));
  INV_X1    g214(.A(G92), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n639), .B1(new_n534), .B2(new_n640), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n555), .A2(KEYINPUT10), .A3(G92), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  AOI22_X1  g219(.A1(new_n633), .A2(new_n634), .B1(new_n644), .B2(new_n632), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(new_n634), .B2(new_n633), .ZN(G284));
  OAI21_X1  g221(.A(new_n645), .B1(new_n634), .B2(new_n633), .ZN(G321));
  OR3_X1    g222(.A1(G168), .A2(KEYINPUT84), .A3(new_n632), .ZN(new_n648));
  OAI21_X1  g223(.A(KEYINPUT84), .B1(G168), .B2(new_n632), .ZN(new_n649));
  INV_X1    g224(.A(G299), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n648), .B(new_n649), .C1(G868), .C2(new_n650), .ZN(G297));
  OAI211_X1 g226(.A(new_n648), .B(new_n649), .C1(G868), .C2(new_n650), .ZN(G280));
  INV_X1    g227(.A(G559), .ZN(new_n653));
  OAI211_X1 g228(.A(new_n638), .B(new_n643), .C1(new_n653), .C2(G860), .ZN(G148));
  NAND3_X1  g229(.A1(new_n638), .A2(new_n653), .A3(new_n643), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(G868), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n656), .B1(new_n583), .B2(G868), .ZN(G323));
  XNOR2_X1  g232(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g233(.A1(new_n469), .A2(new_n467), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT12), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT85), .B(KEYINPUT13), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n662), .A2(G2100), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n483), .A2(G123), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n466), .A2(G111), .ZN(new_n665));
  OAI21_X1  g240(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n478), .A2(new_n480), .ZN(new_n667));
  INV_X1    g242(.A(G135), .ZN(new_n668));
  OAI221_X1 g243(.A(new_n664), .B1(new_n665), .B2(new_n666), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n669), .A2(G2096), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n662), .A2(G2100), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(G2096), .ZN(new_n672));
  NAND4_X1  g247(.A1(new_n663), .A2(new_n670), .A3(new_n671), .A4(new_n672), .ZN(G156));
  INV_X1    g248(.A(KEYINPUT14), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2427), .B(G2438), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G2430), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT15), .B(G2435), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n674), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n678), .B1(new_n677), .B2(new_n676), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2451), .B(G2454), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT16), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1341), .B(G1348), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n679), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G2443), .B(G2446), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G14), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n684), .A2(new_n685), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(G401));
  XOR2_X1   g264(.A(G2084), .B(G2090), .Z(new_n690));
  XNOR2_X1  g265(.A(G2067), .B(G2678), .ZN(new_n691));
  XNOR2_X1  g266(.A(G2072), .B(G2078), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT86), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT18), .Z(new_n695));
  INV_X1    g270(.A(new_n690), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n691), .B(KEYINPUT87), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n692), .B(KEYINPUT88), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n696), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT89), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n692), .B(KEYINPUT17), .Z(new_n702));
  OAI22_X1  g277(.A1(new_n700), .A2(new_n701), .B1(new_n697), .B2(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n701), .B2(new_n700), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n698), .A2(new_n696), .ZN(new_n705));
  AOI211_X1 g280(.A(new_n695), .B(new_n704), .C1(new_n702), .C2(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(G2096), .B(G2100), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(G227));
  XNOR2_X1  g283(.A(G1971), .B(G1976), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(G1956), .B(G2474), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1961), .B(G1966), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n712), .A2(new_n713), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n711), .A2(KEYINPUT91), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n717), .B(new_n718), .Z(new_n719));
  NOR3_X1   g294(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT20), .Z(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(G1991), .B(G1996), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(G1981), .B(G1986), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(G229));
  INV_X1    g303(.A(G16), .ZN(new_n729));
  NOR2_X1   g304(.A1(G171), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G5), .B2(new_n729), .ZN(new_n731));
  INV_X1    g306(.A(G1961), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G29), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT24), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(G34), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n735), .B2(G34), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G160), .B2(G29), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n467), .A2(G105), .ZN(new_n739));
  NAND3_X1  g314(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT26), .ZN(new_n741));
  AOI211_X1 g316(.A(new_n739), .B(new_n741), .C1(G129), .C2(new_n483), .ZN(new_n742));
  INV_X1    g317(.A(G141), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(new_n743), .B2(new_n667), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT98), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(KEYINPUT99), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n744), .B(KEYINPUT98), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT99), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n734), .B1(new_n747), .B2(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n734), .B2(G32), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT27), .B(G1996), .ZN(new_n753));
  OAI221_X1 g328(.A(new_n733), .B1(G2084), .B2(new_n738), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT101), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n481), .A2(KEYINPUT97), .A3(G139), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT97), .ZN(new_n757));
  INV_X1    g332(.A(G139), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n757), .B1(new_n667), .B2(new_n758), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT25), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(new_n466), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n760), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(G29), .ZN(new_n767));
  NOR2_X1   g342(.A1(G29), .A2(G33), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT96), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n767), .A2(G2072), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(G29), .A2(G35), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G162), .B2(G29), .ZN(new_n772));
  XOR2_X1   g347(.A(KEYINPUT104), .B(KEYINPUT29), .Z(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n770), .B1(new_n774), .B2(G2090), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT95), .B(KEYINPUT28), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n734), .A2(G26), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n481), .A2(G140), .ZN(new_n779));
  OAI21_X1  g354(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n780));
  INV_X1    g355(.A(G116), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n780), .B1(new_n781), .B2(G2105), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n483), .B2(G128), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n778), .B1(new_n784), .B2(G29), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G2067), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n669), .A2(new_n734), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n787), .A2(KEYINPUT100), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G2084), .B2(new_n738), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n787), .A2(KEYINPUT100), .ZN(new_n790));
  INV_X1    g365(.A(G28), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n791), .A2(KEYINPUT30), .ZN(new_n792));
  AOI21_X1  g367(.A(G29), .B1(new_n791), .B2(KEYINPUT30), .ZN(new_n793));
  OR2_X1    g368(.A1(KEYINPUT31), .A2(G11), .ZN(new_n794));
  NAND2_X1  g369(.A1(KEYINPUT31), .A2(G11), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n792), .A2(new_n793), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n786), .A2(new_n789), .A3(new_n790), .A4(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(G2072), .B1(new_n767), .B2(new_n769), .ZN(new_n798));
  NOR3_X1   g373(.A1(new_n775), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n583), .A2(new_n729), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n729), .B2(G19), .ZN(new_n801));
  INV_X1    g376(.A(G1341), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n801), .A2(new_n802), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n734), .A2(G27), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT102), .Z(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n503), .B2(G29), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT103), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G2078), .ZN(new_n809));
  INV_X1    g384(.A(new_n731), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n809), .B1(G1961), .B2(new_n810), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n799), .A2(new_n803), .A3(new_n804), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n752), .A2(new_n753), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n729), .A2(G21), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(G168), .B2(new_n729), .ZN(new_n815));
  INV_X1    g390(.A(G1966), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  MUX2_X1   g392(.A(G4), .B(new_n644), .S(G16), .Z(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(G1348), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n818), .A2(G1348), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n813), .A2(new_n817), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  NOR3_X1   g396(.A1(new_n755), .A2(new_n812), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n729), .A2(G23), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(new_n612), .B2(new_n729), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT33), .B(G1976), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n729), .A2(G22), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(G166), .B2(new_n729), .ZN(new_n828));
  INV_X1    g403(.A(G1971), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  MUX2_X1   g405(.A(G6), .B(G305), .S(G16), .Z(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT32), .B(G1981), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n826), .A2(new_n830), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n835), .A2(KEYINPUT34), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(KEYINPUT34), .ZN(new_n837));
  NOR2_X1   g412(.A1(G16), .A2(G24), .ZN(new_n838));
  INV_X1    g413(.A(G290), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n838), .B1(new_n839), .B2(G16), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(G1986), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n840), .A2(G1986), .ZN(new_n842));
  NOR2_X1   g417(.A1(G25), .A2(G29), .ZN(new_n843));
  OR2_X1    g418(.A1(G95), .A2(G2105), .ZN(new_n844));
  OAI211_X1 g419(.A(new_n844), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT92), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n846), .B1(G119), .B2(new_n483), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n481), .A2(G131), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n843), .B1(new_n850), .B2(G29), .ZN(new_n851));
  XNOR2_X1  g426(.A(KEYINPUT35), .B(G1991), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT93), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n851), .B(new_n853), .ZN(new_n854));
  AND3_X1   g429(.A1(new_n842), .A2(KEYINPUT94), .A3(new_n854), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n836), .A2(new_n837), .A3(new_n841), .A4(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT36), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n856), .A2(new_n857), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n774), .A2(G2090), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n729), .A2(G20), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT23), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n862), .B1(new_n650), .B2(new_n729), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(KEYINPUT105), .Z(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(G1956), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n864), .A2(G1956), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n860), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT106), .ZN(new_n868));
  NAND4_X1  g443(.A1(new_n822), .A2(new_n858), .A3(new_n859), .A4(new_n868), .ZN(G150));
  INV_X1    g444(.A(G150), .ZN(G311));
  NOR2_X1   g445(.A1(new_n644), .A2(new_n653), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT38), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT107), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n555), .A2(G93), .ZN(new_n874));
  OAI21_X1  g449(.A(G55), .B1(new_n544), .B2(new_n547), .ZN(new_n875));
  AOI22_X1  g450(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n874), .B(new_n875), .C1(new_n558), .C2(new_n876), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n576), .A2(new_n873), .A3(new_n581), .A4(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n877), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n580), .A2(new_n566), .A3(new_n567), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n576), .A2(new_n581), .A3(new_n877), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(KEYINPUT107), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n872), .B(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT39), .ZN(new_n887));
  AOI21_X1  g462(.A(G860), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n888), .B1(new_n887), .B2(new_n886), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT108), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n877), .A2(G860), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n891), .B(KEYINPUT37), .Z(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(G145));
  XNOR2_X1  g468(.A(new_n669), .B(G160), .ZN(new_n894));
  XNOR2_X1  g469(.A(G162), .B(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n748), .A2(new_n749), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n746), .A2(KEYINPUT99), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n766), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n784), .A2(KEYINPUT109), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n784), .A2(KEYINPUT109), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n503), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n902), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(G164), .A3(new_n900), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n748), .A2(new_n766), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n899), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n903), .A2(new_n905), .ZN(new_n910));
  INV_X1    g485(.A(new_n766), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n911), .B1(new_n747), .B2(new_n750), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n910), .B1(new_n912), .B2(new_n907), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n849), .B(new_n660), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n483), .A2(G130), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n466), .A2(G118), .ZN(new_n916));
  OAI21_X1  g491(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n917));
  INV_X1    g492(.A(G142), .ZN(new_n918));
  OAI221_X1 g493(.A(new_n915), .B1(new_n916), .B2(new_n917), .C1(new_n667), .C2(new_n918), .ZN(new_n919));
  XOR2_X1   g494(.A(new_n914), .B(new_n919), .Z(new_n920));
  AND3_X1   g495(.A1(new_n909), .A2(new_n913), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n920), .B1(new_n909), .B2(new_n913), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n896), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n920), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n912), .A2(new_n910), .A3(new_n907), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n906), .B1(new_n899), .B2(new_n908), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n909), .A2(new_n913), .A3(new_n920), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n927), .A2(new_n895), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(G37), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n923), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(KEYINPUT110), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT110), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n923), .A2(new_n929), .A3(new_n933), .A4(new_n930), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n935), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g511(.A(new_n885), .B(new_n655), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n644), .B(new_n650), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(KEYINPUT41), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n937), .A2(new_n938), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT42), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n528), .B(KEYINPUT111), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n839), .B(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n612), .B(G305), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n944), .B(new_n945), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n946), .A2(KEYINPUT112), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n937), .A2(new_n939), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT42), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n948), .B(new_n949), .C1(new_n938), .C2(new_n937), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n942), .A2(new_n947), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n947), .B1(new_n942), .B2(new_n950), .ZN(new_n952));
  OAI21_X1  g527(.A(G868), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n953), .B1(G868), .B2(new_n879), .ZN(G295));
  OAI21_X1  g529(.A(new_n953), .B1(G868), .B2(new_n879), .ZN(G331));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n956));
  XOR2_X1   g531(.A(new_n938), .B(KEYINPUT41), .Z(new_n957));
  AND2_X1   g532(.A1(new_n883), .A2(KEYINPUT107), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n878), .A2(new_n881), .ZN(new_n959));
  OAI21_X1  g534(.A(G168), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n884), .A2(G286), .A3(new_n881), .A4(new_n878), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n960), .A2(G171), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(G171), .B1(new_n960), .B2(new_n961), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n957), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(G286), .B1(new_n882), .B2(new_n884), .ZN(new_n965));
  INV_X1    g540(.A(new_n961), .ZN(new_n966));
  OAI21_X1  g541(.A(G301), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n960), .A2(G171), .A3(new_n961), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n967), .A2(new_n938), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n964), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(G37), .B1(new_n970), .B2(new_n946), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n972));
  INV_X1    g547(.A(new_n946), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n964), .A2(new_n969), .A3(new_n973), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n971), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n972), .B1(new_n971), .B2(new_n974), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n956), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n970), .A2(new_n946), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n978), .A2(new_n930), .A3(new_n974), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT43), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n971), .A2(new_n972), .A3(new_n974), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n980), .A2(KEYINPUT44), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n977), .A2(new_n982), .ZN(G397));
  XOR2_X1   g558(.A(KEYINPUT113), .B(G1384), .Z(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT45), .B1(new_n503), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n477), .A2(G137), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n464), .A2(new_n988), .A3(G40), .A4(new_n468), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(G290), .A2(G1986), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(KEYINPUT114), .ZN(new_n992));
  INV_X1    g567(.A(G1986), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n992), .B1(new_n993), .B2(new_n839), .ZN(new_n994));
  INV_X1    g569(.A(G1996), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n747), .A2(new_n750), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n784), .A2(G2067), .ZN(new_n997));
  INV_X1    g572(.A(G2067), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n779), .A2(new_n998), .A3(new_n783), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n1000), .B1(new_n748), .B2(G1996), .ZN(new_n1001));
  OR2_X1    g576(.A1(new_n850), .A2(new_n853), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n850), .A2(new_n853), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n996), .A2(new_n1001), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n990), .B1(new_n994), .B2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n1005), .B(KEYINPUT115), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n558), .B1(new_n596), .B2(new_n597), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1007), .B1(new_n555), .B2(G91), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1008), .B(new_n594), .C1(KEYINPUT120), .C2(KEYINPUT57), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n595), .A2(new_n599), .A3(KEYINPUT120), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT57), .ZN(new_n1011));
  NAND3_X1  g586(.A1(G299), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1956), .ZN(new_n1014));
  INV_X1    g589(.A(new_n989), .ZN(new_n1015));
  AOI21_X1  g590(.A(G1384), .B1(new_n493), .B2(new_n502), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT50), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1384), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT69), .B1(new_n461), .B2(new_n488), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n469), .A2(new_n491), .A3(new_n490), .ZN(new_n1021));
  AOI22_X1  g596(.A1(new_n1020), .A2(new_n1021), .B1(KEYINPUT4), .B2(new_n485), .ZN(new_n1022));
  INV_X1    g597(.A(new_n496), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT68), .B1(new_n469), .B2(new_n497), .ZN(new_n1024));
  INV_X1    g599(.A(new_n501), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1023), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1019), .B1(new_n1022), .B2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1027), .A2(KEYINPUT50), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1014), .B1(new_n1018), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT45), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n989), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n985), .ZN(new_n1032));
  XNOR2_X1  g607(.A(KEYINPUT56), .B(G2072), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1013), .B1(new_n1029), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1348), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1036), .B1(new_n1018), .B2(new_n1028), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1027), .A2(new_n989), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n998), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n644), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1013), .A2(new_n1029), .A3(new_n1034), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1035), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT61), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1013), .A2(new_n1029), .A3(new_n1034), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1043), .B1(new_n1044), .B2(new_n1035), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1037), .A2(new_n644), .A3(new_n1039), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT60), .B1(new_n1046), .B2(new_n1040), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n644), .A2(KEYINPUT60), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1048), .A2(new_n1039), .A3(new_n1037), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1029), .A2(new_n1034), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1052), .A2(KEYINPUT61), .A3(new_n1041), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1045), .A2(new_n1047), .A3(new_n1049), .A4(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1031), .A2(new_n995), .A3(new_n1032), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1038), .ZN(new_n1056));
  XOR2_X1   g631(.A(KEYINPUT58), .B(G1341), .Z(new_n1057));
  AOI22_X1  g632(.A1(new_n1055), .A2(KEYINPUT121), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT121), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1031), .A2(new_n1059), .A3(new_n995), .A4(new_n1032), .ZN(new_n1060));
  AOI211_X1 g635(.A(KEYINPUT59), .B(new_n582), .C1(new_n1058), .C2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT59), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1055), .A2(KEYINPUT121), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1063), .A2(new_n1060), .A3(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1062), .B1(new_n1065), .B2(new_n583), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1061), .A2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1042), .B1(new_n1054), .B2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(G303), .A2(KEYINPUT117), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n528), .A2(KEYINPUT80), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1070), .A2(KEYINPUT55), .A3(G8), .A4(new_n604), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT117), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1070), .A2(G8), .A3(new_n604), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT55), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1069), .A2(new_n1073), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT116), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1015), .B1(new_n1016), .B2(KEYINPUT45), .ZN(new_n1079));
  AOI211_X1 g654(.A(new_n1030), .B(new_n984), .C1(new_n493), .C2(new_n502), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1078), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1031), .A2(KEYINPUT116), .A3(new_n1032), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1081), .A2(new_n1082), .A3(new_n829), .ZN(new_n1083));
  OR3_X1    g658(.A1(new_n1018), .A2(new_n1028), .A3(G2090), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(G8), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1077), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT49), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT118), .B(G86), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n520), .A2(new_n525), .A3(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n617), .A2(new_n620), .A3(new_n1090), .A4(new_n624), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1091), .A2(G1981), .ZN(new_n1092));
  NOR2_X1   g667(.A1(G305), .A2(G1981), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1088), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1091), .A2(G1981), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1095), .B(KEYINPUT49), .C1(G1981), .C2(G305), .ZN(new_n1096));
  INV_X1    g671(.A(G8), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1097), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1094), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n555), .A2(G87), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1100), .A2(G1976), .A3(new_n610), .A4(new_n609), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n1098), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT52), .ZN(new_n1103));
  INV_X1    g678(.A(G1976), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(new_n608), .B2(new_n611), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT52), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1105), .A2(new_n1101), .A3(new_n1098), .A4(new_n1106), .ZN(new_n1107));
  AND2_X1   g682(.A1(new_n1103), .A2(new_n1107), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1099), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1097), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1069), .A2(new_n1073), .A3(new_n1076), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1087), .A2(new_n1109), .A3(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(G8), .B1(new_n536), .B2(new_n550), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n816), .B1(new_n1079), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n989), .B1(new_n1027), .B2(KEYINPUT50), .ZN(new_n1117));
  INV_X1    g692(.A(G2084), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1114), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n1018), .A2(new_n1028), .A3(G2084), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1016), .A2(KEYINPUT45), .ZN(new_n1123));
  AOI21_X1  g698(.A(G1966), .B1(new_n1031), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(G8), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT51), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1126), .B1(new_n1114), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1125), .A2(new_n1129), .A3(new_n1114), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1097), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1114), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1128), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1121), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT54), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1135), .B1(new_n560), .B2(new_n563), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n556), .A2(KEYINPUT54), .A3(new_n562), .A4(new_n559), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1139));
  INV_X1    g714(.A(G2078), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT53), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1140), .A2(KEYINPUT53), .ZN(new_n1144));
  NOR3_X1   g719(.A1(new_n1079), .A2(new_n1115), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(G1961), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT123), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n732), .B1(new_n1018), .B2(new_n1028), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT123), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1031), .A2(new_n1123), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1148), .B(new_n1149), .C1(new_n1150), .C2(new_n1144), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1147), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1138), .B1(new_n1143), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n989), .A2(new_n1144), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1032), .A2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1154), .B1(new_n1156), .B2(new_n986), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n987), .A2(KEYINPUT124), .A3(new_n1032), .A4(new_n1155), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1138), .A2(new_n1157), .A3(new_n1158), .A4(new_n1148), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1159), .B1(new_n1142), .B2(new_n1141), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n1134), .A2(new_n1153), .A3(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1068), .A2(new_n1113), .A3(new_n1161), .ZN(new_n1162));
  OAI211_X1 g737(.A(G8), .B(G168), .C1(new_n1122), .C2(new_n1124), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(KEYINPUT119), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT119), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1131), .A2(new_n1165), .A3(G168), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1087), .A2(new_n1167), .A3(new_n1109), .A4(new_n1112), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT63), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1099), .A2(new_n1108), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1171), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1172), .A2(KEYINPUT63), .A3(new_n1087), .A4(new_n1167), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1170), .A2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1112), .A2(new_n1171), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1099), .A2(new_n1104), .A3(new_n612), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1176), .B1(G1981), .B2(G305), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1175), .B1(new_n1177), .B2(new_n1098), .ZN(new_n1178));
  AND3_X1   g753(.A1(new_n1162), .A2(new_n1174), .A3(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT62), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1134), .A2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g756(.A(G301), .B1(new_n1143), .B2(new_n1152), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1113), .A2(KEYINPUT125), .A3(new_n1181), .A4(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT125), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1182), .A2(new_n1087), .A3(new_n1109), .A4(new_n1112), .ZN(new_n1185));
  AOI211_X1 g760(.A(KEYINPUT62), .B(new_n1121), .C1(new_n1130), .C2(new_n1133), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1184), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  OR2_X1    g762(.A1(new_n1134), .A2(new_n1180), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1183), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1006), .B1(new_n1179), .B2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g765(.A(KEYINPUT46), .B1(new_n990), .B2(new_n995), .ZN(new_n1191));
  XOR2_X1   g766(.A(new_n1191), .B(KEYINPUT126), .Z(new_n1192));
  INV_X1    g767(.A(KEYINPUT46), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n746), .B1(new_n1193), .B2(G1996), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n990), .B1(new_n1194), .B2(new_n1000), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1192), .A2(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g771(.A(new_n1196), .B(KEYINPUT47), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT48), .ZN(new_n1198));
  INV_X1    g773(.A(new_n990), .ZN(new_n1199));
  OR3_X1    g774(.A1(new_n992), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1004), .A2(new_n990), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1198), .B1(new_n992), .B2(new_n1199), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n996), .A2(new_n1001), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n999), .B1(new_n1204), .B2(new_n1003), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1205), .A2(new_n990), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1197), .A2(new_n1203), .A3(new_n1206), .ZN(new_n1207));
  OAI21_X1  g782(.A(KEYINPUT127), .B1(new_n1190), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g783(.A(KEYINPUT127), .ZN(new_n1209));
  INV_X1    g784(.A(new_n1207), .ZN(new_n1210));
  INV_X1    g785(.A(new_n1189), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1162), .A2(new_n1174), .A3(new_n1178), .ZN(new_n1212));
  NOR2_X1   g787(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  OAI211_X1 g788(.A(new_n1209), .B(new_n1210), .C1(new_n1213), .C2(new_n1006), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1208), .A2(new_n1214), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g790(.A(G319), .B1(new_n687), .B2(new_n688), .ZN(new_n1217));
  OR2_X1    g791(.A1(G227), .A2(new_n1217), .ZN(new_n1218));
  NOR2_X1   g792(.A1(G229), .A2(new_n1218), .ZN(new_n1219));
  OAI211_X1 g793(.A(new_n935), .B(new_n1219), .C1(new_n975), .C2(new_n976), .ZN(G225));
  INV_X1    g794(.A(G225), .ZN(G308));
endmodule


