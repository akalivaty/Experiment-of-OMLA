//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 1 1 1 0 1 1 0 0 0 1 1 1 1 0 0 1 0 0 1 0 1 0 0 1 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G210), .B1(G237), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  XNOR2_X1  g005(.A(G110), .B(G122), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(G116), .B(G119), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT5), .ZN(new_n195));
  INV_X1    g009(.A(G113), .ZN(new_n196));
  INV_X1    g010(.A(G116), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(KEYINPUT5), .ZN(new_n198));
  INV_X1    g012(.A(G119), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n196), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT2), .B(G113), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  AOI22_X1  g016(.A1(new_n195), .A2(new_n200), .B1(new_n202), .B2(new_n194), .ZN(new_n203));
  INV_X1    g017(.A(G104), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT3), .B1(new_n204), .B2(G107), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n206));
  INV_X1    g020(.A(G107), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(G104), .ZN(new_n208));
  INV_X1    g022(.A(G101), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n204), .A2(G107), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n205), .A2(new_n208), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n204), .A2(G107), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n207), .A2(G104), .ZN(new_n213));
  OAI211_X1 g027(.A(KEYINPUT83), .B(G101), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT83), .ZN(new_n215));
  XNOR2_X1  g029(.A(G104), .B(G107), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n215), .B1(new_n216), .B2(new_n209), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n203), .A2(new_n211), .A3(new_n214), .A4(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n195), .A2(new_n200), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n202), .A2(new_n194), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n217), .A2(new_n211), .A3(new_n214), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n193), .B1(new_n224), .B2(KEYINPUT8), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n205), .A2(new_n208), .A3(new_n210), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G101), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(KEYINPUT4), .A3(new_n211), .ZN(new_n228));
  INV_X1    g042(.A(new_n194), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(new_n201), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(new_n220), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT4), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n226), .A2(new_n232), .A3(G101), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n228), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(new_n218), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT8), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n224), .A2(new_n236), .ZN(new_n237));
  AOI22_X1  g051(.A1(new_n225), .A2(new_n235), .B1(new_n237), .B2(new_n193), .ZN(new_n238));
  INV_X1    g052(.A(G128), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(KEYINPUT1), .ZN(new_n240));
  INV_X1    g054(.A(G146), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G143), .ZN(new_n242));
  INV_X1    g056(.A(G143), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G146), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n240), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n243), .A2(KEYINPUT1), .A3(G146), .ZN(new_n246));
  XNOR2_X1  g060(.A(G143), .B(G146), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n245), .B(new_n246), .C1(G128), .C2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G125), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(KEYINPUT0), .A2(G128), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  XOR2_X1   g066(.A(KEYINPUT0), .B(G128), .Z(new_n253));
  OAI21_X1  g067(.A(new_n252), .B1(new_n253), .B2(new_n247), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n250), .B1(new_n255), .B2(new_n249), .ZN(new_n256));
  INV_X1    g070(.A(G953), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G224), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n258), .A2(KEYINPUT7), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n256), .B(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n191), .B1(new_n238), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n235), .A2(new_n193), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n234), .A2(new_n218), .A3(new_n192), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n262), .A2(KEYINPUT87), .A3(KEYINPUT6), .A4(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n256), .B(new_n258), .ZN(new_n265));
  NAND2_X1  g079(.A1(KEYINPUT87), .A2(KEYINPUT6), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n235), .A2(new_n193), .A3(new_n266), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n264), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n190), .B1(new_n261), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n260), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n225), .A2(new_n235), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n192), .B1(new_n224), .B2(new_n236), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n264), .A2(new_n265), .A3(new_n267), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n273), .A2(new_n191), .A3(new_n189), .A4(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n188), .B1(new_n269), .B2(new_n275), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n257), .A2(G952), .ZN(new_n277));
  INV_X1    g091(.A(G234), .ZN(new_n278));
  INV_X1    g092(.A(G237), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  AOI211_X1 g095(.A(new_n191), .B(new_n257), .C1(G234), .C2(G237), .ZN(new_n282));
  XNOR2_X1  g096(.A(KEYINPUT21), .B(G898), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n276), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(G116), .B(G122), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n207), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT93), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n288), .B(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(G128), .B(G143), .ZN(new_n291));
  INV_X1    g105(.A(G134), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n291), .B(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT14), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n287), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n197), .A2(KEYINPUT14), .A3(G122), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n295), .A2(G107), .A3(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n290), .A2(new_n293), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n291), .A2(KEYINPUT13), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n243), .A2(G128), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n299), .B(G134), .C1(KEYINPUT13), .C2(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n287), .B(new_n207), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n291), .A2(new_n292), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n298), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT9), .B(G234), .ZN(new_n306));
  INV_X1    g120(.A(G217), .ZN(new_n307));
  NOR3_X1   g121(.A1(new_n306), .A2(new_n307), .A3(G953), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n298), .A2(new_n308), .A3(new_n304), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(KEYINPUT94), .A3(new_n191), .ZN(new_n313));
  INV_X1    g127(.A(G478), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n314), .A2(KEYINPUT15), .ZN(new_n315));
  XOR2_X1   g129(.A(new_n313), .B(new_n315), .Z(new_n316));
  XNOR2_X1  g130(.A(G113), .B(G122), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n317), .B(new_n204), .ZN(new_n318));
  INV_X1    g132(.A(G140), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G125), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n249), .A2(G140), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(KEYINPUT16), .ZN(new_n322));
  OR3_X1    g136(.A1(new_n249), .A2(KEYINPUT16), .A3(G140), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n241), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n322), .A2(new_n323), .A3(G146), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G131), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT68), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n329), .A2(G237), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n279), .A2(KEYINPUT68), .ZN(new_n331));
  OAI211_X1 g145(.A(G214), .B(new_n257), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n243), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n279), .A2(KEYINPUT68), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n329), .A2(G237), .ZN(new_n335));
  AOI21_X1  g149(.A(G953), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n336), .A2(G143), .A3(G214), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n328), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n327), .B1(new_n338), .B2(KEYINPUT17), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n333), .A2(new_n328), .A3(new_n337), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT90), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n333), .A2(new_n337), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G131), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT90), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n333), .A2(new_n344), .A3(new_n337), .A4(new_n328), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n341), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n339), .B1(new_n346), .B2(KEYINPUT17), .ZN(new_n347));
  XNOR2_X1  g161(.A(G125), .B(G140), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n348), .A2(KEYINPUT79), .A3(new_n241), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT79), .B1(new_n348), .B2(new_n241), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n348), .A2(new_n241), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n338), .A2(KEYINPUT88), .A3(KEYINPUT18), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT88), .B1(new_n338), .B2(KEYINPUT18), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n354), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT18), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n333), .B(new_n337), .C1(new_n359), .C2(new_n328), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n360), .B(KEYINPUT89), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n318), .B(new_n347), .C1(new_n358), .C2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n342), .A2(KEYINPUT18), .A3(G131), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT88), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n355), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT89), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n360), .B(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n369), .A3(new_n354), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n318), .B1(new_n370), .B2(new_n347), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n191), .B1(new_n363), .B2(new_n371), .ZN(new_n372));
  XOR2_X1   g186(.A(KEYINPUT92), .B(G475), .Z(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n353), .B1(new_n366), .B2(new_n355), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n322), .A2(G146), .A3(new_n323), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n348), .B(KEYINPUT19), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n376), .B1(new_n377), .B2(new_n241), .ZN(new_n378));
  AOI22_X1  g192(.A1(new_n375), .A2(new_n369), .B1(new_n346), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n362), .B1(new_n379), .B2(new_n318), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT20), .ZN(new_n381));
  NOR2_X1   g195(.A1(G475), .A2(G902), .ZN(new_n382));
  XOR2_X1   g196(.A(new_n382), .B(KEYINPUT91), .Z(new_n383));
  AND3_X1   g197(.A1(new_n380), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n381), .B1(new_n380), .B2(new_n383), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n316), .B(new_n374), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n286), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(G221), .B1(new_n306), .B2(G902), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n388), .B(KEYINPUT82), .ZN(new_n389));
  INV_X1    g203(.A(G469), .ZN(new_n390));
  XNOR2_X1  g204(.A(G110), .B(G140), .ZN(new_n391));
  INV_X1    g205(.A(G227), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n392), .A2(G953), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n391), .B(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n240), .A2(new_n242), .A3(new_n244), .ZN(new_n396));
  AOI21_X1  g210(.A(G128), .B1(new_n242), .B2(new_n244), .ZN(new_n397));
  INV_X1    g211(.A(new_n246), .ZN(new_n398));
  NOR3_X1   g212(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(KEYINPUT84), .B1(new_n222), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(KEYINPUT10), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n248), .A2(new_n211), .A3(new_n214), .A4(new_n217), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT10), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(KEYINPUT84), .A3(new_n403), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n254), .A2(new_n233), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n228), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n401), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT11), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n408), .B1(new_n292), .B2(G137), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n292), .A2(G137), .ZN(new_n410));
  INV_X1    g224(.A(G137), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(KEYINPUT11), .A3(G134), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n409), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(KEYINPUT65), .B1(new_n413), .B2(G131), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n413), .A2(KEYINPUT65), .A3(G131), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n409), .A2(new_n412), .A3(new_n328), .A4(new_n410), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT64), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n416), .A2(new_n417), .ZN(new_n419));
  OAI22_X1  g233(.A1(new_n414), .A2(new_n415), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT85), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n407), .A2(new_n422), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n400), .A2(KEYINPUT10), .B1(new_n405), .B2(new_n228), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(new_n404), .A3(new_n421), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n395), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n413), .A2(G131), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT65), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n413), .A2(KEYINPUT65), .A3(G131), .ZN(new_n430));
  AND2_X1   g244(.A1(new_n412), .A2(new_n410), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n431), .A2(KEYINPUT64), .A3(new_n328), .A4(new_n409), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n416), .A2(new_n417), .ZN(new_n433));
  AOI22_X1  g247(.A1(new_n429), .A2(new_n430), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n401), .A2(new_n434), .A3(new_n404), .A4(new_n406), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n222), .A2(new_n399), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n402), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n420), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT12), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT12), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n437), .A2(new_n440), .A3(new_n420), .ZN(new_n441));
  AND4_X1   g255(.A1(new_n435), .A2(new_n439), .A3(new_n441), .A4(new_n395), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n390), .B(new_n191), .C1(new_n426), .C2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(KEYINPUT86), .ZN(new_n444));
  AND4_X1   g258(.A1(new_n404), .A2(new_n421), .A3(new_n401), .A4(new_n406), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n421), .B1(new_n424), .B2(new_n404), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n394), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n435), .A2(new_n439), .A3(new_n441), .A4(new_n395), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT86), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n449), .A2(new_n450), .A3(new_n390), .A4(new_n191), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n444), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n435), .A2(new_n439), .A3(new_n441), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n394), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n423), .A2(new_n395), .A3(new_n425), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n390), .B1(new_n456), .B2(new_n191), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n389), .B1(new_n452), .B2(new_n458), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n387), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n336), .A2(G210), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT27), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT26), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT27), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n336), .A2(new_n464), .A3(G210), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n462), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n463), .B1(new_n462), .B2(new_n465), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n209), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n468), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(G101), .A3(new_n466), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT28), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT71), .ZN(new_n474));
  INV_X1    g288(.A(new_n410), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n292), .A2(G137), .ZN(new_n476));
  OAI21_X1  g290(.A(G131), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n477), .B(new_n248), .C1(new_n418), .C2(new_n419), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n474), .B(new_n478), .C1(new_n434), .C2(new_n255), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT67), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n231), .B(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n415), .A2(new_n414), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n416), .B(KEYINPUT64), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n254), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n474), .B1(new_n485), .B2(new_n478), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n473), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT72), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT72), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n489), .B(new_n473), .C1(new_n482), .C2(new_n486), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT66), .ZN(new_n492));
  NOR3_X1   g306(.A1(new_n434), .A2(new_n492), .A3(new_n255), .ZN(new_n493));
  AOI21_X1  g307(.A(KEYINPUT66), .B1(new_n420), .B2(new_n254), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n478), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n231), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n481), .A2(new_n485), .A3(new_n478), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n473), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n472), .B1(new_n491), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT69), .ZN(new_n500));
  OAI211_X1 g314(.A(KEYINPUT30), .B(new_n478), .C1(new_n434), .C2(new_n255), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n231), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT30), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n502), .B1(new_n495), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n497), .A2(new_n471), .A3(new_n469), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n500), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n505), .ZN(new_n507));
  INV_X1    g321(.A(new_n478), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n492), .B1(new_n434), .B2(new_n255), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n420), .A2(KEYINPUT66), .A3(new_n254), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n511), .A2(KEYINPUT30), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n507), .B(KEYINPUT69), .C1(new_n512), .C2(new_n502), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n506), .A2(KEYINPUT31), .A3(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT70), .B(KEYINPUT31), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n507), .B(new_n515), .C1(new_n512), .C2(new_n502), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n499), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(G472), .A2(G902), .ZN(new_n518));
  AOI21_X1  g332(.A(KEYINPUT32), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n231), .B(KEYINPUT67), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n434), .A2(new_n255), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n521), .B1(new_n522), .B2(new_n508), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n523), .A2(KEYINPUT73), .A3(new_n497), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT73), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n485), .A2(new_n481), .A3(new_n525), .A4(new_n478), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n524), .A2(KEYINPUT28), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT29), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n472), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n527), .A2(new_n488), .A3(new_n490), .A4(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT74), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n530), .B(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n231), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n497), .B1(new_n511), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT28), .ZN(new_n535));
  INV_X1    g349(.A(new_n472), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n535), .A2(new_n488), .A3(new_n490), .A4(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n497), .B1(new_n512), .B2(new_n502), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n472), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n537), .A2(new_n528), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n191), .ZN(new_n541));
  OAI21_X1  g355(.A(G472), .B1(new_n532), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n517), .A2(KEYINPUT32), .A3(new_n518), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n520), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT81), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n326), .B1(new_n349), .B2(new_n350), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT75), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n547), .B1(new_n199), .B2(G128), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT23), .ZN(new_n549));
  INV_X1    g363(.A(G110), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT23), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n547), .B(new_n551), .C1(new_n199), .C2(G128), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n199), .A2(G128), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n549), .A2(new_n550), .A3(new_n552), .A4(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n239), .A2(G119), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n553), .ZN(new_n556));
  XNOR2_X1  g370(.A(KEYINPUT24), .B(G110), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(KEYINPUT78), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT78), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n554), .A2(new_n561), .A3(new_n558), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n546), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT77), .ZN(new_n565));
  INV_X1    g379(.A(new_n556), .ZN(new_n566));
  INV_X1    g380(.A(new_n557), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(G146), .B1(new_n322), .B2(new_n323), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n568), .B1(new_n376), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n549), .A2(new_n552), .A3(new_n553), .ZN(new_n571));
  AOI21_X1  g385(.A(KEYINPUT76), .B1(new_n571), .B2(G110), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n571), .A2(KEYINPUT76), .A3(G110), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n565), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g389(.A1(new_n325), .A2(new_n326), .B1(new_n566), .B2(new_n567), .ZN(new_n576));
  AOI21_X1  g390(.A(KEYINPUT75), .B1(new_n239), .B2(G119), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n553), .B1(new_n577), .B2(new_n551), .ZN(new_n578));
  INV_X1    g392(.A(new_n552), .ZN(new_n579));
  OAI21_X1  g393(.A(G110), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT76), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n576), .A2(new_n565), .A3(new_n574), .A4(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n564), .B1(new_n575), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n257), .A2(G221), .A3(G234), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(KEYINPUT22), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(G137), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n582), .A2(new_n327), .A3(new_n574), .A4(new_n568), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT77), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n583), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n593), .A2(new_n564), .A3(new_n588), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n590), .A2(KEYINPUT25), .A3(new_n191), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(KEYINPUT80), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n588), .B1(new_n593), .B2(new_n564), .ZN(new_n597));
  AOI211_X1 g411(.A(new_n589), .B(new_n563), .C1(new_n592), .C2(new_n583), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT25), .B1(new_n599), .B2(new_n191), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n590), .A2(new_n191), .A3(new_n594), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT80), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT25), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n307), .B1(G234), .B2(new_n191), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n545), .B1(new_n601), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n602), .A2(new_n604), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n609), .A2(KEYINPUT80), .A3(new_n595), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n610), .A2(KEYINPUT81), .A3(new_n606), .A4(new_n605), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n606), .A2(G902), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n599), .A2(new_n612), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n608), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n460), .A2(new_n544), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G101), .ZN(G3));
  NAND2_X1  g430(.A1(new_n517), .A2(new_n191), .ZN(new_n617));
  AOI22_X1  g431(.A1(new_n617), .A2(G472), .B1(new_n517), .B2(new_n518), .ZN(new_n618));
  AND3_X1   g432(.A1(new_n614), .A2(new_n618), .A3(new_n459), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n374), .B1(new_n384), .B2(new_n385), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n305), .A2(KEYINPUT96), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n308), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n305), .A2(KEYINPUT96), .A3(new_n309), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n622), .A2(KEYINPUT33), .A3(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n314), .A2(G902), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT95), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT33), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n626), .B1(new_n312), .B2(new_n627), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n298), .A2(new_n308), .A3(new_n304), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n308), .B1(new_n298), .B2(new_n304), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n626), .B(new_n627), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n624), .B(new_n625), .C1(new_n628), .C2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n312), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n314), .B1(new_n634), .B2(G902), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n620), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n637), .A2(new_n286), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n619), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT34), .B(G104), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  NAND2_X1  g455(.A1(new_n380), .A2(new_n383), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(KEYINPUT20), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n380), .A2(new_n381), .A3(new_n383), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n316), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n645), .A2(new_n646), .A3(new_n374), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n647), .A2(new_n286), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n619), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(new_n649), .B(KEYINPUT97), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT35), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G107), .ZN(G9));
  AOI21_X1  g466(.A(new_n563), .B1(new_n592), .B2(new_n583), .ZN(new_n653));
  OR2_X1    g467(.A1(new_n589), .A2(KEYINPUT36), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n612), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT98), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n608), .A2(new_n611), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n460), .A2(new_n618), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT37), .B(G110), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G12));
  INV_X1    g475(.A(new_n276), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n517), .A2(KEYINPUT32), .A3(new_n518), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n663), .A2(new_n519), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n662), .B1(new_n664), .B2(new_n542), .ZN(new_n665));
  INV_X1    g479(.A(G900), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n282), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n280), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n620), .A2(new_n316), .A3(new_n669), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n658), .A2(new_n459), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n665), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(KEYINPUT99), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(new_n239), .ZN(G30));
  INV_X1    g488(.A(KEYINPUT40), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n668), .B(KEYINPUT39), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n675), .B1(new_n459), .B2(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n457), .B1(new_n444), .B2(new_n451), .ZN(new_n678));
  INV_X1    g492(.A(new_n676), .ZN(new_n679));
  NOR4_X1   g493(.A1(new_n678), .A2(KEYINPUT40), .A3(new_n389), .A4(new_n679), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n269), .A2(new_n275), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT38), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n677), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n506), .A2(new_n513), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n524), .A2(new_n526), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n684), .B1(new_n472), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g500(.A(G472), .B1(new_n686), .B2(G902), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n520), .A2(new_n543), .A3(new_n687), .ZN(new_n688));
  AND3_X1   g502(.A1(new_n608), .A2(new_n611), .A3(new_n657), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n620), .A2(new_n646), .A3(new_n187), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(KEYINPUT100), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT100), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n658), .A2(new_n693), .A3(new_n690), .ZN(new_n694));
  OAI211_X1 g508(.A(new_n683), .B(new_n688), .C1(new_n692), .C2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G143), .ZN(G45));
  AND3_X1   g510(.A1(new_n620), .A2(new_n636), .A3(new_n668), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n658), .A2(new_n697), .A3(new_n459), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n665), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G146), .ZN(G48));
  AOI21_X1  g514(.A(G902), .B1(new_n447), .B2(new_n448), .ZN(new_n701));
  OAI21_X1  g515(.A(KEYINPUT101), .B1(new_n701), .B2(new_n390), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n191), .B1(new_n426), .B2(new_n442), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT101), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n703), .A2(new_n704), .A3(G469), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n706), .A2(new_n452), .A3(new_n388), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(KEYINPUT102), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n708), .A2(new_n544), .A3(new_n614), .A4(new_n638), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT41), .B(G113), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G15));
  NAND4_X1  g525(.A1(new_n708), .A2(new_n544), .A3(new_n614), .A4(new_n648), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G116), .ZN(G18));
  INV_X1    g527(.A(new_n707), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n544), .A2(new_n387), .A3(new_n658), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G119), .ZN(G21));
  AND3_X1   g530(.A1(new_n527), .A2(new_n488), .A3(new_n490), .ZN(new_n717));
  OAI211_X1 g531(.A(new_n514), .B(new_n516), .C1(new_n717), .C2(new_n536), .ZN(new_n718));
  AOI22_X1  g532(.A1(new_n617), .A2(G472), .B1(new_n518), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n620), .A2(new_n646), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n720), .A2(new_n284), .A3(new_n662), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n708), .A2(new_n614), .A3(new_n719), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G122), .ZN(G24));
  INV_X1    g537(.A(KEYINPUT103), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n617), .A2(G472), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n718), .A2(new_n518), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n658), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  AND4_X1   g541(.A1(new_n452), .A2(new_n706), .A3(new_n388), .A4(new_n276), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n697), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n724), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n620), .A2(new_n636), .A3(new_n668), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n731), .A2(new_n707), .A3(new_n662), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n732), .A2(KEYINPUT103), .A3(new_n658), .A4(new_n719), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G125), .ZN(G27));
  AND2_X1   g549(.A1(new_n544), .A2(new_n614), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n390), .A2(new_n191), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n737), .B1(new_n444), .B2(new_n451), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT105), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT104), .B1(new_n454), .B2(new_n455), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n455), .A2(KEYINPUT104), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n739), .B1(new_n742), .B2(G469), .ZN(new_n743));
  NOR4_X1   g557(.A1(new_n740), .A2(new_n741), .A3(KEYINPUT105), .A4(new_n390), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n738), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n681), .A2(new_n187), .ZN(new_n746));
  INV_X1    g560(.A(new_n388), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AND3_X1   g562(.A1(new_n697), .A2(new_n745), .A3(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n736), .A2(KEYINPUT42), .A3(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(new_n544), .A3(new_n614), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT42), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G131), .ZN(G33));
  AND3_X1   g569(.A1(new_n670), .A2(new_n748), .A3(new_n745), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(new_n544), .A3(new_n614), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G134), .ZN(G36));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n374), .B(new_n636), .C1(new_n384), .C2(new_n385), .ZN(new_n760));
  XNOR2_X1  g574(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT106), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(KEYINPUT43), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n645), .A2(new_n374), .A3(new_n636), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n658), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n759), .B1(new_n769), .B2(new_n618), .ZN(new_n770));
  INV_X1    g584(.A(new_n737), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT45), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n740), .A2(new_n741), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n456), .A2(new_n772), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(G469), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n771), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT46), .ZN(new_n777));
  AOI22_X1  g591(.A1(new_n776), .A2(new_n777), .B1(new_n451), .B2(new_n444), .ZN(new_n778));
  OAI211_X1 g592(.A(KEYINPUT46), .B(new_n771), .C1(new_n773), .C2(new_n775), .ZN(new_n779));
  AOI211_X1 g593(.A(new_n747), .B(new_n679), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n746), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n517), .A2(new_n518), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n725), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n783), .A2(KEYINPUT44), .A3(new_n658), .A4(new_n768), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n770), .A2(new_n780), .A3(new_n781), .A4(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G137), .ZN(G39));
  NOR4_X1   g600(.A1(new_n544), .A2(new_n614), .A3(new_n731), .A4(new_n746), .ZN(new_n787));
  INV_X1    g601(.A(new_n778), .ZN(new_n788));
  INV_X1    g602(.A(new_n779), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n388), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(KEYINPUT47), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT47), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n792), .B(new_n388), .C1(new_n788), .C2(new_n789), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n787), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G140), .ZN(G42));
  INV_X1    g609(.A(new_n389), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n682), .A2(new_n796), .A3(new_n187), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(new_n760), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n706), .A2(new_n452), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(KEYINPUT49), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n799), .A2(KEYINPUT49), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n798), .A2(new_n614), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n802), .A2(new_n688), .ZN(new_n803));
  XOR2_X1   g617(.A(new_n803), .B(KEYINPUT107), .Z(new_n804));
  OAI21_X1  g618(.A(new_n665), .B1(new_n671), .B2(new_n698), .ZN(new_n805));
  INV_X1    g619(.A(new_n745), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n669), .A2(new_n747), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n620), .A2(new_n646), .A3(new_n276), .A4(new_n807), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n806), .A2(new_n658), .A3(new_n808), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n809), .A2(KEYINPUT109), .A3(new_n688), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT109), .B1(new_n809), .B2(new_n688), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n734), .B(new_n805), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n809), .A2(new_n688), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT109), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n809), .A2(KEYINPUT109), .A3(new_n688), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n819), .A2(KEYINPUT52), .A3(new_n734), .A4(new_n805), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n814), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n286), .B1(new_n637), .B2(new_n647), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n822), .A2(new_n614), .A3(new_n618), .A4(new_n459), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n615), .A2(new_n659), .A3(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n727), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n749), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n826), .A2(new_n757), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT111), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n658), .A2(new_n459), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n386), .A2(KEYINPUT108), .A3(new_n669), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(new_n746), .ZN(new_n831));
  OAI21_X1  g645(.A(KEYINPUT108), .B1(new_n386), .B2(new_n669), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n829), .A2(new_n544), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n824), .A2(new_n827), .A3(new_n828), .A4(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n833), .A2(new_n826), .A3(new_n757), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n615), .A2(new_n659), .A3(new_n823), .ZN(new_n836));
  OAI21_X1  g650(.A(KEYINPUT111), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AND4_X1   g651(.A1(new_n709), .A2(new_n712), .A3(new_n722), .A4(new_n715), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n834), .A2(new_n837), .A3(new_n754), .A4(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT53), .B1(new_n821), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT52), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n812), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(new_n820), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n835), .A2(new_n836), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n844), .A2(new_n754), .A3(new_n838), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n843), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(KEYINPUT54), .B1(new_n840), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n846), .B1(new_n843), .B2(new_n845), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n844), .A2(new_n838), .A3(new_n846), .A4(new_n754), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n850), .B1(new_n820), .B2(new_n814), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n849), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n791), .A2(new_n793), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n854), .B1(new_n796), .B2(new_n799), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n614), .A2(new_n719), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n280), .B1(new_n763), .B2(new_n767), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n855), .A2(new_n781), .A3(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT50), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n187), .B1(KEYINPUT112), .B2(new_n860), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n682), .A2(new_n714), .A3(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n856), .A2(new_n857), .A3(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n860), .A2(KEYINPUT112), .ZN(new_n864));
  XOR2_X1   g678(.A(new_n863), .B(new_n864), .Z(new_n865));
  NOR3_X1   g679(.A1(new_n707), .A2(new_n280), .A3(new_n746), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(new_n614), .ZN(new_n867));
  NOR4_X1   g681(.A1(new_n867), .A2(new_n688), .A3(new_n620), .A4(new_n636), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n866), .A2(new_n768), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n825), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT113), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n869), .A2(KEYINPUT113), .A3(new_n825), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n868), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n859), .A2(new_n865), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT51), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n859), .A2(KEYINPUT51), .A3(new_n865), .A4(new_n874), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n736), .A2(new_n869), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n879), .B(KEYINPUT48), .Z(new_n880));
  NOR3_X1   g694(.A1(new_n867), .A2(new_n688), .A3(new_n637), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n858), .A2(new_n728), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n277), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n880), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n877), .A2(new_n878), .A3(new_n884), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n848), .A2(new_n853), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(G952), .A2(G953), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n804), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT114), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT114), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n890), .B(new_n804), .C1(new_n886), .C2(new_n887), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n889), .A2(new_n891), .ZN(G75));
  NAND2_X1  g706(.A1(new_n840), .A2(new_n847), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n893), .A2(new_n191), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(G210), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT56), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n264), .A2(new_n267), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(new_n265), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT55), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n895), .A2(new_n896), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n899), .B1(new_n895), .B2(new_n896), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n257), .A2(G952), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(G51));
  XNOR2_X1  g717(.A(new_n737), .B(KEYINPUT57), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n840), .A2(KEYINPUT54), .A3(new_n847), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n904), .B1(new_n906), .B2(new_n848), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n449), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n773), .A2(new_n775), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n894), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n902), .B1(new_n908), .B2(new_n910), .ZN(G54));
  AND2_X1   g725(.A1(KEYINPUT58), .A2(G475), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n840), .A2(G902), .A3(new_n847), .A4(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n380), .ZN(new_n914));
  OR2_X1    g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(new_n902), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n913), .A2(new_n914), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(KEYINPUT115), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT115), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n915), .A2(new_n920), .A3(new_n916), .A4(new_n917), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n919), .A2(new_n921), .ZN(G60));
  OAI21_X1  g736(.A(new_n624), .B1(new_n628), .B2(new_n632), .ZN(new_n923));
  NAND2_X1  g737(.A1(G478), .A2(G902), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT59), .Z(new_n925));
  NOR2_X1   g739(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n893), .A2(new_n852), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n927), .B1(new_n928), .B2(new_n905), .ZN(new_n929));
  OAI21_X1  g743(.A(KEYINPUT116), .B1(new_n929), .B2(new_n902), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n926), .B1(new_n906), .B2(new_n848), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT116), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n931), .A2(new_n932), .A3(new_n916), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n848), .A2(new_n853), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n923), .B1(new_n934), .B2(new_n925), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n930), .A2(new_n933), .A3(new_n935), .ZN(G63));
  NAND2_X1  g750(.A1(G217), .A2(G902), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT60), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n840), .A2(new_n847), .A3(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n599), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n902), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n840), .A2(new_n655), .A3(new_n847), .A4(new_n939), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(KEYINPUT117), .A2(KEYINPUT61), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT117), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT61), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n944), .A2(new_n945), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n948), .B1(new_n944), .B2(new_n945), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n949), .A2(new_n950), .ZN(G66));
  INV_X1    g765(.A(G224), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n283), .A2(new_n952), .A3(new_n257), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n709), .A2(new_n712), .A3(new_n722), .A4(new_n715), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n954), .A2(new_n836), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n953), .B1(new_n955), .B2(new_n257), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n897), .B1(G898), .B2(new_n257), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(G69));
  OAI21_X1  g772(.A(new_n501), .B1(new_n511), .B2(KEYINPUT30), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(new_n377), .Z(new_n960));
  XNOR2_X1  g774(.A(KEYINPUT118), .B(KEYINPUT119), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n392), .A2(G900), .A3(G953), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT121), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n754), .A2(new_n965), .A3(new_n757), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n965), .B1(new_n754), .B2(new_n757), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n734), .A2(new_n805), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n720), .A2(new_n662), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n736), .A2(new_n970), .A3(new_n780), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n794), .A2(new_n785), .A3(new_n971), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n968), .A2(new_n969), .A3(new_n972), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n963), .B(new_n964), .C1(new_n973), .C2(G953), .ZN(new_n974));
  NAND3_X1  g788(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT62), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n695), .A2(new_n734), .A3(new_n805), .A4(new_n976), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n977), .A2(new_n794), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n695), .A2(new_n734), .A3(new_n805), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n979), .A2(KEYINPUT120), .A3(KEYINPUT62), .ZN(new_n980));
  AOI21_X1  g794(.A(KEYINPUT120), .B1(new_n979), .B2(KEYINPUT62), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n978), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n678), .A2(new_n389), .A3(new_n679), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n746), .B1(new_n637), .B2(new_n647), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n736), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n785), .A2(new_n985), .A3(new_n257), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n975), .B(new_n962), .C1(new_n982), .C2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n974), .A2(new_n987), .ZN(G72));
  INV_X1    g802(.A(KEYINPUT125), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n785), .A2(new_n985), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n990), .A2(new_n954), .A3(new_n836), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n978), .B(new_n991), .C1(new_n980), .C2(new_n981), .ZN(new_n992));
  XNOR2_X1  g806(.A(KEYINPUT122), .B(KEYINPUT63), .ZN(new_n993));
  NAND2_X1  g807(.A1(G472), .A2(G902), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n993), .B(new_n994), .Z(new_n995));
  NAND3_X1  g809(.A1(new_n992), .A2(KEYINPUT123), .A3(new_n995), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n538), .B(KEYINPUT124), .ZN(new_n997));
  AND2_X1   g811(.A1(new_n997), .A2(new_n536), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(KEYINPUT123), .B1(new_n992), .B2(new_n995), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n989), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n992), .A2(new_n995), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT123), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n1004), .A2(KEYINPUT125), .A3(new_n996), .A4(new_n998), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1001), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n972), .A2(new_n969), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n1007), .B(new_n955), .C1(new_n966), .C2(new_n967), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1008), .A2(new_n995), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n997), .A2(new_n536), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n849), .A2(new_n851), .ZN(new_n1011));
  INV_X1    g825(.A(new_n995), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT126), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n684), .B1(new_n1013), .B2(new_n539), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n538), .A2(KEYINPUT126), .A3(new_n472), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1012), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  AOI221_X4 g830(.A(new_n902), .B1(new_n1009), .B2(new_n1010), .C1(new_n1011), .C2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1006), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT127), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n1006), .A2(new_n1017), .A3(KEYINPUT127), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1020), .A2(new_n1021), .ZN(G57));
endmodule


