//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 0 1 1 0 0 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n781, new_n783, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n990, new_n991;
  INV_X1    g000(.A(G71gat), .ZN(new_n202));
  INV_X1    g001(.A(G78gat), .ZN(new_n203));
  OAI211_X1 g002(.A(new_n202), .B(new_n203), .C1(KEYINPUT97), .C2(KEYINPUT9), .ZN(new_n204));
  NAND2_X1  g003(.A1(G71gat), .A2(G78gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT9), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AOI22_X1  g006(.A1(new_n204), .A2(new_n205), .B1(new_n207), .B2(KEYINPUT97), .ZN(new_n208));
  AND2_X1   g007(.A1(G57gat), .A2(G64gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(G57gat), .A2(G64gat), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT96), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  OR2_X1    g010(.A1(G57gat), .A2(G64gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT96), .ZN(new_n213));
  NAND2_X1  g012(.A1(G57gat), .A2(G64gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n208), .A2(new_n211), .A3(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n209), .A2(new_n210), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT9), .ZN(new_n218));
  OR3_X1    g017(.A1(KEYINPUT95), .A2(G71gat), .A3(G78gat), .ZN(new_n219));
  OAI21_X1  g018(.A(KEYINPUT95), .B1(G71gat), .B2(G78gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n218), .A2(new_n221), .A3(new_n205), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n216), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT21), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G231gat), .A2(G233gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n225), .B(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G127gat), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G15gat), .B(G22gat), .ZN(new_n230));
  OR2_X1    g029(.A1(new_n230), .A2(G1gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT93), .ZN(new_n232));
  AOI21_X1  g031(.A(G8gat), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT16), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n230), .B1(new_n234), .B2(G1gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n231), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n233), .B(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n237), .B1(new_n224), .B2(new_n223), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n238), .B(KEYINPUT98), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n229), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(G155gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(G183gat), .B(G211gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n240), .B(new_n244), .ZN(new_n245));
  AND2_X1   g044(.A1(G43gat), .A2(G50gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(G43gat), .A2(G50gat), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT15), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(new_n248), .B(KEYINPUT90), .Z(new_n249));
  OAI21_X1  g048(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(KEYINPUT88), .ZN(new_n251));
  OR3_X1    g050(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n252));
  AOI22_X1  g051(.A1(new_n251), .A2(new_n252), .B1(G29gat), .B2(G36gat), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT15), .ZN(new_n254));
  XOR2_X1   g053(.A(KEYINPUT92), .B(G50gat), .Z(new_n255));
  NOR2_X1   g054(.A1(new_n255), .A2(G43gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT91), .B(G43gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n257), .A2(G50gat), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n254), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n249), .A2(new_n253), .A3(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n248), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(new_n252), .ZN(new_n263));
  OR2_X1    g062(.A1(new_n251), .A2(KEYINPUT89), .ZN(new_n264));
  AOI22_X1  g063(.A1(new_n251), .A2(KEYINPUT89), .B1(G29gat), .B2(G36gat), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT100), .ZN(new_n269));
  NAND2_X1  g068(.A1(G99gat), .A2(G106gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT8), .ZN(new_n271));
  NAND2_X1  g070(.A1(G85gat), .A2(G92gat), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT7), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G85gat), .ZN(new_n275));
  INV_X1    g074(.A(G92gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n271), .A2(new_n274), .A3(new_n277), .A4(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G99gat), .B(G106gat), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  AND3_X1   g081(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI22_X1  g084(.A1(KEYINPUT8), .A2(new_n270), .B1(new_n275), .B2(new_n276), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n280), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n269), .B1(new_n282), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n285), .A2(new_n280), .A3(new_n286), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT100), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  AND2_X1   g091(.A1(G232gat), .A2(G233gat), .ZN(new_n293));
  AOI22_X1  g092(.A1(new_n268), .A2(new_n292), .B1(KEYINPUT41), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT17), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n295), .B1(new_n261), .B2(new_n266), .ZN(new_n296));
  INV_X1    g095(.A(new_n266), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n297), .A2(KEYINPUT17), .A3(new_n260), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n296), .A2(new_n298), .A3(new_n291), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  XOR2_X1   g099(.A(G190gat), .B(G218gat), .Z(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n293), .A2(KEYINPUT41), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n303), .B(KEYINPUT99), .ZN(new_n304));
  XNOR2_X1  g103(.A(G134gat), .B(G162gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n304), .B(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n301), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n294), .A2(new_n307), .A3(new_n299), .ZN(new_n308));
  AND3_X1   g107(.A1(new_n302), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n306), .B1(new_n302), .B2(new_n308), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n245), .A2(new_n311), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n215), .A2(new_n211), .ZN(new_n313));
  AOI22_X1  g112(.A1(new_n217), .A2(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n313), .A2(new_n208), .B1(new_n314), .B2(new_n221), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT10), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT102), .B1(new_n316), .B2(new_n291), .ZN(new_n317));
  AND3_X1   g116(.A1(new_n216), .A2(KEYINPUT10), .A3(new_n222), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT102), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n318), .A2(new_n319), .A3(new_n288), .A4(new_n290), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n279), .A2(new_n281), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n216), .A2(new_n222), .A3(new_n289), .A4(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT101), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n282), .A2(new_n287), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT101), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n315), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT10), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n291), .A2(new_n223), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n321), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(G230gat), .A2(G233gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n324), .A2(new_n327), .B1(new_n291), .B2(new_n223), .ZN(new_n335));
  OR2_X1    g134(.A1(new_n335), .A2(new_n333), .ZN(new_n336));
  AND2_X1   g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G120gat), .B(G148gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(G176gat), .B(G204gat), .ZN(new_n339));
  XOR2_X1   g138(.A(new_n338), .B(new_n339), .Z(new_n340));
  OR2_X1    g139(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n335), .A2(new_n329), .B1(new_n317), .B2(new_n320), .ZN(new_n342));
  INV_X1    g141(.A(new_n333), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n336), .B(new_n340), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT103), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n334), .A2(KEYINPUT103), .A3(new_n336), .A4(new_n340), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n341), .A2(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n312), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(KEYINPUT71), .A2(KEYINPUT36), .ZN(new_n352));
  INV_X1    g151(.A(G183gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT27), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT27), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(G183gat), .ZN(new_n356));
  INV_X1    g155(.A(G190gat), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n354), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT28), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n358), .B(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(G183gat), .A2(G190gat), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NOR2_X1   g161(.A1(G169gat), .A2(G176gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n363), .B(KEYINPUT26), .ZN(new_n364));
  NAND2_X1  g163(.A1(G169gat), .A2(G176gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT65), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT65), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n367), .A2(G169gat), .A3(G176gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n362), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n360), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n361), .A2(KEYINPUT24), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT24), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n373), .A2(G183gat), .A3(G190gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n353), .A2(new_n357), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT25), .B1(new_n363), .B2(KEYINPUT23), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  AOI221_X4 g179(.A(KEYINPUT66), .B1(new_n363), .B2(KEYINPUT23), .C1(new_n366), .C2(new_n368), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT66), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n363), .A2(KEYINPUT23), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n382), .B1(new_n369), .B2(new_n383), .ZN(new_n384));
  NOR3_X1   g183(.A1(new_n380), .A2(new_n381), .A3(new_n384), .ZN(new_n385));
  OR2_X1    g184(.A1(G169gat), .A2(G176gat), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT23), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n369), .A2(new_n383), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT64), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n392), .A2(new_n353), .A3(new_n357), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n375), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT25), .B1(new_n390), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n371), .B1(new_n385), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT69), .ZN(new_n397));
  OR2_X1    g196(.A1(new_n228), .A2(G134gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n228), .A2(G134gat), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT1), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT67), .ZN(new_n402));
  INV_X1    g201(.A(G120gat), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n402), .B1(new_n403), .B2(G113gat), .ZN(new_n404));
  INV_X1    g203(.A(G113gat), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n405), .A2(KEYINPUT67), .A3(G120gat), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n404), .B(new_n406), .C1(new_n405), .C2(G120gat), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n405), .A2(G120gat), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n403), .A2(G113gat), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n400), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n398), .A2(new_n399), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n401), .A2(new_n407), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n396), .A2(new_n397), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n369), .A2(new_n383), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT66), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n378), .B1(new_n375), .B2(new_n376), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n369), .A2(new_n382), .A3(new_n383), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT25), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n353), .A2(KEYINPUT24), .ZN(new_n421));
  AOI22_X1  g220(.A1(new_n421), .A2(G190gat), .B1(KEYINPUT24), .B2(new_n361), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n393), .A2(new_n391), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n420), .B1(new_n424), .B2(new_n389), .ZN(new_n425));
  AOI22_X1  g224(.A1(new_n419), .A2(new_n425), .B1(new_n360), .B2(new_n370), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT69), .B1(new_n426), .B2(new_n412), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n414), .A2(new_n427), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n412), .B(new_n371), .C1(new_n385), .C2(new_n395), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT68), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT68), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n426), .A2(new_n431), .A3(new_n412), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n428), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(G227gat), .A2(G233gat), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT34), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  AOI22_X1  g236(.A1(new_n427), .A2(new_n414), .B1(new_n430), .B2(new_n432), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT34), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n438), .A2(new_n439), .A3(new_n435), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT33), .B1(new_n434), .B2(new_n436), .ZN(new_n441));
  XNOR2_X1  g240(.A(G15gat), .B(G43gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n442), .B(KEYINPUT70), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n443), .B(new_n202), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n444), .B(G99gat), .Z(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n437), .B(new_n440), .C1(new_n441), .C2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT33), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n448), .B1(new_n438), .B2(new_n435), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n439), .B1(new_n438), .B2(new_n435), .ZN(new_n450));
  AND4_X1   g249(.A1(new_n439), .A2(new_n428), .A3(new_n433), .A4(new_n435), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n449), .B(new_n445), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n434), .A2(new_n436), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT32), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n447), .A2(new_n452), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n455), .B1(new_n447), .B2(new_n452), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n352), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n447), .A2(new_n452), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n454), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n447), .A2(new_n452), .A3(new_n455), .ZN(new_n461));
  XNOR2_X1  g260(.A(KEYINPUT71), .B(KEYINPUT36), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(G78gat), .B(G106gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n465), .B(KEYINPUT82), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n466), .B(G50gat), .ZN(new_n467));
  XOR2_X1   g266(.A(KEYINPUT81), .B(KEYINPUT31), .Z(new_n468));
  XNOR2_X1  g267(.A(new_n467), .B(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n469), .B(KEYINPUT84), .ZN(new_n470));
  XOR2_X1   g269(.A(G141gat), .B(G148gat), .Z(new_n471));
  XNOR2_X1  g270(.A(G155gat), .B(G162gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(G155gat), .A2(G162gat), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT76), .B1(new_n473), .B2(KEYINPUT2), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n471), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n472), .B1(new_n471), .B2(new_n474), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G211gat), .B(G218gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n478), .B(KEYINPUT72), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n480));
  INV_X1    g279(.A(G197gat), .ZN(new_n481));
  INV_X1    g280(.A(G204gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(G197gat), .A2(G204gat), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n480), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n479), .B(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT29), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT3), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n477), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n471), .A2(new_n474), .ZN(new_n491));
  INV_X1    g290(.A(new_n472), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n471), .A2(new_n472), .A3(new_n474), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(new_n489), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n486), .B1(new_n487), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT83), .B1(new_n490), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(G22gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(G228gat), .ZN(new_n500));
  INV_X1    g299(.A(G233gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  OAI211_X1 g302(.A(KEYINPUT83), .B(G22gat), .C1(new_n490), .C2(new_n496), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n499), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n503), .B1(new_n499), .B2(new_n504), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n470), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n499), .A2(new_n504), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n502), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT84), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n469), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(new_n512), .A3(new_n505), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n508), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(G226gat), .A2(G233gat), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT73), .ZN(new_n517));
  AOI221_X4 g316(.A(new_n517), .B1(new_n360), .B2(new_n370), .C1(new_n419), .C2(new_n425), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n419), .A2(new_n425), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT73), .B1(new_n519), .B2(new_n371), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n516), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT74), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT74), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n523), .B(new_n516), .C1(new_n518), .C2(new_n520), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n516), .B1(new_n396), .B2(new_n487), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n522), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n486), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n516), .A2(KEYINPUT29), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n530), .B1(new_n518), .B2(new_n520), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n426), .A2(new_n516), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n528), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(G8gat), .B(G36gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(G64gat), .B(G92gat), .ZN(new_n536));
  XOR2_X1   g335(.A(new_n535), .B(new_n536), .Z(new_n537));
  NAND4_X1  g336(.A1(new_n529), .A2(new_n534), .A3(KEYINPUT30), .A4(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n537), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n525), .B1(new_n521), .B2(KEYINPUT74), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n486), .B1(new_n540), .B2(new_n524), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n539), .B1(new_n541), .B2(new_n533), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  AOI211_X1 g342(.A(new_n533), .B(new_n539), .C1(new_n527), .C2(new_n528), .ZN(new_n544));
  OAI21_X1  g343(.A(KEYINPUT75), .B1(new_n544), .B2(KEYINPUT30), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n529), .A2(new_n534), .A3(new_n537), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT75), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT30), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n543), .B1(new_n545), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(KEYINPUT3), .B1(new_n475), .B2(new_n476), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n413), .A2(new_n551), .A3(new_n495), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n401), .A2(new_n407), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n410), .A2(new_n411), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n553), .A2(new_n493), .A3(new_n494), .A4(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT4), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G225gat), .A2(G233gat), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n477), .A2(KEYINPUT4), .A3(new_n412), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n552), .A2(new_n557), .A3(new_n558), .A4(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT79), .ZN(new_n561));
  XOR2_X1   g360(.A(KEYINPUT78), .B(KEYINPUT5), .Z(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  OR3_X1    g362(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n561), .B1(new_n560), .B2(new_n563), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT77), .B1(new_n477), .B2(new_n412), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n566), .B1(new_n477), .B2(new_n412), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n413), .B(KEYINPUT77), .C1(new_n476), .C2(new_n475), .ZN(new_n568));
  INV_X1    g367(.A(new_n558), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n560), .A2(new_n563), .ZN(new_n571));
  AOI22_X1  g370(.A1(new_n564), .A2(new_n565), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G1gat), .B(G29gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT0), .ZN(new_n574));
  XNOR2_X1  g373(.A(G57gat), .B(G85gat), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n574), .B(new_n575), .Z(new_n576));
  OAI21_X1  g375(.A(KEYINPUT80), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(KEYINPUT6), .B1(new_n572), .B2(new_n576), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n571), .A2(new_n570), .ZN(new_n579));
  INV_X1    g378(.A(new_n565), .ZN(new_n580));
  NOR3_X1   g379(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT80), .ZN(new_n583));
  INV_X1    g382(.A(new_n576), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n577), .A2(new_n578), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n582), .A2(KEYINPUT6), .A3(new_n584), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n514), .B1(new_n550), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(KEYINPUT85), .B1(new_n464), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n543), .ZN(new_n591));
  NOR3_X1   g390(.A1(new_n544), .A2(KEYINPUT75), .A3(KEYINPUT30), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n547), .B1(new_n546), .B2(new_n548), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n588), .B(new_n591), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n508), .A2(new_n513), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT85), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n458), .A2(new_n463), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT38), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n528), .B1(new_n540), .B2(new_n524), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n396), .A2(new_n517), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n426), .A2(KEYINPUT73), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI22_X1  g403(.A1(new_n604), .A2(new_n530), .B1(new_n516), .B2(new_n426), .ZN(new_n605));
  OAI21_X1  g404(.A(KEYINPUT37), .B1(new_n605), .B2(new_n486), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n600), .B1(new_n601), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n539), .A2(KEYINPUT37), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n607), .B1(new_n542), .B2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT6), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n610), .B1(new_n582), .B2(new_n584), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n572), .A2(new_n576), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n546), .B(new_n587), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n529), .A2(new_n534), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n615), .A2(KEYINPUT37), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n539), .B1(new_n615), .B2(KEYINPUT37), .ZN(new_n617));
  OAI21_X1  g416(.A(KEYINPUT38), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n595), .B1(new_n614), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT87), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n552), .A2(new_n557), .A3(new_n559), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(new_n569), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n567), .A2(new_n568), .ZN(new_n623));
  OAI211_X1 g422(.A(KEYINPUT39), .B(new_n622), .C1(new_n623), .C2(new_n569), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n622), .A2(KEYINPUT39), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n624), .A2(new_n576), .A3(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT40), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(KEYINPUT86), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT86), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n626), .A2(new_n630), .A3(new_n627), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n612), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n626), .A2(new_n627), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n620), .B1(new_n550), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n634), .A2(new_n633), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n638), .B1(new_n629), .B2(new_n631), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n637), .A2(new_n639), .A3(KEYINPUT87), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n619), .A2(new_n636), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n590), .A2(new_n599), .A3(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n456), .A2(new_n457), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n514), .ZN(new_n644));
  OAI21_X1  g443(.A(KEYINPUT35), .B1(new_n644), .B2(new_n594), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n633), .A2(new_n578), .ZN(new_n646));
  AOI21_X1  g445(.A(KEYINPUT35), .B1(new_n646), .B2(new_n587), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n550), .A2(new_n643), .A3(new_n514), .A4(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n642), .A2(new_n649), .ZN(new_n650));
  OR2_X1    g449(.A1(new_n267), .A2(new_n237), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n296), .A2(new_n298), .A3(new_n237), .ZN(new_n652));
  NAND2_X1  g451(.A1(G229gat), .A2(G233gat), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT18), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n651), .A2(new_n652), .A3(KEYINPUT18), .A4(new_n653), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n267), .B(new_n237), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n653), .B(KEYINPUT13), .Z(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n656), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(G113gat), .B(G141gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G197gat), .ZN(new_n663));
  XOR2_X1   g462(.A(KEYINPUT11), .B(G169gat), .Z(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT12), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n661), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n656), .A2(new_n660), .A3(new_n666), .A4(new_n657), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n650), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT94), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n650), .A2(KEYINPUT94), .A3(new_n670), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n351), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n588), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(G1gat), .ZN(G1324gat));
  INV_X1    g477(.A(KEYINPUT42), .ZN(new_n679));
  AOI21_X1  g478(.A(KEYINPUT94), .B1(new_n650), .B2(new_n670), .ZN(new_n680));
  INV_X1    g479(.A(new_n670), .ZN(new_n681));
  AOI211_X1 g480(.A(new_n672), .B(new_n681), .C1(new_n642), .C2(new_n649), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n637), .B(new_n350), .C1(new_n680), .C2(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(KEYINPUT16), .B(G8gat), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n679), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(KEYINPUT104), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n687), .B(new_n679), .C1(new_n683), .C2(new_n684), .ZN(new_n688));
  OR3_X1    g487(.A1(new_n683), .A2(new_n679), .A3(new_n684), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n683), .A2(G8gat), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n686), .A2(new_n688), .A3(new_n689), .A4(new_n690), .ZN(G1325gat));
  INV_X1    g490(.A(G15gat), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n675), .A2(new_n692), .A3(new_n643), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n598), .A2(KEYINPUT105), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n458), .A2(new_n463), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  OAI211_X1 g497(.A(new_n350), .B(new_n698), .C1(new_n680), .C2(new_n682), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(G15gat), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n693), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT106), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n693), .A2(new_n700), .A3(KEYINPUT106), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(G1326gat));
  NAND2_X1  g504(.A1(new_n675), .A2(new_n595), .ZN(new_n706));
  XNOR2_X1  g505(.A(KEYINPUT43), .B(G22gat), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1327gat));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n311), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n650), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n464), .A2(new_n589), .ZN(new_n713));
  AOI22_X1  g512(.A1(new_n641), .A2(new_n713), .B1(new_n645), .B2(new_n648), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n710), .B1(new_n714), .B2(new_n311), .ZN(new_n715));
  INV_X1    g514(.A(new_n245), .ZN(new_n716));
  INV_X1    g515(.A(new_n349), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n718), .A2(new_n681), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n712), .A2(new_n715), .A3(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n709), .B1(new_n721), .B2(new_n588), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n720), .A2(KEYINPUT107), .A3(new_n676), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n722), .A2(G29gat), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n673), .A2(new_n674), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n718), .A2(new_n311), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT45), .ZN(new_n728));
  OR2_X1    g527(.A1(new_n588), .A2(G29gat), .ZN(new_n729));
  OR3_X1    g528(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n728), .B1(new_n727), .B2(new_n729), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n724), .A2(new_n730), .A3(new_n731), .ZN(G1328gat));
  NOR2_X1   g531(.A1(new_n550), .A2(G36gat), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n725), .A2(new_n726), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(KEYINPUT46), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT108), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n734), .A2(new_n737), .A3(KEYINPUT46), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT46), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n725), .A2(new_n739), .A3(new_n726), .A4(new_n733), .ZN(new_n740));
  OAI21_X1  g539(.A(G36gat), .B1(new_n721), .B2(new_n550), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n736), .A2(new_n738), .A3(new_n740), .A4(new_n741), .ZN(G1329gat));
  INV_X1    g541(.A(new_n257), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n743), .B1(new_n721), .B2(new_n598), .ZN(new_n744));
  INV_X1    g543(.A(new_n643), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n745), .A2(new_n743), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n726), .B(new_n746), .C1(new_n680), .C2(new_n682), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n744), .A2(KEYINPUT47), .A3(new_n747), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n712), .A2(new_n715), .A3(new_n698), .A4(new_n719), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT109), .ZN(new_n750));
  AND3_X1   g549(.A1(new_n749), .A2(new_n750), .A3(new_n743), .ZN(new_n751));
  INV_X1    g550(.A(new_n747), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n750), .B1(new_n749), .B2(new_n743), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n751), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n748), .B1(new_n754), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n756));
  INV_X1    g555(.A(new_n255), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n514), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n725), .A2(new_n756), .A3(new_n726), .A4(new_n758), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n726), .B(new_n758), .C1(new_n680), .C2(new_n682), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT110), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n712), .A2(new_n715), .A3(new_n595), .A4(new_n719), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n757), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n759), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT48), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n762), .A2(KEYINPUT111), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n757), .B1(new_n762), .B2(KEYINPUT111), .ZN(new_n768));
  OAI211_X1 g567(.A(KEYINPUT48), .B(new_n760), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n766), .A2(new_n769), .ZN(G1331gat));
  NOR4_X1   g569(.A1(new_n714), .A2(new_n670), .A3(new_n312), .A4(new_n717), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n676), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g572(.A(new_n550), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT112), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n777));
  XOR2_X1   g576(.A(new_n776), .B(new_n777), .Z(G1333gat));
  AOI21_X1  g577(.A(new_n202), .B1(new_n771), .B2(new_n698), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n745), .A2(G71gat), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n779), .B1(new_n771), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g581(.A1(new_n771), .A2(new_n595), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(G78gat), .ZN(G1335gat));
  AND2_X1   g583(.A1(new_n712), .A2(new_n715), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n245), .A2(new_n717), .A3(new_n670), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(G85gat), .B1(new_n787), .B2(new_n588), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n714), .A2(new_n311), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n245), .A2(new_n670), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n789), .A2(KEYINPUT51), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT51), .B1(new_n789), .B2(new_n790), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n676), .A2(new_n275), .A3(new_n349), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n788), .B1(new_n793), .B2(new_n794), .ZN(G1336gat));
  NAND3_X1  g594(.A1(new_n785), .A2(new_n637), .A3(new_n786), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(G92gat), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n550), .A2(G92gat), .A3(new_n717), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n799), .B1(new_n791), .B2(new_n792), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n793), .ZN(new_n802));
  XOR2_X1   g601(.A(new_n799), .B(KEYINPUT113), .Z(new_n803));
  AOI22_X1  g602(.A1(new_n802), .A2(new_n803), .B1(new_n796), .B2(G92gat), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n801), .B1(new_n804), .B2(new_n798), .ZN(G1337gat));
  OAI21_X1  g604(.A(KEYINPUT114), .B1(new_n787), .B2(new_n697), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(G99gat), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n787), .A2(KEYINPUT114), .A3(new_n697), .ZN(new_n808));
  OR3_X1    g607(.A1(new_n745), .A2(G99gat), .A3(new_n717), .ZN(new_n809));
  OAI22_X1  g608(.A1(new_n807), .A2(new_n808), .B1(new_n793), .B2(new_n809), .ZN(G1338gat));
  NAND4_X1  g609(.A1(new_n712), .A2(new_n715), .A3(new_n595), .A4(new_n786), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(G106gat), .ZN(new_n812));
  OR3_X1    g611(.A1(new_n514), .A2(new_n717), .A3(G106gat), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n812), .B1(new_n793), .B2(new_n813), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g614(.A(new_n311), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n321), .A2(new_n331), .A3(new_n343), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n334), .A2(KEYINPUT54), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n343), .B1(new_n321), .B2(new_n331), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n340), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT55), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n818), .A2(KEYINPUT55), .A3(new_n821), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n348), .A2(KEYINPUT115), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT115), .B1(new_n348), .B2(new_n824), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n670), .B(new_n823), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n658), .A2(new_n659), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n653), .B1(new_n651), .B2(new_n652), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n665), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n349), .A2(new_n669), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n816), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n825), .A2(new_n826), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n669), .B(new_n830), .C1(new_n309), .C2(new_n310), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n833), .A2(new_n822), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n716), .B1(new_n832), .B2(new_n835), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n312), .A2(new_n670), .A3(new_n349), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n836), .A2(KEYINPUT116), .A3(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(KEYINPUT116), .B1(new_n836), .B2(new_n838), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n550), .A2(new_n676), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n842), .A2(new_n514), .A3(new_n643), .A4(new_n844), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n845), .A2(new_n405), .A3(new_n681), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n836), .A2(new_n838), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT116), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n644), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n849), .A2(new_n676), .A3(new_n850), .A4(new_n839), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n852));
  OR2_X1    g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n852), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n853), .A2(new_n550), .A3(new_n854), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n855), .A2(new_n681), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n846), .B1(new_n856), .B2(new_n405), .ZN(G1340gat));
  NAND2_X1  g656(.A1(new_n349), .A2(new_n403), .ZN(new_n858));
  XOR2_X1   g657(.A(new_n858), .B(KEYINPUT118), .Z(new_n859));
  NAND4_X1  g658(.A1(new_n853), .A2(new_n550), .A3(new_n854), .A4(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(G120gat), .B1(new_n845), .B2(new_n717), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n860), .A2(new_n861), .A3(KEYINPUT119), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(G1341gat));
  OAI21_X1  g665(.A(G127gat), .B1(new_n845), .B2(new_n716), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n245), .A2(new_n228), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n867), .B1(new_n855), .B2(new_n868), .ZN(G1342gat));
  NOR2_X1   g668(.A1(new_n311), .A2(G134gat), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n853), .A2(new_n550), .A3(new_n854), .A4(new_n870), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n871), .A2(KEYINPUT56), .ZN(new_n872));
  OAI21_X1  g671(.A(G134gat), .B1(new_n845), .B2(new_n311), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(KEYINPUT56), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(G1343gat));
  INV_X1    g674(.A(KEYINPUT121), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n849), .A2(new_n877), .A3(new_n595), .A4(new_n839), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n844), .A2(new_n598), .ZN(new_n879));
  OR3_X1    g678(.A1(new_n833), .A2(new_n822), .A3(new_n834), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n823), .A2(new_n348), .A3(new_n824), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n831), .B1(new_n681), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n311), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n245), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n595), .B1(new_n884), .B2(new_n837), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n879), .B1(new_n885), .B2(KEYINPUT57), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n878), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n876), .B1(new_n887), .B2(new_n681), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n878), .A2(new_n886), .A3(KEYINPUT121), .A4(new_n670), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n888), .A2(G141gat), .A3(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT58), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT120), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n842), .A2(new_n892), .A3(new_n676), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n849), .A2(new_n839), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT120), .B1(new_n894), .B2(new_n588), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n698), .A2(new_n637), .A3(new_n514), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n893), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n681), .A2(G141gat), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n890), .B(new_n891), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(G141gat), .B1(new_n887), .B2(new_n681), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n900), .B1(new_n897), .B2(new_n898), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(KEYINPUT58), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n899), .A2(new_n902), .ZN(G1344gat));
  INV_X1    g702(.A(new_n897), .ZN(new_n904));
  INV_X1    g703(.A(G148gat), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n904), .A2(new_n905), .A3(new_n349), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n907));
  INV_X1    g706(.A(new_n879), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n514), .A2(new_n877), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n840), .A2(new_n841), .A3(new_n910), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n885), .A2(new_n877), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n349), .B(new_n908), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n905), .B1(new_n913), .B2(KEYINPUT122), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n849), .A2(new_n839), .A3(new_n909), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n885), .A2(new_n877), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n917), .A2(new_n918), .A3(new_n349), .A4(new_n908), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n907), .B1(new_n914), .B2(new_n919), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n887), .A2(new_n717), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n921), .A2(KEYINPUT59), .A3(new_n905), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n906), .B1(new_n920), .B2(new_n922), .ZN(G1345gat));
  OAI21_X1  g722(.A(G155gat), .B1(new_n887), .B2(new_n716), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n716), .A2(G155gat), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n924), .B1(new_n897), .B2(new_n925), .ZN(G1346gat));
  INV_X1    g725(.A(G162gat), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n887), .A2(new_n927), .A3(new_n311), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n904), .A2(new_n816), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n928), .B1(new_n929), .B2(new_n927), .ZN(G1347gat));
  NOR3_X1   g729(.A1(new_n745), .A2(new_n676), .A3(new_n550), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n842), .A2(new_n514), .A3(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(G169gat), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n932), .A2(new_n933), .A3(new_n681), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n850), .A2(new_n637), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT123), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n842), .A2(new_n588), .A3(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(new_n670), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n934), .B1(new_n933), .B2(new_n939), .ZN(G1348gat));
  OAI21_X1  g739(.A(G176gat), .B1(new_n932), .B2(new_n717), .ZN(new_n941));
  OR2_X1    g740(.A1(new_n717), .A2(G176gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n941), .B1(new_n937), .B2(new_n942), .ZN(G1349gat));
  AND3_X1   g742(.A1(new_n245), .A2(new_n354), .A3(new_n356), .ZN(new_n944));
  AOI22_X1  g743(.A1(new_n938), .A2(new_n944), .B1(KEYINPUT124), .B2(KEYINPUT60), .ZN(new_n945));
  OR2_X1    g744(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n946));
  OAI21_X1  g745(.A(G183gat), .B1(new_n932), .B2(new_n716), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n946), .B1(new_n945), .B2(new_n947), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n948), .A2(new_n949), .ZN(G1350gat));
  OAI21_X1  g749(.A(G190gat), .B1(new_n932), .B2(new_n311), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT61), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n938), .A2(new_n357), .A3(new_n816), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(G1351gat));
  NAND3_X1  g753(.A1(new_n697), .A2(new_n588), .A3(new_n637), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n917), .A2(new_n956), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n957), .A2(new_n481), .A3(new_n681), .ZN(new_n958));
  AOI211_X1 g757(.A(new_n550), .B(new_n514), .C1(new_n694), .C2(new_n696), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n849), .A2(new_n588), .A3(new_n839), .A4(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(G197gat), .B1(new_n961), .B2(new_n670), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n958), .A2(new_n962), .ZN(G1352gat));
  NOR2_X1   g762(.A1(new_n717), .A2(G204gat), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n960), .A2(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n967));
  AOI21_X1  g766(.A(KEYINPUT125), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT125), .ZN(new_n969));
  NOR4_X1   g768(.A1(new_n960), .A2(new_n969), .A3(KEYINPUT62), .A4(new_n965), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n842), .A2(new_n588), .A3(new_n959), .A4(new_n964), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(KEYINPUT62), .ZN(new_n973));
  AOI211_X1 g772(.A(new_n717), .B(new_n955), .C1(new_n915), .C2(new_n916), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n973), .B1(new_n974), .B2(new_n482), .ZN(new_n975));
  OAI21_X1  g774(.A(KEYINPUT126), .B1(new_n971), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n917), .A2(new_n349), .A3(new_n956), .ZN(new_n977));
  AOI22_X1  g776(.A1(new_n977), .A2(G204gat), .B1(KEYINPUT62), .B2(new_n972), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT126), .ZN(new_n979));
  OAI211_X1 g778(.A(new_n978), .B(new_n979), .C1(new_n968), .C2(new_n970), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n976), .A2(new_n980), .ZN(G1353gat));
  OAI21_X1  g780(.A(G211gat), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n982));
  INV_X1    g781(.A(new_n982), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n983), .B1(new_n957), .B2(new_n716), .ZN(new_n984));
  AND2_X1   g783(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n985));
  OR2_X1    g784(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OR3_X1    g785(.A1(new_n960), .A2(G211gat), .A3(new_n716), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n984), .A2(new_n985), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n986), .A2(new_n987), .A3(new_n988), .ZN(G1354gat));
  OAI21_X1  g788(.A(G218gat), .B1(new_n957), .B2(new_n311), .ZN(new_n990));
  OR3_X1    g789(.A1(new_n960), .A2(G218gat), .A3(new_n311), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(G1355gat));
endmodule


