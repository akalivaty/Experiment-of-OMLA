

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581;

  XNOR2_X1 U320 ( .A(KEYINPUT47), .B(KEYINPUT114), .ZN(n382) );
  INV_X1 U321 ( .A(n335), .ZN(n316) );
  XNOR2_X1 U322 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U323 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U324 ( .A(n426), .B(KEYINPUT55), .ZN(n427) );
  XNOR2_X1 U325 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U326 ( .A(n428), .B(n427), .ZN(n447) );
  INV_X1 U327 ( .A(G190GAT), .ZN(n449) );
  XNOR2_X1 U328 ( .A(n448), .B(KEYINPUT121), .ZN(n562) );
  XNOR2_X1 U329 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U330 ( .A(n452), .B(n451), .ZN(G1351GAT) );
  XOR2_X1 U331 ( .A(KEYINPUT21), .B(KEYINPUT90), .Z(n289) );
  XNOR2_X1 U332 ( .A(G218GAT), .B(KEYINPUT89), .ZN(n288) );
  XNOR2_X1 U333 ( .A(n289), .B(n288), .ZN(n290) );
  XOR2_X1 U334 ( .A(n290), .B(G211GAT), .Z(n292) );
  XNOR2_X1 U335 ( .A(G197GAT), .B(G204GAT), .ZN(n291) );
  XNOR2_X1 U336 ( .A(n292), .B(n291), .ZN(n389) );
  XOR2_X1 U337 ( .A(KEYINPUT75), .B(G162GAT), .Z(n352) );
  XOR2_X1 U338 ( .A(G78GAT), .B(G148GAT), .Z(n294) );
  XNOR2_X1 U339 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n293) );
  XNOR2_X1 U340 ( .A(n294), .B(n293), .ZN(n308) );
  XOR2_X1 U341 ( .A(n352), .B(n308), .Z(n296) );
  NAND2_X1 U342 ( .A1(G228GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U343 ( .A(n296), .B(n295), .ZN(n298) );
  XNOR2_X1 U344 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n297) );
  XNOR2_X1 U345 ( .A(n297), .B(KEYINPUT2), .ZN(n422) );
  XOR2_X1 U346 ( .A(n298), .B(n422), .Z(n300) );
  XNOR2_X1 U347 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n299) );
  XNOR2_X1 U348 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U349 ( .A(n301), .B(KEYINPUT22), .Z(n303) );
  XOR2_X1 U350 ( .A(G141GAT), .B(G22GAT), .Z(n366) );
  XNOR2_X1 U351 ( .A(G50GAT), .B(n366), .ZN(n302) );
  XNOR2_X1 U352 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U353 ( .A(n389), .B(n304), .ZN(n466) );
  XOR2_X1 U354 ( .A(KEYINPUT32), .B(KEYINPUT73), .Z(n306) );
  XNOR2_X1 U355 ( .A(G204GAT), .B(KEYINPUT74), .ZN(n305) );
  XOR2_X1 U356 ( .A(n306), .B(n305), .Z(n321) );
  XNOR2_X1 U357 ( .A(G176GAT), .B(G92GAT), .ZN(n307) );
  XNOR2_X1 U358 ( .A(n307), .B(G64GAT), .ZN(n397) );
  XNOR2_X1 U359 ( .A(n308), .B(n397), .ZN(n314) );
  XOR2_X1 U360 ( .A(KEYINPUT33), .B(KEYINPUT71), .Z(n310) );
  NAND2_X1 U361 ( .A1(G230GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U362 ( .A(n310), .B(n309), .ZN(n312) );
  INV_X1 U363 ( .A(KEYINPUT31), .ZN(n311) );
  XNOR2_X1 U364 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U365 ( .A(n314), .B(n313), .ZN(n319) );
  XOR2_X1 U366 ( .A(G120GAT), .B(G71GAT), .Z(n438) );
  XOR2_X1 U367 ( .A(G99GAT), .B(G85GAT), .Z(n351) );
  XNOR2_X1 U368 ( .A(n438), .B(n351), .ZN(n317) );
  XNOR2_X1 U369 ( .A(G57GAT), .B(KEYINPUT70), .ZN(n315) );
  XNOR2_X1 U370 ( .A(n315), .B(KEYINPUT13), .ZN(n335) );
  XNOR2_X1 U371 ( .A(n321), .B(n320), .ZN(n377) );
  XOR2_X1 U372 ( .A(KEYINPUT78), .B(KEYINPUT14), .Z(n323) );
  XNOR2_X1 U373 ( .A(KEYINPUT81), .B(KEYINPUT12), .ZN(n322) );
  XNOR2_X1 U374 ( .A(n323), .B(n322), .ZN(n340) );
  XOR2_X1 U375 ( .A(G78GAT), .B(G155GAT), .Z(n325) );
  XNOR2_X1 U376 ( .A(G22GAT), .B(G211GAT), .ZN(n324) );
  XNOR2_X1 U377 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U378 ( .A(G64GAT), .B(G71GAT), .Z(n327) );
  XNOR2_X1 U379 ( .A(G8GAT), .B(G127GAT), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U381 ( .A(n329), .B(n328), .Z(n334) );
  XOR2_X1 U382 ( .A(KEYINPUT79), .B(KEYINPUT15), .Z(n331) );
  NAND2_X1 U383 ( .A1(G231GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U384 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U385 ( .A(KEYINPUT80), .B(n332), .ZN(n333) );
  XNOR2_X1 U386 ( .A(n334), .B(n333), .ZN(n336) );
  XOR2_X1 U387 ( .A(n336), .B(n335), .Z(n338) );
  XOR2_X1 U388 ( .A(G15GAT), .B(G1GAT), .Z(n373) );
  XOR2_X1 U389 ( .A(G183GAT), .B(KEYINPUT77), .Z(n399) );
  XNOR2_X1 U390 ( .A(n373), .B(n399), .ZN(n337) );
  XNOR2_X1 U391 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U392 ( .A(n340), .B(n339), .Z(n548) );
  XOR2_X1 U393 ( .A(G29GAT), .B(KEYINPUT7), .Z(n342) );
  XNOR2_X1 U394 ( .A(G43GAT), .B(G36GAT), .ZN(n341) );
  XNOR2_X1 U395 ( .A(n342), .B(n341), .ZN(n344) );
  XOR2_X1 U396 ( .A(G50GAT), .B(KEYINPUT8), .Z(n343) );
  XNOR2_X1 U397 ( .A(n344), .B(n343), .ZN(n368) );
  INV_X1 U398 ( .A(n368), .ZN(n348) );
  XOR2_X1 U399 ( .A(KEYINPUT76), .B(KEYINPUT10), .Z(n346) );
  XNOR2_X1 U400 ( .A(G92GAT), .B(KEYINPUT9), .ZN(n345) );
  XNOR2_X1 U401 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U402 ( .A(n348), .B(n347), .ZN(n360) );
  XOR2_X1 U403 ( .A(KEYINPUT65), .B(G106GAT), .Z(n350) );
  XNOR2_X1 U404 ( .A(G190GAT), .B(G134GAT), .ZN(n349) );
  XNOR2_X1 U405 ( .A(n350), .B(n349), .ZN(n356) );
  XOR2_X1 U406 ( .A(KEYINPUT11), .B(n351), .Z(n354) );
  XNOR2_X1 U407 ( .A(G218GAT), .B(n352), .ZN(n353) );
  XNOR2_X1 U408 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U409 ( .A(n356), .B(n355), .Z(n358) );
  NAND2_X1 U410 ( .A1(G232GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U411 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U412 ( .A(n360), .B(n359), .ZN(n552) );
  XNOR2_X1 U413 ( .A(KEYINPUT36), .B(n552), .ZN(n579) );
  NOR2_X1 U414 ( .A1(n548), .A2(n579), .ZN(n361) );
  XOR2_X1 U415 ( .A(KEYINPUT45), .B(n361), .Z(n362) );
  NOR2_X1 U416 ( .A1(n377), .A2(n362), .ZN(n376) );
  XOR2_X1 U417 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n364) );
  NAND2_X1 U418 ( .A1(G229GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U419 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U420 ( .A(n366), .B(n365), .Z(n367) );
  XNOR2_X1 U421 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U422 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n370) );
  XNOR2_X1 U423 ( .A(G197GAT), .B(G113GAT), .ZN(n369) );
  XNOR2_X1 U424 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U425 ( .A(n372), .B(n371), .Z(n375) );
  XOR2_X1 U426 ( .A(G169GAT), .B(G8GAT), .Z(n400) );
  XNOR2_X1 U427 ( .A(n400), .B(n373), .ZN(n374) );
  XNOR2_X1 U428 ( .A(n375), .B(n374), .ZN(n567) );
  XOR2_X1 U429 ( .A(KEYINPUT69), .B(n567), .Z(n524) );
  NAND2_X1 U430 ( .A1(n376), .A2(n524), .ZN(n385) );
  XNOR2_X1 U431 ( .A(n377), .B(KEYINPUT41), .ZN(n544) );
  NOR2_X1 U432 ( .A1(n567), .A2(n544), .ZN(n378) );
  XNOR2_X1 U433 ( .A(n378), .B(KEYINPUT46), .ZN(n379) );
  INV_X1 U434 ( .A(n548), .ZN(n576) );
  NOR2_X1 U435 ( .A1(n379), .A2(n576), .ZN(n380) );
  XNOR2_X1 U436 ( .A(n380), .B(KEYINPUT113), .ZN(n381) );
  INV_X1 U437 ( .A(n552), .ZN(n534) );
  NOR2_X1 U438 ( .A1(n381), .A2(n534), .ZN(n383) );
  NAND2_X1 U439 ( .A1(n385), .A2(n384), .ZN(n386) );
  XNOR2_X1 U440 ( .A(n386), .B(KEYINPUT48), .ZN(n538) );
  XOR2_X1 U441 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n388) );
  NAND2_X1 U442 ( .A1(G226GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U443 ( .A(n388), .B(n387), .ZN(n390) );
  XOR2_X1 U444 ( .A(n390), .B(n389), .Z(n396) );
  XNOR2_X1 U445 ( .A(KEYINPUT87), .B(KEYINPUT19), .ZN(n391) );
  XNOR2_X1 U446 ( .A(n391), .B(KEYINPUT86), .ZN(n392) );
  XOR2_X1 U447 ( .A(n392), .B(KEYINPUT17), .Z(n394) );
  XNOR2_X1 U448 ( .A(KEYINPUT18), .B(G190GAT), .ZN(n393) );
  XNOR2_X1 U449 ( .A(n394), .B(n393), .ZN(n446) );
  XNOR2_X1 U450 ( .A(G36GAT), .B(n446), .ZN(n395) );
  XNOR2_X1 U451 ( .A(n396), .B(n395), .ZN(n398) );
  XOR2_X1 U452 ( .A(n398), .B(n397), .Z(n402) );
  XNOR2_X1 U453 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U454 ( .A(n402), .B(n401), .ZN(n459) );
  NAND2_X1 U455 ( .A1(n538), .A2(n459), .ZN(n404) );
  XOR2_X1 U456 ( .A(KEYINPUT54), .B(KEYINPUT118), .Z(n403) );
  XNOR2_X1 U457 ( .A(n404), .B(n403), .ZN(n425) );
  XOR2_X1 U458 ( .A(G85GAT), .B(G162GAT), .Z(n406) );
  XNOR2_X1 U459 ( .A(G29GAT), .B(G141GAT), .ZN(n405) );
  XNOR2_X1 U460 ( .A(n406), .B(n405), .ZN(n410) );
  XOR2_X1 U461 ( .A(KEYINPUT91), .B(KEYINPUT5), .Z(n408) );
  XNOR2_X1 U462 ( .A(G120GAT), .B(G148GAT), .ZN(n407) );
  XNOR2_X1 U463 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U464 ( .A(n410), .B(n409), .Z(n415) );
  XOR2_X1 U465 ( .A(KEYINPUT1), .B(G57GAT), .Z(n412) );
  NAND2_X1 U466 ( .A1(G225GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U467 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U468 ( .A(KEYINPUT6), .B(n413), .ZN(n414) );
  XNOR2_X1 U469 ( .A(n415), .B(n414), .ZN(n419) );
  XOR2_X1 U470 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n417) );
  XNOR2_X1 U471 ( .A(G1GAT), .B(KEYINPUT4), .ZN(n416) );
  XNOR2_X1 U472 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U473 ( .A(n419), .B(n418), .Z(n424) );
  XOR2_X1 U474 ( .A(G127GAT), .B(KEYINPUT0), .Z(n421) );
  XNOR2_X1 U475 ( .A(G113GAT), .B(G134GAT), .ZN(n420) );
  XNOR2_X1 U476 ( .A(n421), .B(n420), .ZN(n437) );
  XNOR2_X1 U477 ( .A(n437), .B(n422), .ZN(n423) );
  XNOR2_X1 U478 ( .A(n424), .B(n423), .ZN(n540) );
  NAND2_X1 U479 ( .A1(n425), .A2(n540), .ZN(n565) );
  NOR2_X1 U480 ( .A1(n466), .A2(n565), .ZN(n428) );
  XNOR2_X1 U481 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n426) );
  XOR2_X1 U482 ( .A(KEYINPUT64), .B(G176GAT), .Z(n430) );
  XNOR2_X1 U483 ( .A(G43GAT), .B(G99GAT), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U485 ( .A(G183GAT), .B(KEYINPUT83), .Z(n432) );
  XNOR2_X1 U486 ( .A(G15GAT), .B(KEYINPUT88), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U488 ( .A(n434), .B(n433), .Z(n444) );
  XOR2_X1 U489 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n436) );
  XNOR2_X1 U490 ( .A(G169GAT), .B(KEYINPUT85), .ZN(n435) );
  XNOR2_X1 U491 ( .A(n436), .B(n435), .ZN(n442) );
  XOR2_X1 U492 ( .A(n438), .B(n437), .Z(n440) );
  NAND2_X1 U493 ( .A1(G227GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U494 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U495 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U496 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U497 ( .A(n446), .B(n445), .ZN(n455) );
  NAND2_X1 U498 ( .A1(n447), .A2(n455), .ZN(n448) );
  NAND2_X1 U499 ( .A1(n562), .A2(n534), .ZN(n452) );
  XOR2_X1 U500 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n450) );
  NOR2_X1 U501 ( .A1(n524), .A2(n377), .ZN(n485) );
  XOR2_X1 U502 ( .A(KEYINPUT82), .B(KEYINPUT16), .Z(n454) );
  NAND2_X1 U503 ( .A1(n552), .A2(n576), .ZN(n453) );
  XNOR2_X1 U504 ( .A(n454), .B(n453), .ZN(n471) );
  INV_X1 U505 ( .A(n455), .ZN(n527) );
  NAND2_X1 U506 ( .A1(n466), .A2(n527), .ZN(n456) );
  XNOR2_X1 U507 ( .A(n456), .B(KEYINPUT26), .ZN(n566) );
  XNOR2_X1 U508 ( .A(n459), .B(KEYINPUT96), .ZN(n457) );
  XNOR2_X1 U509 ( .A(n457), .B(KEYINPUT27), .ZN(n467) );
  INV_X1 U510 ( .A(n467), .ZN(n458) );
  NOR2_X1 U511 ( .A1(n566), .A2(n458), .ZN(n541) );
  INV_X1 U512 ( .A(n459), .ZN(n513) );
  NOR2_X1 U513 ( .A1(n527), .A2(n513), .ZN(n460) );
  NOR2_X1 U514 ( .A1(n466), .A2(n460), .ZN(n461) );
  XOR2_X1 U515 ( .A(KEYINPUT25), .B(n461), .Z(n462) );
  NOR2_X1 U516 ( .A1(n541), .A2(n462), .ZN(n463) );
  XNOR2_X1 U517 ( .A(KEYINPUT97), .B(n463), .ZN(n464) );
  NAND2_X1 U518 ( .A1(n464), .A2(n540), .ZN(n470) );
  XOR2_X1 U519 ( .A(KEYINPUT66), .B(KEYINPUT28), .Z(n465) );
  XNOR2_X1 U520 ( .A(n466), .B(n465), .ZN(n521) );
  NAND2_X1 U521 ( .A1(n467), .A2(n521), .ZN(n468) );
  NOR2_X1 U522 ( .A1(n540), .A2(n468), .ZN(n525) );
  NAND2_X1 U523 ( .A1(n525), .A2(n527), .ZN(n469) );
  NAND2_X1 U524 ( .A1(n470), .A2(n469), .ZN(n482) );
  AND2_X1 U525 ( .A1(n471), .A2(n482), .ZN(n499) );
  NAND2_X1 U526 ( .A1(n485), .A2(n499), .ZN(n480) );
  NOR2_X1 U527 ( .A1(n540), .A2(n480), .ZN(n473) );
  XNOR2_X1 U528 ( .A(KEYINPUT34), .B(KEYINPUT98), .ZN(n472) );
  XNOR2_X1 U529 ( .A(n473), .B(n472), .ZN(n474) );
  XOR2_X1 U530 ( .A(G1GAT), .B(n474), .Z(G1324GAT) );
  NOR2_X1 U531 ( .A1(n513), .A2(n480), .ZN(n476) );
  XNOR2_X1 U532 ( .A(G8GAT), .B(KEYINPUT99), .ZN(n475) );
  XNOR2_X1 U533 ( .A(n476), .B(n475), .ZN(G1325GAT) );
  NOR2_X1 U534 ( .A1(n527), .A2(n480), .ZN(n478) );
  XNOR2_X1 U535 ( .A(KEYINPUT100), .B(KEYINPUT35), .ZN(n477) );
  XNOR2_X1 U536 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U537 ( .A(G15GAT), .B(n479), .ZN(G1326GAT) );
  NOR2_X1 U538 ( .A1(n521), .A2(n480), .ZN(n481) );
  XOR2_X1 U539 ( .A(G22GAT), .B(n481), .Z(G1327GAT) );
  NOR2_X1 U540 ( .A1(n579), .A2(n576), .ZN(n483) );
  NAND2_X1 U541 ( .A1(n483), .A2(n482), .ZN(n484) );
  XNOR2_X1 U542 ( .A(KEYINPUT37), .B(n484), .ZN(n510) );
  NAND2_X1 U543 ( .A1(n510), .A2(n485), .ZN(n487) );
  XNOR2_X1 U544 ( .A(KEYINPUT102), .B(KEYINPUT38), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n487), .B(n486), .ZN(n496) );
  NOR2_X1 U546 ( .A1(n540), .A2(n496), .ZN(n490) );
  XOR2_X1 U547 ( .A(KEYINPUT101), .B(KEYINPUT39), .Z(n488) );
  XNOR2_X1 U548 ( .A(G29GAT), .B(n488), .ZN(n489) );
  XNOR2_X1 U549 ( .A(n490), .B(n489), .ZN(G1328GAT) );
  NOR2_X1 U550 ( .A1(n513), .A2(n496), .ZN(n492) );
  XNOR2_X1 U551 ( .A(G36GAT), .B(KEYINPUT103), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(G1329GAT) );
  NOR2_X1 U553 ( .A1(n527), .A2(n496), .ZN(n494) );
  XNOR2_X1 U554 ( .A(KEYINPUT104), .B(KEYINPUT40), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U556 ( .A(G43GAT), .B(n495), .Z(G1330GAT) );
  NOR2_X1 U557 ( .A1(n521), .A2(n496), .ZN(n498) );
  XNOR2_X1 U558 ( .A(G50GAT), .B(KEYINPUT105), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n498), .B(n497), .ZN(G1331GAT) );
  INV_X1 U560 ( .A(n544), .ZN(n557) );
  AND2_X1 U561 ( .A1(n567), .A2(n557), .ZN(n509) );
  NAND2_X1 U562 ( .A1(n509), .A2(n499), .ZN(n506) );
  NOR2_X1 U563 ( .A1(n540), .A2(n506), .ZN(n501) );
  XNOR2_X1 U564 ( .A(KEYINPUT106), .B(KEYINPUT42), .ZN(n500) );
  XNOR2_X1 U565 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U566 ( .A(G57GAT), .B(n502), .Z(G1332GAT) );
  NOR2_X1 U567 ( .A1(n513), .A2(n506), .ZN(n504) );
  XNOR2_X1 U568 ( .A(G64GAT), .B(KEYINPUT107), .ZN(n503) );
  XNOR2_X1 U569 ( .A(n504), .B(n503), .ZN(G1333GAT) );
  NOR2_X1 U570 ( .A1(n527), .A2(n506), .ZN(n505) );
  XOR2_X1 U571 ( .A(G71GAT), .B(n505), .Z(G1334GAT) );
  NOR2_X1 U572 ( .A1(n521), .A2(n506), .ZN(n508) );
  XNOR2_X1 U573 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n507) );
  XNOR2_X1 U574 ( .A(n508), .B(n507), .ZN(G1335GAT) );
  NAND2_X1 U575 ( .A1(n510), .A2(n509), .ZN(n520) );
  NOR2_X1 U576 ( .A1(n540), .A2(n520), .ZN(n511) );
  XOR2_X1 U577 ( .A(G85GAT), .B(n511), .Z(n512) );
  XNOR2_X1 U578 ( .A(KEYINPUT108), .B(n512), .ZN(G1336GAT) );
  NOR2_X1 U579 ( .A1(n513), .A2(n520), .ZN(n515) );
  XNOR2_X1 U580 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U582 ( .A(G92GAT), .B(n516), .ZN(G1337GAT) );
  NOR2_X1 U583 ( .A1(n527), .A2(n520), .ZN(n517) );
  XOR2_X1 U584 ( .A(G99GAT), .B(n517), .Z(G1338GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT111), .B(KEYINPUT44), .Z(n519) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(KEYINPUT112), .ZN(n518) );
  XNOR2_X1 U587 ( .A(n519), .B(n518), .ZN(n523) );
  NOR2_X1 U588 ( .A1(n521), .A2(n520), .ZN(n522) );
  XOR2_X1 U589 ( .A(n523), .B(n522), .Z(G1339GAT) );
  INV_X1 U590 ( .A(n524), .ZN(n555) );
  NAND2_X1 U591 ( .A1(n538), .A2(n525), .ZN(n526) );
  NOR2_X1 U592 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U593 ( .A(KEYINPUT115), .B(n528), .Z(n535) );
  NAND2_X1 U594 ( .A1(n555), .A2(n535), .ZN(n529) );
  XNOR2_X1 U595 ( .A(n529), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U596 ( .A(G120GAT), .B(KEYINPUT49), .Z(n531) );
  NAND2_X1 U597 ( .A1(n535), .A2(n557), .ZN(n530) );
  XNOR2_X1 U598 ( .A(n531), .B(n530), .ZN(G1341GAT) );
  NAND2_X1 U599 ( .A1(n576), .A2(n535), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n532), .B(KEYINPUT50), .ZN(n533) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n533), .ZN(G1342GAT) );
  XOR2_X1 U602 ( .A(G134GAT), .B(KEYINPUT51), .Z(n537) );
  NAND2_X1 U603 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n537), .B(n536), .ZN(G1343GAT) );
  INV_X1 U605 ( .A(n538), .ZN(n539) );
  NOR2_X1 U606 ( .A1(n540), .A2(n539), .ZN(n542) );
  NAND2_X1 U607 ( .A1(n542), .A2(n541), .ZN(n551) );
  NOR2_X1 U608 ( .A1(n567), .A2(n551), .ZN(n543) );
  XOR2_X1 U609 ( .A(G141GAT), .B(n543), .Z(G1344GAT) );
  NOR2_X1 U610 ( .A1(n544), .A2(n551), .ZN(n546) );
  XNOR2_X1 U611 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(n547), .ZN(G1345GAT) );
  NOR2_X1 U614 ( .A1(n548), .A2(n551), .ZN(n549) );
  XOR2_X1 U615 ( .A(KEYINPUT116), .B(n549), .Z(n550) );
  XNOR2_X1 U616 ( .A(G155GAT), .B(n550), .ZN(G1346GAT) );
  NOR2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n554) );
  XNOR2_X1 U618 ( .A(G162GAT), .B(KEYINPUT117), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(G1347GAT) );
  NAND2_X1 U620 ( .A1(n555), .A2(n562), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n556), .B(G169GAT), .ZN(G1348GAT) );
  XNOR2_X1 U622 ( .A(KEYINPUT122), .B(KEYINPUT57), .ZN(n561) );
  XOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT56), .Z(n559) );
  NAND2_X1 U624 ( .A1(n562), .A2(n557), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n561), .B(n560), .ZN(G1349GAT) );
  XOR2_X1 U627 ( .A(G183GAT), .B(KEYINPUT123), .Z(n564) );
  NAND2_X1 U628 ( .A1(n562), .A2(n576), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(G1350GAT) );
  NOR2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n575) );
  INV_X1 U631 ( .A(n575), .ZN(n578) );
  NOR2_X1 U632 ( .A1(n567), .A2(n578), .ZN(n569) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n571) );
  XOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n573) );
  NAND2_X1 U638 ( .A1(n575), .A2(n377), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(n574), .ZN(G1353GAT) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n577), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U644 ( .A(KEYINPUT62), .B(n580), .Z(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

