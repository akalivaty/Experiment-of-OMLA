//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986;
  INV_X1    g000(.A(KEYINPUT20), .ZN(new_n187));
  NOR2_X1   g001(.A1(G475), .A2(G902), .ZN(new_n188));
  NOR2_X1   g002(.A1(G237), .A2(G953), .ZN(new_n189));
  AND3_X1   g003(.A1(new_n189), .A2(G143), .A3(G214), .ZN(new_n190));
  AOI21_X1  g004(.A(G143), .B1(new_n189), .B2(G214), .ZN(new_n191));
  OAI21_X1  g005(.A(G131), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT17), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n189), .A2(G214), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G131), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n189), .A2(G143), .A3(G214), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n197), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  AND2_X1   g014(.A1(new_n192), .A2(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n194), .B1(new_n201), .B2(new_n193), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT16), .ZN(new_n204));
  INV_X1    g018(.A(G140), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G125), .ZN(new_n206));
  OR2_X1    g020(.A1(KEYINPUT75), .A2(G125), .ZN(new_n207));
  NAND2_X1  g021(.A1(KEYINPUT75), .A2(G125), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI211_X1 g023(.A(KEYINPUT76), .B(new_n206), .C1(new_n209), .C2(new_n205), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT76), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n207), .A2(new_n211), .A3(G140), .A4(new_n208), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n204), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n209), .A2(new_n204), .A3(new_n205), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n203), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  AND2_X1   g030(.A1(KEYINPUT75), .A2(G125), .ZN(new_n217));
  NOR2_X1   g031(.A1(KEYINPUT75), .A2(G125), .ZN(new_n218));
  NOR3_X1   g032(.A1(new_n217), .A2(new_n218), .A3(new_n205), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n206), .A2(KEYINPUT76), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n212), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT16), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(G146), .A3(new_n214), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n202), .A2(new_n216), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n197), .A2(new_n199), .ZN(new_n225));
  NAND2_X1  g039(.A1(KEYINPUT18), .A2(G131), .ZN(new_n226));
  OR3_X1    g040(.A1(new_n225), .A2(KEYINPUT91), .A3(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n226), .B1(new_n225), .B2(KEYINPUT91), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(G125), .B(G140), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(new_n203), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n231), .B1(new_n221), .B2(new_n203), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(G113), .B(G122), .ZN(new_n234));
  INV_X1    g048(.A(G104), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g050(.A(new_n236), .B(KEYINPUT93), .Z(new_n237));
  AND3_X1   g051(.A1(new_n224), .A2(new_n233), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT92), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT19), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n239), .B1(new_n221), .B2(new_n240), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n210), .A2(KEYINPUT92), .A3(KEYINPUT19), .A4(new_n212), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n230), .A2(new_n240), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n241), .A2(new_n203), .A3(new_n242), .A4(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n201), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n223), .A3(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n236), .B1(new_n246), .B2(new_n233), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n187), .B(new_n188), .C1(new_n238), .C2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT94), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n224), .A2(new_n233), .A3(new_n237), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n223), .A2(new_n245), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n251), .A2(new_n244), .B1(new_n232), .B2(new_n229), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n250), .B1(new_n252), .B2(new_n236), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT94), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n253), .A2(new_n254), .A3(new_n187), .A4(new_n188), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n188), .B1(new_n238), .B2(new_n247), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(KEYINPUT20), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n249), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(G234), .A2(G237), .ZN(new_n259));
  INV_X1    g073(.A(G953), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n259), .A2(G952), .A3(new_n260), .ZN(new_n261));
  AND3_X1   g075(.A1(new_n259), .A2(G902), .A3(G953), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT21), .B(G898), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT9), .B(G234), .ZN(new_n266));
  INV_X1    g080(.A(G217), .ZN(new_n267));
  NOR3_X1   g081(.A1(new_n266), .A2(new_n267), .A3(G953), .ZN(new_n268));
  INV_X1    g082(.A(G122), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G116), .ZN(new_n270));
  INV_X1    g084(.A(G116), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G122), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G107), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n273), .B(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n196), .A2(G128), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT13), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G128), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G143), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n276), .A2(new_n277), .ZN(new_n282));
  OAI21_X1  g096(.A(G134), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n276), .A2(new_n280), .ZN(new_n284));
  INV_X1    g098(.A(G134), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n275), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n284), .B(new_n285), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n273), .A2(new_n274), .ZN(new_n289));
  OR2_X1    g103(.A1(new_n272), .A2(KEYINPUT14), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n272), .A2(KEYINPUT14), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n290), .A2(new_n291), .A3(new_n270), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G107), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n288), .A2(new_n289), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n268), .B1(new_n287), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n287), .A2(new_n294), .A3(new_n268), .ZN(new_n297));
  AOI21_X1  g111(.A(G902), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G478), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n299), .A2(KEYINPUT15), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  OR2_X1    g115(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n298), .A2(new_n301), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G902), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n236), .B1(new_n224), .B2(new_n233), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n306), .B1(new_n238), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G475), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n258), .A2(new_n265), .A3(new_n305), .A4(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT95), .ZN(new_n311));
  OR2_X1    g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n311), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(G110), .B(G140), .ZN(new_n315));
  INV_X1    g129(.A(G227), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n316), .A2(G953), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n315), .B(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n203), .A2(G143), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n196), .A2(G146), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(G128), .ZN(new_n322));
  OR2_X1    g136(.A1(KEYINPUT68), .A2(KEYINPUT1), .ZN(new_n323));
  NAND2_X1  g137(.A1(KEYINPUT68), .A2(KEYINPUT1), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT69), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  AND2_X1   g140(.A1(KEYINPUT68), .A2(KEYINPUT1), .ZN(new_n327));
  NOR2_X1   g141(.A1(KEYINPUT68), .A2(KEYINPUT1), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(G143), .B(G146), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT69), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n329), .A2(new_n330), .A3(new_n331), .A4(G128), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n326), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n320), .A2(new_n321), .ZN(new_n334));
  AOI22_X1  g148(.A1(new_n323), .A2(new_n324), .B1(G143), .B2(new_n203), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n334), .B1(new_n335), .B2(new_n279), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT82), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n338), .B1(new_n274), .B2(G104), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n274), .A2(G104), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n235), .A2(KEYINPUT82), .A3(G107), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G101), .ZN(new_n343));
  INV_X1    g157(.A(G101), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n235), .A2(G107), .ZN(new_n345));
  AND3_X1   g159(.A1(new_n274), .A2(KEYINPUT3), .A3(G104), .ZN(new_n346));
  AOI21_X1  g160(.A(KEYINPUT3), .B1(new_n274), .B2(G104), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n344), .B(new_n345), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n337), .A2(KEYINPUT10), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT10), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n203), .A2(G143), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT1), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n354), .B1(new_n330), .B2(G128), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n355), .B1(new_n326), .B2(new_n332), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n352), .B1(new_n356), .B2(new_n349), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G101), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n359), .A2(KEYINPUT4), .A3(new_n348), .ZN(new_n360));
  NOR2_X1   g174(.A1(KEYINPUT0), .A2(G128), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT64), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n334), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(KEYINPUT0), .A2(G128), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n364), .B1(new_n361), .B2(KEYINPUT64), .ZN(new_n365));
  OAI22_X1  g179(.A1(new_n363), .A2(new_n365), .B1(new_n364), .B2(new_n334), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  XOR2_X1   g181(.A(KEYINPUT81), .B(KEYINPUT4), .Z(new_n368));
  NAND3_X1  g182(.A1(new_n358), .A2(G101), .A3(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n360), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n351), .A2(new_n357), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT11), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n372), .B1(new_n285), .B2(G137), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n285), .A2(G137), .ZN(new_n374));
  INV_X1    g188(.A(G137), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n375), .A2(KEYINPUT11), .A3(G134), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n373), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT66), .ZN(new_n378));
  AND3_X1   g192(.A1(new_n377), .A2(new_n378), .A3(G131), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n378), .B1(new_n377), .B2(G131), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n373), .A2(new_n376), .A3(new_n198), .A4(new_n374), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT65), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n382), .B(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(KEYINPUT83), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n377), .A2(G131), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT66), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n377), .A2(new_n378), .A3(G131), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n376), .A2(new_n374), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n390), .A2(new_n383), .A3(new_n198), .A4(new_n373), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n382), .A2(KEYINPUT65), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT83), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n389), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n385), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n319), .B1(new_n371), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT87), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI211_X1 g213(.A(KEYINPUT87), .B(new_n319), .C1(new_n371), .C2(new_n396), .ZN(new_n400));
  AND2_X1   g214(.A1(new_n382), .A2(KEYINPUT65), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n382), .A2(KEYINPUT65), .ZN(new_n402));
  OAI22_X1  g216(.A1(new_n380), .A2(new_n379), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n371), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n399), .A2(new_n400), .A3(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n371), .A2(new_n396), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n333), .A2(new_n349), .A3(new_n336), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n407), .B1(new_n349), .B2(new_n356), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT85), .ZN(new_n409));
  XOR2_X1   g223(.A(KEYINPUT84), .B(KEYINPUT12), .Z(new_n410));
  AOI21_X1  g224(.A(new_n410), .B1(new_n389), .B2(new_n393), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n408), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n409), .B1(new_n408), .B2(new_n411), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n333), .A2(new_n349), .A3(new_n336), .ZN(new_n415));
  INV_X1    g229(.A(new_n355), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n349), .B1(new_n333), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(KEYINPUT86), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT86), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n407), .B(new_n419), .C1(new_n349), .C2(new_n356), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n418), .A2(new_n403), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT12), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n406), .B1(new_n414), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n318), .B(KEYINPUT80), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n405), .B(G469), .C1(new_n424), .C2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G469), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n397), .B1(new_n414), .B2(new_n423), .ZN(new_n428));
  OR2_X1    g242(.A1(new_n371), .A2(new_n396), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n319), .B1(new_n429), .B2(new_n404), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n427), .B(new_n306), .C1(new_n428), .C2(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n427), .A2(new_n306), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n426), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(G221), .B1(new_n266), .B2(G902), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(KEYINPUT79), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT88), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT88), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n434), .A2(new_n439), .A3(new_n436), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G119), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G116), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n271), .A2(G119), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(KEYINPUT2), .B(G113), .ZN(new_n446));
  OR2_X1    g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n446), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n360), .A2(new_n369), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n443), .A2(new_n444), .A3(KEYINPUT5), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n451), .B(G113), .C1(KEYINPUT5), .C2(new_n443), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n350), .A2(new_n447), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(G110), .B(G122), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(KEYINPUT89), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n450), .A2(new_n453), .A3(new_n456), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(KEYINPUT6), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n209), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n337), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n366), .A2(new_n461), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n260), .A2(G224), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n462), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n209), .B1(new_n333), .B2(new_n336), .ZN(new_n467));
  OAI211_X1 g281(.A(G224), .B(new_n260), .C1(new_n467), .C2(new_n463), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT6), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n454), .A2(new_n470), .A3(new_n457), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n460), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT7), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n465), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n466), .A2(new_n468), .A3(new_n474), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n462), .A2(new_n464), .A3(new_n473), .A4(new_n465), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n452), .A2(new_n447), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(new_n349), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n456), .B(KEYINPUT8), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n475), .A2(new_n459), .A3(new_n476), .A4(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n472), .A2(new_n306), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(G210), .B1(G237), .B2(G902), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n472), .A2(new_n481), .A3(new_n306), .A4(new_n483), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(G214), .B1(G237), .B2(G902), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT90), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n488), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n492), .B1(new_n485), .B2(new_n486), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT90), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n314), .A2(new_n441), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT78), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n367), .B1(new_n381), .B2(new_n384), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT67), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n499), .B1(new_n375), .B2(G134), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n285), .A2(G137), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n375), .A2(G134), .ZN(new_n503));
  OAI21_X1  g317(.A(G131), .B1(new_n503), .B2(new_n499), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n505), .B1(new_n391), .B2(new_n392), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n337), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT30), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n498), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n508), .B1(new_n498), .B2(new_n507), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n449), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AOI22_X1  g325(.A1(new_n403), .A2(new_n367), .B1(new_n337), .B2(new_n506), .ZN(new_n512));
  INV_X1    g326(.A(new_n449), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n189), .A2(G210), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n515), .B(KEYINPUT27), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT26), .B(G101), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n516), .B(new_n517), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n511), .A2(KEYINPUT70), .A3(new_n514), .A4(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT31), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n520), .A2(KEYINPUT70), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n521), .A2(KEYINPUT31), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  AND2_X1   g337(.A1(new_n337), .A2(new_n506), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n366), .B1(new_n389), .B2(new_n393), .ZN(new_n525));
  NOR3_X1   g339(.A1(new_n524), .A2(new_n525), .A3(new_n449), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT30), .B1(new_n524), .B2(new_n525), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n498), .A2(new_n507), .A3(new_n508), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n526), .B1(new_n529), .B2(new_n449), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n530), .A2(KEYINPUT70), .A3(KEYINPUT31), .A4(new_n518), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n523), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT28), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n514), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT71), .B1(new_n512), .B2(new_n513), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n498), .A2(new_n507), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT71), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(new_n537), .A3(new_n449), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n526), .B1(new_n535), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n534), .B1(new_n539), .B2(new_n533), .ZN(new_n540));
  INV_X1    g354(.A(new_n518), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n532), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT32), .ZN(new_n544));
  NOR2_X1   g358(.A1(G472), .A2(G902), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  AOI22_X1  g360(.A1(new_n523), .A2(new_n531), .B1(new_n540), .B2(new_n541), .ZN(new_n547));
  INV_X1    g361(.A(new_n545), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT32), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n511), .ZN(new_n551));
  OAI211_X1 g365(.A(KEYINPUT72), .B(new_n541), .C1(new_n551), .C2(new_n526), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT72), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n553), .B1(new_n530), .B2(new_n518), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n534), .B(new_n518), .C1(new_n539), .C2(new_n533), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT29), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n552), .A2(new_n554), .A3(new_n555), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n536), .A2(new_n449), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT73), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(new_n514), .A3(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n536), .A2(KEYINPUT73), .A3(new_n449), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n560), .A2(KEYINPUT28), .A3(new_n561), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n562), .A2(KEYINPUT29), .A3(new_n534), .A4(new_n518), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n557), .A2(new_n306), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(G472), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n550), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n267), .B1(G234), .B2(new_n306), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n216), .A2(new_n223), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT24), .B(G110), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(KEYINPUT74), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n442), .A2(G128), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n442), .A2(G128), .ZN(new_n574));
  AND2_X1   g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n279), .A2(KEYINPUT23), .A3(G119), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n577), .B(new_n574), .C1(new_n572), .C2(KEYINPUT23), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(G110), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n569), .A2(new_n581), .ZN(new_n582));
  OAI22_X1  g396(.A1(new_n571), .A2(new_n575), .B1(G110), .B2(new_n578), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n223), .A2(new_n231), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n260), .A2(G221), .A3(G234), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(KEYINPUT77), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT22), .B(G137), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n586), .B(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n582), .A2(new_n584), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n588), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n580), .B1(new_n216), .B2(new_n223), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n223), .A2(new_n231), .A3(new_n583), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n589), .A2(new_n593), .A3(new_n306), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT25), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n589), .A2(new_n593), .A3(KEYINPUT25), .A4(new_n306), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n568), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n589), .A2(new_n593), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n567), .A2(G902), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n497), .B1(new_n566), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n546), .A2(new_n549), .B1(new_n564), .B2(G472), .ZN(new_n603));
  INV_X1    g417(.A(new_n601), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n603), .A2(KEYINPUT78), .A3(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n496), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G101), .ZN(G3));
  OAI21_X1  g421(.A(G472), .B1(new_n547), .B2(G902), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n608), .B1(new_n548), .B2(new_n547), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n609), .A2(new_n604), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n610), .A2(new_n441), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n258), .A2(new_n309), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT33), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n296), .A2(new_n613), .A3(new_n297), .ZN(new_n614));
  INV_X1    g428(.A(new_n297), .ZN(new_n615));
  OAI21_X1  g429(.A(KEYINPUT33), .B1(new_n615), .B2(new_n295), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n614), .A2(new_n616), .A3(G478), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n298), .A2(new_n299), .ZN(new_n618));
  NAND2_X1  g432(.A1(G478), .A2(G902), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n612), .A2(new_n493), .A3(new_n265), .A4(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n611), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT96), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT34), .B(G104), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G6));
  AOI22_X1  g441(.A1(new_n257), .A2(new_n248), .B1(new_n308), .B2(G475), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n493), .A2(new_n304), .A3(new_n265), .A4(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n611), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT35), .B(G107), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G9));
  NAND2_X1  g447(.A1(new_n582), .A2(new_n584), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n590), .A2(KEYINPUT36), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n600), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n596), .A2(new_n597), .ZN(new_n638));
  OAI211_X1 g452(.A(KEYINPUT97), .B(new_n637), .C1(new_n638), .C2(new_n568), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT97), .ZN(new_n640));
  INV_X1    g454(.A(new_n637), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n640), .B1(new_n641), .B2(new_n598), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n609), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n496), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT37), .B(G110), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G12));
  NAND3_X1  g461(.A1(new_n639), .A2(new_n642), .A3(new_n493), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n648), .B1(new_n550), .B2(new_n565), .ZN(new_n649));
  INV_X1    g463(.A(new_n261), .ZN(new_n650));
  INV_X1    g464(.A(new_n262), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n650), .B1(new_n651), .B2(G900), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT98), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n628), .A2(new_n304), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n655), .B1(new_n438), .B2(new_n440), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n649), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G128), .ZN(G30));
  XOR2_X1   g472(.A(new_n653), .B(KEYINPUT39), .Z(new_n659));
  NAND2_X1  g473(.A1(new_n441), .A2(new_n659), .ZN(new_n660));
  OR2_X1    g474(.A1(new_n660), .A2(KEYINPUT40), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(KEYINPUT40), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n560), .A2(new_n541), .A3(new_n561), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n663), .A2(KEYINPUT99), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n530), .A2(new_n518), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n663), .A2(KEYINPUT99), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g481(.A(G472), .B1(new_n667), .B2(G902), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n550), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n487), .B(KEYINPUT38), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n671), .A2(new_n304), .A3(new_n612), .A4(new_n488), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n641), .A2(new_n598), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n670), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n661), .A2(new_n662), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G143), .ZN(G45));
  NAND3_X1  g491(.A1(new_n612), .A2(new_n621), .A3(new_n654), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n678), .B1(new_n438), .B2(new_n440), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n649), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(KEYINPUT100), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT100), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n649), .A2(new_n679), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G146), .ZN(G48));
  NOR2_X1   g499(.A1(new_n603), .A2(new_n604), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n428), .A2(new_n430), .ZN(new_n687));
  OAI21_X1  g501(.A(G469), .B1(new_n687), .B2(G902), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n688), .A2(new_n435), .A3(new_n431), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n622), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT41), .B(G113), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G15));
  NOR2_X1   g507(.A1(new_n629), .A2(new_n689), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n686), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G116), .ZN(G18));
  AOI21_X1  g510(.A(new_n689), .B1(new_n312), .B2(new_n313), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n649), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(KEYINPUT101), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT101), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n697), .A2(new_n649), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G119), .ZN(G21));
  AND2_X1   g517(.A1(new_n523), .A2(new_n531), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n518), .B1(new_n562), .B2(new_n534), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n545), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  AND2_X1   g520(.A1(new_n608), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n612), .A2(new_n493), .A3(new_n304), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n708), .A2(new_n264), .ZN(new_n709));
  INV_X1    g523(.A(new_n689), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n707), .A2(new_n709), .A3(new_n601), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G122), .ZN(G24));
  AOI211_X1 g526(.A(new_n653), .B(new_n620), .C1(new_n258), .C2(new_n309), .ZN(new_n713));
  AND4_X1   g527(.A1(new_n608), .A2(new_n713), .A3(new_n674), .A4(new_n706), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n689), .A2(new_n489), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G125), .ZN(G27));
  NOR2_X1   g531(.A1(new_n487), .A2(new_n492), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n718), .A2(new_n435), .A3(new_n434), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n603), .A2(new_n604), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g534(.A(KEYINPUT42), .B1(new_n720), .B2(new_n713), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n550), .A2(KEYINPUT102), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT102), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n546), .A2(new_n549), .A3(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n722), .A2(new_n565), .A3(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT42), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n719), .A2(new_n726), .A3(new_n678), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n725), .A2(new_n601), .A3(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT103), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n725), .A2(KEYINPUT103), .A3(new_n601), .A4(new_n727), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n721), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(KEYINPUT104), .B(G131), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G33));
  INV_X1    g548(.A(new_n655), .ZN(new_n735));
  AOI21_X1  g549(.A(KEYINPUT105), .B1(new_n720), .B2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n719), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n566), .A2(new_n601), .A3(new_n735), .A4(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT105), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OR2_X1    g554(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G134), .ZN(G36));
  INV_X1    g556(.A(new_n718), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n258), .A2(new_n309), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n621), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT43), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n747), .A2(new_n609), .A3(new_n674), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n743), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n750), .B1(new_n749), .B2(new_n748), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n751), .A2(KEYINPUT107), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(KEYINPUT107), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n405), .B1(new_n424), .B2(new_n425), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n755));
  OR2_X1    g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n427), .B1(new_n754), .B2(new_n755), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OR2_X1    g572(.A1(new_n758), .A2(new_n432), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT46), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n431), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n759), .A2(new_n760), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n435), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT106), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n765), .A2(new_n766), .A3(new_n659), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n766), .B1(new_n765), .B2(new_n659), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n752), .B(new_n753), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G137), .ZN(G39));
  INV_X1    g584(.A(KEYINPUT47), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n764), .A2(new_n771), .ZN(new_n772));
  OAI211_X1 g586(.A(KEYINPUT47), .B(new_n435), .C1(new_n762), .C2(new_n763), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n678), .A2(new_n601), .A3(new_n743), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n774), .A2(new_n603), .A3(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G140), .ZN(G42));
  AND2_X1   g591(.A1(new_n688), .A2(new_n431), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT49), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n601), .A2(new_n488), .A3(new_n436), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n671), .A2(new_n780), .A3(new_n745), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n670), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n491), .A2(new_n265), .A3(new_n494), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n612), .A2(new_n620), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n784), .B1(new_n304), .B2(new_n612), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n786), .A2(new_n441), .A3(new_n610), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n566), .B(new_n601), .C1(new_n690), .C2(new_n694), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n787), .A2(new_n711), .A3(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n789), .A2(new_n702), .A3(new_n606), .A4(new_n645), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n714), .A2(new_n737), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT108), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n304), .A2(new_n653), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n628), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n792), .B1(new_n743), .B2(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n718), .A2(KEYINPUT108), .A3(new_n628), .A4(new_n793), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n643), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(new_n566), .A3(new_n441), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n791), .B(new_n798), .C1(new_n736), .C2(new_n740), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n790), .A2(new_n732), .A3(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT110), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n649), .A2(new_n679), .A3(new_n682), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n682), .B1(new_n649), .B2(new_n679), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n708), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n434), .A2(new_n435), .A3(new_n654), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n669), .A2(new_n673), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n657), .A2(new_n807), .A3(new_n716), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n801), .B1(new_n804), .B2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n657), .A2(new_n807), .A3(new_n716), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n684), .A2(new_n811), .A3(KEYINPUT110), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n809), .A2(new_n810), .A3(new_n812), .ZN(new_n813));
  AOI22_X1  g627(.A1(new_n649), .A2(new_n656), .B1(new_n714), .B2(new_n715), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n814), .B(new_n807), .C1(new_n802), .C2(new_n803), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT109), .B1(new_n815), .B2(new_n810), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT109), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n684), .A2(new_n811), .A3(new_n817), .A4(KEYINPUT52), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n800), .B1(new_n813), .B2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n820), .A2(KEYINPUT111), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n809), .A2(new_n812), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT52), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n809), .A2(new_n812), .A3(new_n810), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(KEYINPUT53), .A3(new_n800), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n822), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT111), .B1(new_n820), .B2(new_n821), .ZN(new_n829));
  OAI21_X1  g643(.A(KEYINPUT54), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT112), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT51), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n707), .A2(new_n601), .ZN(new_n833));
  AND4_X1   g647(.A1(new_n261), .A2(new_n833), .A3(new_n747), .A4(new_n710), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n671), .A2(new_n488), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT50), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n834), .A2(KEYINPUT50), .A3(new_n835), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AND4_X1   g654(.A1(new_n261), .A2(new_n747), .A3(new_n710), .A4(new_n718), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n707), .A2(new_n674), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n710), .A2(new_n601), .A3(new_n261), .A4(new_n718), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n844), .A2(new_n669), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n612), .A2(new_n621), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n841), .A2(new_n843), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n840), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT113), .ZN(new_n849));
  INV_X1    g663(.A(new_n778), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n772), .B(new_n773), .C1(new_n436), .C2(new_n850), .ZN(new_n851));
  AND4_X1   g665(.A1(new_n261), .A2(new_n833), .A3(new_n747), .A4(new_n718), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n848), .A2(KEYINPUT113), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n832), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(G952), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n744), .A2(new_n620), .ZN(new_n858));
  AOI211_X1 g672(.A(new_n857), .B(G953), .C1(new_n845), .C2(new_n858), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n834), .A2(KEYINPUT115), .A3(new_n493), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT115), .B1(new_n834), .B2(new_n493), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n862), .A2(KEYINPUT116), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n862), .A2(KEYINPUT116), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n725), .A2(new_n601), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n841), .A2(new_n865), .ZN(new_n866));
  XOR2_X1   g680(.A(new_n866), .B(KEYINPUT48), .Z(new_n867));
  NOR3_X1   g681(.A1(new_n863), .A2(new_n864), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n856), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n848), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n832), .B1(new_n851), .B2(new_n852), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT114), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n872), .B(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n869), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT112), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n876), .B(KEYINPUT54), .C1(new_n828), .C2(new_n829), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n800), .B(KEYINPUT53), .C1(new_n813), .C2(new_n819), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n732), .A2(new_n799), .ZN(new_n880));
  INV_X1    g694(.A(new_n790), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n882), .B1(new_n825), .B2(new_n824), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n878), .B(new_n879), .C1(new_n883), .C2(KEYINPUT53), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n831), .A2(new_n875), .A3(new_n877), .A4(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT117), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n884), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n888), .B1(new_n830), .B2(KEYINPUT112), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n889), .A2(KEYINPUT117), .A3(new_n877), .A4(new_n875), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n857), .A2(new_n260), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n782), .B1(new_n887), .B2(new_n892), .ZN(G75));
  NOR2_X1   g707(.A1(new_n260), .A2(G952), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n879), .B1(new_n883), .B2(KEYINPUT53), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n896), .A2(G902), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT56), .B1(new_n897), .B2(G210), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n460), .A2(new_n471), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT118), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT55), .Z(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(new_n469), .Z(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n895), .B1(new_n898), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n897), .A2(G210), .ZN(new_n905));
  OR2_X1    g719(.A1(new_n903), .A2(KEYINPUT120), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n903), .A2(KEYINPUT120), .ZN(new_n907));
  XNOR2_X1  g721(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n905), .A2(new_n906), .A3(new_n907), .A4(new_n908), .ZN(new_n909));
  OR2_X1    g723(.A1(new_n909), .A2(KEYINPUT121), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(KEYINPUT121), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n904), .B1(new_n910), .B2(new_n911), .ZN(G51));
  XNOR2_X1  g726(.A(new_n896), .B(new_n878), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n432), .B(KEYINPUT57), .Z(new_n914));
  OAI22_X1  g728(.A1(new_n913), .A2(new_n914), .B1(new_n430), .B2(new_n428), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n897), .A2(new_n758), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n894), .B1(new_n915), .B2(new_n916), .ZN(G54));
  NAND3_X1  g731(.A1(new_n897), .A2(KEYINPUT58), .A3(G475), .ZN(new_n918));
  INV_X1    g732(.A(new_n253), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n918), .A2(new_n919), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n920), .A2(new_n921), .A3(new_n894), .ZN(G60));
  AND2_X1   g736(.A1(new_n614), .A2(new_n616), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n619), .B(KEYINPUT59), .Z(new_n924));
  OR2_X1    g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n895), .B1(new_n913), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n889), .A2(new_n877), .ZN(new_n927));
  INV_X1    g741(.A(new_n924), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n926), .B1(new_n929), .B2(new_n923), .ZN(G63));
  NAND2_X1  g744(.A1(G217), .A2(G902), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT122), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT60), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n896), .A2(new_n636), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n895), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n896), .A2(new_n933), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n599), .B(KEYINPUT123), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n938), .B1(KEYINPUT124), .B2(KEYINPUT61), .ZN(new_n939));
  XOR2_X1   g753(.A(KEYINPUT124), .B(KEYINPUT61), .Z(new_n940));
  OAI21_X1  g754(.A(new_n939), .B1(new_n938), .B2(new_n940), .ZN(G66));
  NAND2_X1  g755(.A1(G224), .A2(G953), .ZN(new_n942));
  OAI22_X1  g756(.A1(new_n790), .A2(G953), .B1(new_n263), .B2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(G898), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n900), .B1(new_n944), .B2(G953), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n943), .B(new_n945), .ZN(G69));
  AND2_X1   g760(.A1(new_n730), .A2(new_n731), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n769), .B1(new_n721), .B2(new_n947), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n805), .B(new_n865), .C1(new_n767), .C2(new_n768), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n684), .A2(new_n814), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n949), .A2(new_n741), .A3(new_n776), .A4(new_n950), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n948), .A2(new_n951), .A3(G953), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n529), .B(new_n953), .Z(new_n954));
  INV_X1    g768(.A(G900), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n954), .B1(new_n955), .B2(new_n260), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n952), .A2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n950), .A2(new_n676), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT62), .Z(new_n960));
  NOR3_X1   g774(.A1(new_n660), .A2(new_n743), .A3(new_n785), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n961), .B1(new_n602), .B2(new_n605), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n960), .A2(new_n769), .A3(new_n776), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n260), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n954), .B(KEYINPUT125), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(G953), .B1(new_n316), .B2(new_n955), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT126), .ZN(new_n968));
  OR2_X1    g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n958), .A2(new_n966), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n967), .A2(new_n968), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(G72));
  NAND2_X1  g786(.A1(G472), .A2(G902), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT63), .Z(new_n974));
  OAI21_X1  g788(.A(new_n974), .B1(new_n963), .B2(new_n790), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n530), .A2(new_n541), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n894), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n974), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n948), .A2(new_n951), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n978), .B1(new_n979), .B2(new_n881), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n530), .A2(new_n541), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT127), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n977), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  OR2_X1    g797(.A1(new_n828), .A2(new_n829), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n552), .A2(new_n554), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n978), .B1(new_n985), .B2(new_n665), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n983), .B1(new_n984), .B2(new_n986), .ZN(G57));
endmodule


