//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 0 0 0 0 0 0 0 1 1 0 0 0 1 1 0 1 0 1 0 0 0 1 0 0 1 0 1 1 1 0 0 0 0 0 0 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n809, new_n811, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n202));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT24), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT66), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G183gat), .B2(G190gat), .ZN(new_n206));
  INV_X1    g005(.A(G183gat), .ZN(new_n207));
  INV_X1    g006(.A(G190gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n207), .A2(new_n208), .A3(KEYINPUT66), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n204), .A2(new_n206), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  INV_X1    g010(.A(G169gat), .ZN(new_n212));
  INV_X1    g011(.A(G176gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n212), .A2(new_n213), .A3(KEYINPUT23), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n215), .B1(G169gat), .B2(G176gat), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n210), .A2(new_n211), .A3(new_n214), .A4(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT64), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(G183gat), .B2(G190gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n207), .A2(new_n208), .A3(KEYINPUT64), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(G169gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n222), .A2(KEYINPUT23), .A3(new_n213), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT25), .B1(G169gat), .B2(G176gat), .ZN(new_n224));
  AND3_X1   g023(.A1(new_n223), .A2(new_n216), .A3(new_n224), .ZN(new_n225));
  AOI22_X1  g024(.A1(new_n217), .A2(KEYINPUT25), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n207), .A2(KEYINPUT27), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n227), .A2(KEYINPUT67), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n207), .A2(KEYINPUT27), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(KEYINPUT67), .ZN(new_n230));
  NOR2_X1   g029(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n228), .A2(new_n229), .A3(new_n230), .A4(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n227), .A2(new_n229), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT28), .B1(new_n233), .B2(G190gat), .ZN(new_n234));
  AND3_X1   g033(.A1(new_n212), .A2(new_n213), .A3(KEYINPUT26), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT26), .B1(new_n212), .B2(new_n213), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n211), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n232), .A2(new_n203), .A3(new_n234), .A4(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n226), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(G127gat), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT68), .B1(new_n240), .B2(G134gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(G134gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(G134gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G127gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n245), .A2(KEYINPUT68), .ZN(new_n246));
  XNOR2_X1  g045(.A(G113gat), .B(G120gat), .ZN(new_n247));
  OAI22_X1  g046(.A1(new_n243), .A2(new_n246), .B1(new_n247), .B2(KEYINPUT1), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(KEYINPUT69), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n245), .A2(new_n242), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT70), .B(KEYINPUT1), .ZN(new_n251));
  OR3_X1    g050(.A1(new_n247), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n239), .A2(new_n253), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n226), .A2(new_n249), .A3(new_n252), .A4(new_n238), .ZN(new_n255));
  AND2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(G227gat), .ZN(new_n257));
  INV_X1    g056(.A(G233gat), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(KEYINPUT32), .B1(new_n256), .B2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G15gat), .B(G43gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(G71gat), .B(G99gat), .ZN(new_n263));
  XOR2_X1   g062(.A(new_n262), .B(new_n263), .Z(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT33), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n202), .B1(new_n261), .B2(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n260), .B1(new_n254), .B2(new_n255), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT32), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n270), .A2(KEYINPUT72), .A3(new_n265), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n254), .A2(new_n260), .A3(new_n255), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(KEYINPUT34), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT73), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n276));
  OR3_X1    g075(.A1(new_n268), .A2(new_n276), .A3(KEYINPUT33), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n276), .B1(new_n268), .B2(KEYINPUT33), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n277), .A2(new_n261), .A3(new_n278), .A4(new_n264), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n272), .A2(new_n275), .A3(new_n279), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n274), .A2(KEYINPUT73), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n281), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n283), .A2(new_n272), .A3(new_n275), .A4(new_n279), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n282), .A2(KEYINPUT36), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT36), .B1(new_n282), .B2(new_n284), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT30), .ZN(new_n289));
  XNOR2_X1  g088(.A(G8gat), .B(G36gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(G64gat), .B(G92gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT22), .ZN(new_n293));
  INV_X1    g092(.A(G211gat), .ZN(new_n294));
  INV_X1    g093(.A(G218gat), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G197gat), .ZN(new_n297));
  INV_X1    g096(.A(G204gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g098(.A1(G197gat), .A2(G204gat), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n296), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n301), .A2(KEYINPUT74), .ZN(new_n302));
  XNOR2_X1  g101(.A(G211gat), .B(G218gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G226gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n305), .A2(new_n258), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  OR2_X1    g106(.A1(new_n239), .A2(KEYINPUT75), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n239), .A2(KEYINPUT75), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n239), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n306), .A2(KEYINPUT29), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n304), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n311), .A2(new_n306), .ZN(new_n316));
  INV_X1    g115(.A(new_n304), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n308), .A2(new_n309), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n316), .B(new_n317), .C1(new_n318), .C2(new_n313), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n292), .B1(new_n315), .B2(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n320), .A2(KEYINPUT76), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT76), .ZN(new_n322));
  AOI211_X1 g121(.A(new_n322), .B(new_n292), .C1(new_n315), .C2(new_n319), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n289), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n315), .A2(new_n319), .ZN(new_n325));
  INV_X1    g124(.A(new_n292), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n327), .B1(KEYINPUT30), .B2(new_n320), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT81), .ZN(new_n330));
  XOR2_X1   g129(.A(G155gat), .B(G162gat), .Z(new_n331));
  INV_X1    g130(.A(KEYINPUT77), .ZN(new_n332));
  XOR2_X1   g131(.A(G141gat), .B(G148gat), .Z(new_n333));
  AOI21_X1  g132(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G155gat), .ZN(new_n335));
  INV_X1    g134(.A(G162gat), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT2), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  XOR2_X1   g137(.A(new_n334), .B(new_n338), .Z(new_n339));
  NOR2_X1   g138(.A1(new_n253), .A2(new_n339), .ZN(new_n340));
  XOR2_X1   g139(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT79), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT79), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n340), .A2(new_n344), .A3(new_n341), .ZN(new_n345));
  OAI21_X1  g144(.A(KEYINPUT4), .B1(new_n253), .B2(new_n339), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n343), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n339), .A2(KEYINPUT3), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n334), .B(new_n338), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT3), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n348), .A2(new_n253), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(G225gat), .A2(G233gat), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n354), .A2(KEYINPUT5), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n347), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n340), .A2(KEYINPUT4), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n341), .B1(new_n253), .B2(new_n339), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n357), .A2(new_n352), .A3(new_n358), .A4(new_n353), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n253), .B(new_n339), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(new_n354), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n359), .A2(new_n361), .A3(KEYINPUT5), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n356), .A2(new_n362), .ZN(new_n363));
  XOR2_X1   g162(.A(G1gat), .B(G29gat), .Z(new_n364));
  XNOR2_X1  g163(.A(new_n364), .B(G85gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT0), .B(G57gat), .ZN(new_n366));
  XOR2_X1   g165(.A(new_n365), .B(new_n366), .Z(new_n367));
  NAND2_X1  g166(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT6), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n330), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n367), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n371), .B1(new_n356), .B2(new_n362), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n372), .A2(KEYINPUT81), .A3(KEYINPUT6), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT80), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n372), .A2(KEYINPUT6), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n356), .A2(new_n371), .A3(new_n362), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n376), .A2(new_n375), .A3(new_n377), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n329), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT29), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n351), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n304), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n350), .B1(new_n304), .B2(KEYINPUT29), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(new_n339), .ZN(new_n386));
  AND2_X1   g185(.A1(G228gat), .A2(G233gat), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n384), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  OR2_X1    g188(.A1(new_n301), .A2(new_n303), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT29), .B1(new_n301), .B2(new_n303), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT3), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n349), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n393), .B1(new_n383), .B2(new_n304), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n394), .A2(new_n387), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n389), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT84), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(G22gat), .ZN(new_n398));
  OR2_X1    g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(G50gat), .ZN(new_n401));
  XOR2_X1   g200(.A(G78gat), .B(G106gat), .Z(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n403), .B1(new_n396), .B2(new_n398), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n399), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT85), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n399), .A2(KEYINPUT85), .A3(new_n404), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(G22gat), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n396), .A2(new_n410), .ZN(new_n411));
  NOR3_X1   g210(.A1(new_n389), .A2(new_n395), .A3(G22gat), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n403), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT83), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OAI211_X1 g214(.A(KEYINPUT83), .B(new_n403), .C1(new_n411), .C2(new_n412), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n409), .A2(new_n417), .ZN(new_n418));
  OAI211_X1 g217(.A(KEYINPUT86), .B(new_n288), .C1(new_n381), .C2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT86), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n372), .A2(KEYINPUT81), .A3(KEYINPUT6), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT81), .B1(new_n372), .B2(KEYINPUT6), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n368), .A2(new_n369), .A3(new_n377), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT80), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n423), .A2(new_n380), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n329), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n418), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n287), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n285), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n420), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n353), .B1(new_n347), .B2(new_n352), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT39), .B1(new_n360), .B2(new_n354), .ZN(new_n433));
  OR2_X1    g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT39), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n367), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT87), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n436), .A2(new_n437), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n434), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT40), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n372), .B1(new_n324), .B2(new_n328), .ZN(new_n443));
  OAI211_X1 g242(.A(KEYINPUT40), .B(new_n434), .C1(new_n438), .C2(new_n439), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n423), .A2(KEYINPUT89), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT89), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n374), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n446), .A2(new_n448), .A3(new_n424), .ZN(new_n449));
  OR2_X1    g248(.A1(new_n310), .A2(new_n314), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT88), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n450), .A2(new_n451), .A3(new_n317), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n316), .B1(new_n318), .B2(new_n313), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n452), .B1(new_n317), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n451), .B1(new_n450), .B2(new_n317), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT37), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT38), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT37), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n326), .B1(new_n325), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n456), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  OR2_X1    g259(.A1(new_n321), .A2(new_n323), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n459), .B1(new_n458), .B2(new_n325), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT38), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n460), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n445), .B(new_n418), .C1(new_n449), .C2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n419), .A2(new_n431), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n282), .A2(new_n284), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n329), .A2(KEYINPUT35), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n449), .A2(new_n467), .A3(new_n418), .A4(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n426), .A2(new_n427), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n418), .A2(new_n467), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT35), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n466), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(G113gat), .B(G141gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n475), .B(new_n297), .ZN(new_n476));
  XNOR2_X1  g275(.A(KEYINPUT11), .B(G169gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n476), .B(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n478), .B(KEYINPUT12), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(G8gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(G15gat), .B(G22gat), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT16), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n482), .B1(new_n483), .B2(G1gat), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n481), .B1(new_n484), .B2(KEYINPUT91), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n484), .B1(G1gat), .B2(new_n482), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n485), .B(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT14), .ZN(new_n488));
  INV_X1    g287(.A(G29gat), .ZN(new_n489));
  INV_X1    g288(.A(G36gat), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n493), .B1(new_n489), .B2(new_n490), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT15), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n491), .A2(new_n492), .B1(G29gat), .B2(G36gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT15), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(G43gat), .B(G50gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n500), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(KEYINPUT90), .A2(KEYINPUT17), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT90), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT17), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n501), .A2(new_n503), .A3(new_n504), .A4(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n502), .B1(new_n496), .B2(new_n498), .ZN(new_n509));
  INV_X1    g308(.A(new_n503), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n505), .B(new_n506), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n487), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n509), .A2(new_n510), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(new_n487), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(G229gat), .A2(G233gat), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  NOR3_X1   g316(.A1(new_n512), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT18), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n487), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n501), .A2(new_n503), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(new_n514), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n516), .B(KEYINPUT13), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n527), .B1(new_n518), .B2(KEYINPUT18), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n480), .B1(new_n520), .B2(new_n528), .ZN(new_n529));
  OR2_X1    g328(.A1(new_n518), .A2(KEYINPUT18), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n530), .A2(new_n519), .A3(new_n527), .A4(new_n479), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G230gat), .A2(G233gat), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G57gat), .B(G64gat), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(G71gat), .ZN(new_n538));
  INV_X1    g337(.A(G78gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G71gat), .A2(G78gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT9), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n537), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n541), .B(new_n540), .C1(new_n536), .C2(new_n543), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G99gat), .B(G106gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(G85gat), .A2(G92gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(KEYINPUT92), .A2(KEYINPUT7), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g350(.A1(KEYINPUT92), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n552));
  OR2_X1    g351(.A1(G85gat), .A2(G92gat), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(KEYINPUT93), .B1(G99gat), .B2(G106gat), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(KEYINPUT93), .A2(G99gat), .A3(G106gat), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n557), .A2(KEYINPUT8), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n548), .B1(new_n555), .B2(new_n559), .ZN(new_n560));
  AND3_X1   g359(.A1(KEYINPUT93), .A2(G99gat), .A3(G106gat), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT8), .ZN(new_n562));
  NOR3_X1   g361(.A1(new_n561), .A2(new_n556), .A3(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(G99gat), .B(G106gat), .Z(new_n564));
  NOR3_X1   g363(.A1(new_n563), .A2(new_n554), .A3(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n547), .B1(new_n560), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT10), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n564), .B1(new_n563), .B2(new_n554), .ZN(new_n568));
  NOR2_X1   g367(.A1(G85gat), .A2(G92gat), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n569), .B1(new_n549), .B2(new_n550), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n559), .A2(new_n548), .A3(new_n552), .A4(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n568), .A2(new_n571), .A3(new_n546), .A4(new_n545), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n566), .A2(new_n567), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT94), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n574), .B1(new_n560), .B2(new_n565), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n568), .A2(new_n571), .A3(KEYINPUT94), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n547), .A2(new_n567), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n535), .B1(new_n573), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT95), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n566), .A2(new_n572), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n580), .B1(new_n581), .B2(new_n535), .ZN(new_n582));
  AOI211_X1 g381(.A(KEYINPUT95), .B(new_n534), .C1(new_n566), .C2(new_n572), .ZN(new_n583));
  NOR3_X1   g382(.A1(new_n579), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G120gat), .B(G148gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(G176gat), .B(G204gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n584), .A2(KEYINPUT96), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT96), .B1(new_n584), .B2(new_n588), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n584), .A2(new_n588), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n533), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT21), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n547), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n547), .A2(new_n596), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n521), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n600), .B1(new_n521), .B2(new_n599), .ZN(new_n601));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(new_n207), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(G211gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n601), .B(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(G127gat), .B(G155gat), .Z(new_n606));
  XOR2_X1   g405(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n605), .B(new_n608), .Z(new_n609));
  NAND2_X1  g408(.A1(new_n508), .A2(new_n511), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n575), .A2(new_n576), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(G134gat), .B(G162gat), .Z(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  AND2_X1   g413(.A1(G232gat), .A2(G233gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(KEYINPUT41), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n616), .B1(new_n522), .B2(new_n611), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n612), .A2(new_n614), .A3(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n611), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n620), .B1(new_n508), .B2(new_n511), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n613), .B1(new_n621), .B2(new_n617), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n615), .A2(KEYINPUT41), .ZN(new_n623));
  XNOR2_X1  g422(.A(G190gat), .B(G218gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  AND3_X1   g424(.A1(new_n619), .A2(new_n622), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n625), .B1(new_n619), .B2(new_n622), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n609), .A2(new_n628), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n474), .A2(new_n595), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n426), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g432(.A1(new_n630), .A2(new_n329), .ZN(new_n634));
  OAI21_X1  g433(.A(KEYINPUT42), .B1(new_n634), .B2(new_n481), .ZN(new_n635));
  XOR2_X1   g434(.A(KEYINPUT16), .B(G8gat), .Z(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  MUX2_X1   g436(.A(KEYINPUT42), .B(new_n635), .S(new_n637), .Z(G1325gat));
  NAND2_X1  g437(.A1(new_n630), .A2(new_n430), .ZN(new_n639));
  AOI21_X1  g438(.A(G15gat), .B1(new_n282), .B2(new_n284), .ZN(new_n640));
  AOI22_X1  g439(.A1(new_n639), .A2(G15gat), .B1(new_n630), .B2(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n641), .B(KEYINPUT97), .Z(G1326gat));
  INV_X1    g441(.A(new_n418), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n630), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT43), .B(G22gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(G1327gat));
  NAND2_X1  g445(.A1(new_n474), .A2(new_n628), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n595), .A2(new_n609), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n649), .A2(new_n489), .A3(new_n631), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT45), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT44), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n652), .B1(new_n474), .B2(new_n628), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n428), .A2(new_n430), .ZN(new_n654));
  AOI22_X1  g453(.A1(new_n465), .A2(new_n654), .B1(new_n469), .B2(new_n472), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n628), .A2(KEYINPUT98), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n628), .A2(KEYINPUT98), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NOR3_X1   g457(.A1(new_n655), .A2(KEYINPUT44), .A3(new_n658), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n653), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n648), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(G29gat), .B1(new_n662), .B2(new_n426), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n651), .A2(new_n663), .ZN(G1328gat));
  NAND3_X1  g463(.A1(new_n649), .A2(new_n490), .A3(new_n329), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(KEYINPUT46), .Z(new_n666));
  OAI21_X1  g465(.A(G36gat), .B1(new_n662), .B2(new_n427), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(G1329gat));
  OAI211_X1 g467(.A(new_n430), .B(new_n661), .C1(new_n653), .C2(new_n659), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(G43gat), .ZN(new_n670));
  INV_X1    g469(.A(G43gat), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n649), .A2(new_n671), .A3(new_n467), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT47), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n670), .A2(KEYINPUT47), .A3(new_n672), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(G1330gat));
  OAI211_X1 g476(.A(new_n643), .B(new_n661), .C1(new_n653), .C2(new_n659), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(G50gat), .ZN(new_n679));
  INV_X1    g478(.A(G50gat), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n643), .A2(new_n680), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n647), .A2(new_n648), .A3(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT99), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT48), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT100), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n686), .B1(new_n683), .B2(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n682), .B1(new_n678), .B2(G50gat), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n689), .B1(new_n690), .B2(new_n688), .ZN(new_n691));
  OAI21_X1  g490(.A(KEYINPUT99), .B1(new_n690), .B2(KEYINPUT48), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n687), .A2(new_n691), .A3(new_n692), .ZN(G1331gat));
  NOR2_X1   g492(.A1(new_n655), .A2(new_n532), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n694), .A2(new_n594), .A3(new_n629), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n695), .A2(new_n426), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT101), .B(G57gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1332gat));
  NOR2_X1   g497(.A1(new_n695), .A2(new_n427), .ZN(new_n699));
  NOR2_X1   g498(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n700));
  AND2_X1   g499(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n699), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n702), .B1(new_n699), .B2(new_n700), .ZN(G1333gat));
  OAI21_X1  g502(.A(G71gat), .B1(new_n695), .B2(new_n288), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n467), .A2(new_n538), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n704), .B1(new_n695), .B2(new_n705), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g506(.A1(new_n695), .A2(new_n418), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(new_n539), .ZN(G1335gat));
  INV_X1    g508(.A(KEYINPUT51), .ZN(new_n710));
  INV_X1    g509(.A(new_n609), .ZN(new_n711));
  INV_X1    g510(.A(new_n628), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n710), .B1(new_n694), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n465), .A2(new_n654), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n473), .ZN(new_n716));
  AND4_X1   g515(.A1(new_n710), .A2(new_n716), .A3(new_n533), .A4(new_n713), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n594), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n426), .A2(G85gat), .A3(new_n719), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT103), .Z(new_n721));
  NAND2_X1  g520(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n711), .A2(new_n532), .A3(new_n719), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n660), .A2(new_n631), .A3(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT102), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(G85gat), .B1(new_n724), .B2(new_n725), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n722), .B1(new_n726), .B2(new_n727), .ZN(G1336gat));
  NAND3_X1  g527(.A1(new_n716), .A2(new_n533), .A3(new_n713), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(KEYINPUT104), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n714), .B2(new_n717), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n729), .A2(KEYINPUT104), .A3(new_n710), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n427), .A2(G92gat), .A3(new_n719), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n329), .B(new_n723), .C1(new_n653), .C2(new_n659), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(G92gat), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(KEYINPUT52), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT52), .B1(new_n718), .B2(new_n733), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n736), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n740), .ZN(G1337gat));
  NAND3_X1  g540(.A1(new_n660), .A2(new_n430), .A3(new_n723), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(G99gat), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n719), .A2(G99gat), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n718), .A2(new_n467), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(G1338gat));
  NOR3_X1   g545(.A1(new_n418), .A2(G106gat), .A3(new_n719), .ZN(new_n747));
  XOR2_X1   g546(.A(new_n747), .B(KEYINPUT105), .Z(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT106), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n731), .A2(new_n732), .A3(new_n749), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n643), .B(new_n723), .C1(new_n653), .C2(new_n659), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G106gat), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(KEYINPUT53), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n718), .A2(new_n748), .ZN(new_n755));
  XNOR2_X1  g554(.A(KEYINPUT107), .B(KEYINPUT53), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n752), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n754), .A2(new_n757), .ZN(G1339gat));
  INV_X1    g557(.A(KEYINPUT54), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n588), .B1(new_n579), .B2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  AND3_X1   g560(.A1(new_n573), .A2(new_n578), .A3(new_n535), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n573), .A2(new_n578), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n534), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT108), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n762), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n573), .A2(new_n578), .A3(new_n535), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT54), .B1(new_n767), .B2(KEYINPUT108), .ZN(new_n768));
  OAI21_X1  g567(.A(KEYINPUT109), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n759), .B1(new_n762), .B2(new_n765), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT109), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n767), .B1(new_n579), .B2(KEYINPUT108), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n761), .B1(new_n769), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(KEYINPUT110), .B1(new_n774), .B2(KEYINPUT55), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n591), .B1(new_n774), .B2(KEYINPUT55), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n771), .B1(new_n770), .B2(new_n772), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n760), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT110), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n775), .A2(new_n776), .A3(new_n532), .A4(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT111), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n512), .A2(new_n515), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n784), .B1(new_n785), .B2(new_n516), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n523), .A2(new_n514), .A3(new_n525), .ZN(new_n787));
  OAI211_X1 g586(.A(KEYINPUT111), .B(new_n517), .C1(new_n512), .C2(new_n515), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n478), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n790), .A2(new_n531), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n594), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n783), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT112), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n783), .A2(KEYINPUT112), .A3(new_n792), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n795), .A2(new_n658), .A3(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n791), .A2(new_n775), .A3(new_n776), .A4(new_n782), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n798), .A2(new_n658), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n711), .B1(new_n797), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n629), .A2(new_n533), .A3(new_n719), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n631), .A2(new_n427), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n804), .A2(new_n471), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n532), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n594), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g609(.A1(new_n806), .A2(new_n711), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g611(.A1(new_n806), .A2(new_n628), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n813), .A2(G134gat), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(KEYINPUT56), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n813), .A2(G134gat), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(KEYINPUT113), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(G1343gat));
  INV_X1    g617(.A(new_n658), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n819), .B1(new_n793), .B2(new_n794), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n799), .B1(new_n820), .B2(new_n796), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n802), .B1(new_n821), .B2(new_n711), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n805), .A2(new_n430), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n533), .A2(G141gat), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n822), .A2(new_n823), .A3(new_n643), .A4(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT58), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(KEYINPUT57), .B1(new_n822), .B2(new_n643), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n643), .A2(KEYINPUT57), .ZN(new_n829));
  OAI21_X1  g628(.A(KEYINPUT114), .B1(new_n774), .B2(KEYINPUT55), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT114), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n779), .A2(new_n831), .A3(new_n781), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n830), .A2(new_n776), .A3(new_n532), .A4(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n628), .B1(new_n833), .B2(new_n792), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n609), .B1(new_n834), .B2(new_n799), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n835), .A2(KEYINPUT115), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n803), .B1(new_n835), .B2(KEYINPUT115), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n829), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n532), .B(new_n823), .C1(new_n828), .C2(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n827), .B1(new_n839), .B2(G141gat), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(KEYINPUT117), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n823), .B1(new_n828), .B2(new_n838), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(KEYINPUT116), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n844), .B(new_n823), .C1(new_n828), .C2(new_n838), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n532), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n804), .A2(new_n418), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n823), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  AOI22_X1  g649(.A1(new_n847), .A2(G141gat), .B1(new_n850), .B2(new_n824), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n841), .B1(new_n851), .B2(new_n826), .ZN(G1344gat));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n853));
  AOI211_X1 g652(.A(new_n853), .B(G148gat), .C1(new_n850), .C2(new_n594), .ZN(new_n854));
  OAI211_X1 g653(.A(KEYINPUT57), .B(new_n643), .C1(new_n801), .C2(new_n803), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(KEYINPUT119), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n822), .A2(new_n857), .A3(KEYINPUT57), .A4(new_n643), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n798), .A2(new_n712), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n609), .B1(new_n834), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n418), .B1(new_n860), .B2(new_n802), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n861), .A2(KEYINPUT57), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n856), .A2(new_n858), .A3(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n823), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT118), .ZN(new_n865));
  AOI211_X1 g664(.A(new_n853), .B(new_n719), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n863), .B(new_n866), .C1(new_n865), .C2(new_n864), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n719), .B1(new_n843), .B2(new_n845), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n867), .B1(new_n868), .B2(KEYINPUT59), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n854), .B1(new_n869), .B2(G148gat), .ZN(G1345gat));
  AOI21_X1  g669(.A(G155gat), .B1(new_n850), .B2(new_n711), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n609), .A2(new_n335), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n871), .B1(new_n846), .B2(new_n872), .ZN(G1346gat));
  NAND3_X1  g672(.A1(new_n850), .A2(new_n336), .A3(new_n628), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n658), .B1(new_n843), .B2(new_n845), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n874), .B1(new_n875), .B2(new_n336), .ZN(G1347gat));
  NOR3_X1   g675(.A1(new_n631), .A2(new_n471), .A3(new_n427), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n822), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n532), .ZN(new_n879));
  MUX2_X1   g678(.A(new_n222), .B(G169gat), .S(new_n879), .Z(G1348gat));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n594), .ZN(new_n881));
  XNOR2_X1  g680(.A(KEYINPUT120), .B(G176gat), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n881), .B(new_n882), .ZN(G1349gat));
  NAND2_X1  g682(.A1(new_n878), .A2(new_n711), .ZN(new_n884));
  OR3_X1    g683(.A1(new_n884), .A2(KEYINPUT121), .A3(new_n233), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n884), .A2(new_n233), .ZN(new_n886));
  AOI21_X1  g685(.A(KEYINPUT121), .B1(new_n884), .B2(G183gat), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g688(.A1(new_n878), .A2(new_n208), .A3(new_n819), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n878), .A2(new_n628), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(G190gat), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n892), .A2(KEYINPUT61), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n892), .A2(KEYINPUT61), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n890), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT122), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n895), .B(new_n896), .ZN(G1351gat));
  NOR3_X1   g696(.A1(new_n430), .A2(new_n631), .A3(new_n427), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n848), .A2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT123), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n848), .A2(KEYINPUT123), .A3(new_n898), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g702(.A(KEYINPUT124), .B(G197gat), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n903), .A2(new_n532), .A3(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n863), .ZN(new_n907));
  XOR2_X1   g706(.A(new_n898), .B(KEYINPUT125), .Z(new_n908));
  NOR3_X1   g707(.A1(new_n907), .A2(new_n533), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n906), .B1(new_n909), .B2(new_n905), .ZN(G1352gat));
  NOR3_X1   g709(.A1(new_n899), .A2(G204gat), .A3(new_n719), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT62), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n907), .A2(new_n719), .A3(new_n908), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n912), .B1(new_n298), .B2(new_n913), .ZN(G1353gat));
  NAND3_X1  g713(.A1(new_n903), .A2(new_n294), .A3(new_n711), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n898), .A2(new_n711), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n863), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(KEYINPUT63), .B1(new_n917), .B2(G211gat), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT63), .ZN(new_n919));
  AOI211_X1 g718(.A(new_n919), .B(new_n294), .C1(new_n863), .C2(new_n916), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n915), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(KEYINPUT126), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT126), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n915), .B(new_n923), .C1(new_n918), .C2(new_n920), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(G1354gat));
  OAI21_X1  g724(.A(KEYINPUT127), .B1(new_n907), .B2(new_n908), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(new_n628), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n907), .A2(KEYINPUT127), .A3(new_n908), .ZN(new_n928));
  OAI21_X1  g727(.A(G218gat), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n903), .A2(new_n295), .A3(new_n819), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1355gat));
endmodule


