//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 0 0 1 0 0 0 1 0 0 1 1 0 0 1 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1223, new_n1224,
    new_n1225, new_n1227, new_n1228, new_n1229, new_n1230, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(new_n204));
  INV_X1    g0004(.A(G50), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n209));
  INV_X1    g0009(.A(G116), .ZN(new_n210));
  INV_X1    g0010(.A(G270), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  INV_X1    g0014(.A(G97), .ZN(new_n215));
  INV_X1    g0015(.A(G257), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n213), .B1(new_n202), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI211_X1 g0017(.A(new_n212), .B(new_n217), .C1(G58), .C2(G232), .ZN(new_n218));
  INV_X1    g0018(.A(G1), .ZN(new_n219));
  INV_X1    g0019(.A(G20), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT1), .Z(new_n223));
  NAND2_X1  g0023(.A1(new_n203), .A2(G50), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  NOR3_X1   g0025(.A1(new_n224), .A2(new_n220), .A3(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(G250), .ZN(new_n227));
  INV_X1    g0027(.A(G13), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n221), .A2(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(G264), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n227), .B(new_n229), .C1(new_n216), .C2(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT0), .ZN(new_n232));
  NOR3_X1   g0032(.A1(new_n223), .A2(new_n226), .A3(new_n232), .ZN(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G264), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(new_n211), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G107), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n210), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  NAND2_X1  g0048(.A1(new_n220), .A2(G33), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  OR2_X1    g0050(.A1(KEYINPUT8), .A2(G58), .ZN(new_n251));
  NAND2_X1  g0051(.A1(KEYINPUT8), .A2(G58), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n251), .A2(KEYINPUT65), .A3(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(KEYINPUT65), .B1(new_n251), .B2(new_n252), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n250), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n220), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G150), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n220), .B1(new_n204), .B2(new_n205), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n256), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n225), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n219), .A2(G20), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(new_n228), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(G50), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n266), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n268), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(new_n205), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n267), .A2(new_n272), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT9), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n219), .B1(G41), .B2(G45), .ZN(new_n280));
  INV_X1    g0080(.A(G274), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT3), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n284), .A2(new_n285), .A3(G223), .A4(G1698), .ZN(new_n286));
  INV_X1    g0086(.A(G1698), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n284), .A2(new_n285), .A3(G222), .A4(new_n287), .ZN(new_n288));
  AND2_X1   g0088(.A1(new_n284), .A2(new_n285), .ZN(new_n289));
  INV_X1    g0089(.A(G77), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n286), .B(new_n288), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n225), .B1(G33), .B2(G41), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n282), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT64), .ZN(new_n294));
  INV_X1    g0094(.A(G41), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n294), .B1(new_n257), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n225), .ZN(new_n297));
  NAND3_X1  g0097(.A1(KEYINPUT64), .A2(G33), .A3(G41), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n299), .A2(new_n280), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G226), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n293), .A2(G190), .A3(new_n301), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n267), .A2(KEYINPUT9), .A3(new_n272), .A4(new_n276), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n293), .A2(new_n301), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G200), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n279), .A2(new_n302), .A3(new_n303), .A4(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT10), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n303), .A2(new_n305), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT10), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n308), .A2(new_n309), .A3(new_n302), .A4(new_n279), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n284), .A2(new_n285), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G107), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n284), .A2(new_n285), .A3(G238), .A4(G1698), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n284), .A2(new_n285), .A3(G232), .A4(new_n287), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT66), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT66), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n313), .A2(new_n318), .A3(new_n314), .A4(new_n315), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n317), .A2(new_n292), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n282), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n300), .A2(G244), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G169), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT15), .B(G87), .ZN(new_n326));
  OR3_X1    g0126(.A1(new_n326), .A2(KEYINPUT67), .A3(new_n249), .ZN(new_n327));
  NAND2_X1  g0127(.A1(G20), .A2(G77), .ZN(new_n328));
  OAI21_X1  g0128(.A(KEYINPUT67), .B1(new_n326), .B2(new_n249), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT8), .B(G58), .ZN(new_n330));
  OR2_X1    g0130(.A1(new_n330), .A2(new_n258), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n327), .A2(new_n328), .A3(new_n329), .A4(new_n331), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n332), .A2(new_n266), .B1(new_n290), .B2(new_n269), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(new_n290), .B2(new_n274), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n325), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT68), .ZN(new_n336));
  OR2_X1    g0136(.A1(new_n323), .A2(G179), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT68), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n325), .A2(new_n334), .A3(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n336), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n304), .A2(new_n324), .ZN(new_n341));
  INV_X1    g0141(.A(G179), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n293), .A2(new_n342), .A3(new_n301), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n277), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n323), .A2(G200), .ZN(new_n345));
  INV_X1    g0145(.A(G190), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n345), .B1(new_n346), .B2(new_n323), .ZN(new_n347));
  OR2_X1    g0147(.A1(new_n347), .A2(new_n334), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n311), .A2(new_n340), .A3(new_n344), .A4(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT69), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n340), .A2(new_n348), .ZN(new_n352));
  INV_X1    g0152(.A(new_n344), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n353), .B1(new_n307), .B2(new_n310), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n352), .A2(KEYINPUT69), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n284), .A2(new_n285), .A3(G226), .A4(new_n287), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n284), .A2(new_n285), .A3(G232), .A4(G1698), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G33), .A2(G97), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n282), .B1(new_n360), .B2(new_n292), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n300), .A2(G238), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT13), .ZN(new_n363));
  AND3_X1   g0163(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n363), .B1(new_n361), .B2(new_n362), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(KEYINPUT14), .B1(new_n366), .B2(new_n324), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT14), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n368), .B(G169), .C1(new_n364), .C2(new_n365), .ZN(new_n369));
  INV_X1    g0169(.A(new_n366), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n367), .B(new_n369), .C1(new_n342), .C2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n202), .A2(G20), .ZN(new_n372));
  NOR3_X1   g0172(.A1(new_n372), .A2(G1), .A3(new_n228), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n373), .A2(KEYINPUT12), .ZN(new_n374));
  OAI221_X1 g0174(.A(new_n372), .B1(new_n249), .B2(new_n290), .C1(new_n205), .C2(new_n258), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n375), .A2(new_n266), .ZN(new_n376));
  XOR2_X1   g0176(.A(KEYINPUT70), .B(KEYINPUT11), .Z(new_n377));
  AND2_X1   g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n376), .A2(new_n377), .ZN(new_n379));
  OAI22_X1  g0179(.A1(new_n274), .A2(new_n202), .B1(KEYINPUT12), .B2(new_n373), .ZN(new_n380));
  OR4_X1    g0180(.A1(new_n374), .A2(new_n378), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n371), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n381), .B1(new_n370), .B2(G200), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n366), .A2(G190), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT71), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT71), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n382), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G58), .A2(G68), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n220), .B1(new_n203), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT74), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(G159), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n258), .A2(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n392), .A2(new_n393), .ZN(new_n398));
  NOR3_X1   g0198(.A1(new_n395), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  AND2_X1   g0199(.A1(KEYINPUT72), .A2(G33), .ZN(new_n400));
  NOR2_X1   g0200(.A1(KEYINPUT72), .A2(G33), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT3), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n284), .A2(KEYINPUT73), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  OAI211_X1 g0204(.A(KEYINPUT73), .B(KEYINPUT3), .C1(new_n400), .C2(new_n401), .ZN(new_n405));
  AOI21_X1  g0205(.A(G20), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT7), .ZN(new_n407));
  OAI21_X1  g0207(.A(G68), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  AOI211_X1 g0208(.A(KEYINPUT7), .B(G20), .C1(new_n404), .C2(new_n405), .ZN(new_n409));
  OAI211_X1 g0209(.A(KEYINPUT16), .B(new_n399), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT75), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT72), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n257), .ZN(new_n414));
  NAND2_X1  g0214(.A1(KEYINPUT72), .A2(G33), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n285), .B1(new_n416), .B2(KEYINPUT3), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n417), .A2(KEYINPUT7), .A3(new_n220), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n407), .B1(new_n289), .B2(G20), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n399), .B1(new_n420), .B2(new_n202), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT16), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n283), .B1(new_n414), .B2(new_n415), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT73), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(new_n283), .B2(G33), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n405), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n220), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT7), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n406), .A2(new_n407), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(new_n430), .A3(G68), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n431), .A2(KEYINPUT75), .A3(KEYINPUT16), .A4(new_n399), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n412), .A2(new_n423), .A3(new_n432), .A4(new_n266), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT65), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n330), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n253), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n436), .A2(new_n270), .ZN(new_n437));
  INV_X1    g0237(.A(new_n274), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n437), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  XOR2_X1   g0239(.A(new_n439), .B(KEYINPUT76), .Z(new_n440));
  NAND2_X1  g0240(.A1(new_n300), .A2(G232), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n426), .B1(new_n416), .B2(KEYINPUT3), .ZN(new_n443));
  INV_X1    g0243(.A(new_n405), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT77), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n445), .A2(new_n446), .A3(G223), .A4(new_n287), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n405), .B(new_n287), .C1(new_n424), .C2(new_n426), .ZN(new_n448));
  INV_X1    g0248(.A(G223), .ZN(new_n449));
  OAI21_X1  g0249(.A(KEYINPUT77), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n404), .A2(G226), .A3(G1698), .A4(new_n405), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G33), .A2(G87), .ZN(new_n452));
  XNOR2_X1  g0252(.A(new_n452), .B(KEYINPUT78), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n447), .A2(new_n450), .A3(new_n451), .A4(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n442), .B1(new_n454), .B2(new_n292), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n455), .A2(new_n346), .A3(new_n321), .ZN(new_n456));
  AOI21_X1  g0256(.A(G200), .B1(new_n455), .B2(new_n321), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n433), .B(new_n440), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT17), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n433), .A2(new_n440), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT17), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n455), .A2(new_n346), .A3(new_n321), .ZN(new_n462));
  AOI211_X1 g0262(.A(new_n282), .B(new_n442), .C1(new_n454), .C2(new_n292), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n462), .B1(new_n463), .B2(G200), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n460), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n454), .A2(new_n292), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n466), .A2(G179), .A3(new_n321), .A4(new_n441), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(new_n463), .B2(new_n324), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n433), .A2(new_n440), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT18), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n468), .A2(new_n469), .A3(KEYINPUT18), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n459), .A2(new_n465), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n356), .A2(new_n390), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT79), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n356), .A2(new_n390), .A3(new_n474), .A4(KEYINPUT79), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  XOR2_X1   g0279(.A(KEYINPUT80), .B(KEYINPUT4), .Z(new_n480));
  INV_X1    g0280(.A(G244), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n480), .B1(new_n448), .B2(new_n481), .ZN(new_n482));
  AND2_X1   g0282(.A1(KEYINPUT4), .A2(G244), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n289), .A2(new_n287), .A3(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n284), .A2(new_n285), .A3(G250), .A4(G1698), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G283), .ZN(new_n486));
  AND3_X1   g0286(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n482), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT81), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n482), .A2(new_n487), .A3(KEYINPUT81), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n490), .A2(new_n292), .A3(new_n491), .ZN(new_n492));
  AND2_X1   g0292(.A1(KEYINPUT5), .A2(G41), .ZN(new_n493));
  NOR2_X1   g0293(.A1(KEYINPUT5), .A2(G41), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n219), .B(G45), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  OR2_X1    g0295(.A1(new_n495), .A2(new_n281), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n299), .A2(G257), .A3(new_n495), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n492), .A2(G190), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n258), .A2(new_n290), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT6), .ZN(new_n501));
  INV_X1    g0301(.A(G107), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n215), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(G97), .A2(G107), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n501), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n502), .A2(KEYINPUT6), .A3(G97), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OR2_X1    g0307(.A1(new_n507), .A2(new_n220), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n500), .B(new_n508), .C1(new_n420), .C2(new_n502), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n509), .A2(new_n266), .B1(new_n215), .B2(new_n269), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n219), .A2(G33), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n270), .A2(new_n273), .A3(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G97), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n498), .A2(new_n510), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n492), .A2(new_n496), .A3(new_n497), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT82), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT82), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n492), .A2(new_n518), .A3(new_n496), .A4(new_n497), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(G200), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n510), .A2(new_n514), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n492), .A2(new_n342), .A3(new_n496), .A4(new_n497), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n516), .A2(new_n324), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n515), .A2(new_n520), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n299), .A2(new_n495), .A3(G270), .ZN(new_n526));
  XNOR2_X1  g0326(.A(new_n526), .B(KEYINPUT84), .ZN(new_n527));
  INV_X1    g0327(.A(new_n292), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n230), .A2(G1698), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n216), .A2(new_n287), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n404), .A2(new_n405), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n312), .A2(G303), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n528), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n496), .ZN(new_n534));
  NOR3_X1   g0334(.A1(new_n527), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n270), .A2(G116), .A3(new_n273), .A4(new_n511), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n228), .A2(G1), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n537), .A2(G20), .A3(new_n210), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n265), .A2(new_n225), .B1(G20), .B2(new_n210), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n486), .B(new_n220), .C1(G33), .C2(new_n215), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n539), .A2(KEYINPUT20), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT20), .B1(new_n539), .B2(new_n540), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n536), .B(new_n538), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G169), .ZN(new_n544));
  OAI21_X1  g0344(.A(KEYINPUT21), .B1(new_n535), .B2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT84), .ZN(new_n546));
  XNOR2_X1  g0346(.A(new_n526), .B(new_n546), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n531), .A2(new_n532), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n547), .B(new_n496), .C1(new_n528), .C2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT21), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n549), .A2(new_n550), .A3(G169), .A4(new_n543), .ZN(new_n551));
  INV_X1    g0351(.A(new_n543), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n552), .A2(new_n342), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n545), .A2(new_n551), .B1(new_n535), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n549), .A2(G200), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n555), .B(new_n552), .C1(new_n346), .C2(new_n549), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n404), .A2(new_n220), .A3(G68), .A4(new_n405), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT19), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n558), .A2(new_n220), .A3(G33), .A4(G97), .ZN(new_n559));
  INV_X1    g0359(.A(G87), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n504), .A2(new_n560), .B1(new_n359), .B2(new_n220), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n559), .B1(new_n561), .B2(new_n558), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n273), .B1(new_n557), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n326), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n270), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n512), .A2(new_n326), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(KEYINPUT83), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT83), .ZN(new_n570));
  NOR4_X1   g0370(.A1(new_n563), .A2(new_n570), .A3(new_n567), .A4(new_n565), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n219), .A2(G45), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n299), .A2(G250), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n214), .A2(new_n287), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n481), .A2(G1698), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n404), .A2(new_n405), .A3(new_n575), .A4(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n416), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G116), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n574), .B1(new_n580), .B2(new_n292), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n573), .A2(new_n281), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n581), .A2(G179), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n528), .B1(new_n577), .B2(new_n579), .ZN(new_n585));
  NOR3_X1   g0385(.A1(new_n585), .A2(new_n582), .A3(new_n574), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n584), .B1(new_n586), .B2(new_n324), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n572), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(G200), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n589), .B1(new_n581), .B2(new_n583), .ZN(new_n590));
  NOR4_X1   g0390(.A1(new_n585), .A2(new_n346), .A3(new_n582), .A4(new_n574), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n566), .B1(new_n560), .B2(new_n512), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n554), .A2(new_n556), .A3(new_n588), .A4(new_n595), .ZN(new_n596));
  OR3_X1    g0396(.A1(new_n560), .A2(KEYINPUT22), .A3(G20), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n597), .A2(new_n312), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n404), .A2(new_n220), .A3(G87), .A4(new_n405), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT22), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT85), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT85), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n599), .A2(new_n602), .A3(KEYINPUT22), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n598), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n578), .A2(new_n220), .A3(G116), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n220), .A2(G107), .ZN(new_n606));
  XNOR2_X1  g0406(.A(new_n606), .B(KEYINPUT23), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(KEYINPUT24), .B1(new_n604), .B2(new_n608), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n599), .A2(new_n602), .A3(KEYINPUT22), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n602), .B1(new_n599), .B2(KEYINPUT22), .ZN(new_n611));
  OAI22_X1  g0411(.A1(new_n610), .A2(new_n611), .B1(new_n312), .B2(new_n597), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT24), .ZN(new_n613));
  INV_X1    g0413(.A(new_n608), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n273), .B1(new_n609), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n537), .A2(new_n606), .ZN(new_n617));
  NAND2_X1  g0417(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n620));
  XNOR2_X1  g0420(.A(new_n619), .B(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n621), .B1(G107), .B2(new_n513), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n216), .A2(G1698), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n227), .A2(new_n287), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n404), .A2(new_n405), .A3(new_n624), .A4(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n578), .A2(G294), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n528), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n299), .A2(G264), .A3(new_n495), .ZN(new_n629));
  NOR4_X1   g0429(.A1(new_n628), .A2(G190), .A3(new_n534), .A4(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n496), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n630), .B1(new_n632), .B2(new_n589), .ZN(new_n633));
  NOR3_X1   g0433(.A1(new_n616), .A2(new_n623), .A3(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n596), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n632), .A2(new_n324), .ZN(new_n636));
  INV_X1    g0436(.A(new_n632), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n342), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n636), .B(new_n638), .C1(new_n616), .C2(new_n623), .ZN(new_n639));
  AND4_X1   g0439(.A1(new_n479), .A2(new_n525), .A3(new_n635), .A4(new_n639), .ZN(G372));
  AOI22_X1  g0440(.A1(new_n572), .A2(new_n587), .B1(new_n592), .B2(new_n594), .ZN(new_n641));
  XOR2_X1   g0441(.A(KEYINPUT88), .B(KEYINPUT26), .Z(new_n642));
  NAND4_X1  g0442(.A1(new_n523), .A2(new_n641), .A3(new_n524), .A4(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n524), .A2(new_n521), .A3(new_n522), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n593), .A2(KEYINPUT87), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT87), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n566), .B(new_n646), .C1(new_n560), .C2(new_n512), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n592), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n566), .A2(new_n568), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n587), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n644), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n643), .B1(new_n652), .B2(KEYINPUT26), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n639), .A2(new_n554), .ZN(new_n654));
  INV_X1    g0454(.A(new_n651), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n520), .A2(new_n515), .ZN(new_n657));
  INV_X1    g0457(.A(new_n616), .ZN(new_n658));
  INV_X1    g0458(.A(new_n633), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(new_n659), .A3(new_n622), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n657), .A2(new_n644), .A3(new_n660), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n653), .B(new_n650), .C1(new_n656), .C2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n479), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n459), .A2(new_n465), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n382), .A2(new_n340), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(new_n385), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n472), .A2(new_n473), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n353), .B1(new_n668), .B2(new_n311), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n663), .A2(new_n669), .ZN(G369));
  NAND2_X1  g0470(.A1(new_n537), .A2(new_n220), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(KEYINPUT89), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n672), .A2(KEYINPUT89), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n673), .A2(G213), .A3(new_n674), .A4(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n639), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n678), .B1(new_n616), .B2(new_n623), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n660), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n680), .B1(new_n639), .B2(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n554), .A2(new_n678), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(new_n680), .ZN(new_n686));
  INV_X1    g0486(.A(new_n554), .ZN(new_n687));
  INV_X1    g0487(.A(new_n678), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(new_n552), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n554), .A2(new_n556), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n690), .B1(new_n691), .B2(new_n689), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G330), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n683), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n686), .A2(new_n695), .ZN(G399));
  NOR2_X1   g0496(.A1(new_n229), .A2(G41), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR4_X1   g0498(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(G1), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n224), .B2(new_n698), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n701), .B(KEYINPUT28), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT29), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n662), .A2(new_n703), .A3(new_n688), .ZN(new_n704));
  INV_X1    g0504(.A(new_n650), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n657), .A2(new_n644), .A3(new_n660), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n651), .B1(new_n639), .B2(new_n554), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n642), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n588), .A2(new_n595), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n709), .B1(new_n644), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT91), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n652), .A2(KEYINPUT26), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT91), .ZN(new_n714));
  OAI211_X1 g0514(.A(new_n714), .B(new_n709), .C1(new_n644), .C2(new_n710), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n712), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n678), .B1(new_n708), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n704), .B1(new_n717), .B2(new_n703), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n635), .A2(new_n525), .A3(new_n639), .A4(new_n688), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n535), .A2(G179), .A3(new_n586), .A4(new_n631), .ZN(new_n720));
  OAI21_X1  g0520(.A(KEYINPUT90), .B1(new_n516), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(KEYINPUT30), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n637), .A2(G179), .A3(new_n586), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n723), .A2(new_n516), .A3(new_n549), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT30), .ZN(new_n725));
  OAI211_X1 g0525(.A(KEYINPUT90), .B(new_n725), .C1(new_n516), .C2(new_n720), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n722), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n678), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n719), .A2(KEYINPUT31), .A3(new_n728), .ZN(new_n729));
  OR2_X1    g0529(.A1(new_n728), .A2(KEYINPUT31), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n729), .A2(G330), .A3(new_n730), .ZN(new_n731));
  OR2_X1    g0531(.A1(new_n718), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n702), .B1(new_n733), .B2(G1), .ZN(new_n734));
  XOR2_X1   g0534(.A(new_n734), .B(KEYINPUT92), .Z(G364));
  NOR2_X1   g0535(.A1(new_n228), .A2(G20), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n219), .B1(new_n736), .B2(G45), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n697), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n225), .B1(G20), .B2(new_n324), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n220), .A2(new_n342), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n742), .A2(new_n346), .A3(G200), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT33), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n744), .B1(new_n745), .B2(G317), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n746), .B1(new_n745), .B2(G317), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G179), .A2(G200), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n220), .B1(new_n748), .B2(G190), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI211_X1 g0550(.A(new_n289), .B(new_n747), .C1(G294), .C2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n220), .A2(new_n346), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n752), .A2(G179), .A3(new_n589), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G322), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n742), .A2(G190), .A3(G200), .ZN(new_n756));
  XNOR2_X1  g0556(.A(new_n756), .B(KEYINPUT96), .ZN(new_n757));
  XNOR2_X1  g0557(.A(KEYINPUT97), .B(G326), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n220), .A2(G190), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n589), .A2(G179), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G283), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n760), .A2(G179), .A3(new_n589), .ZN(new_n765));
  INV_X1    g0565(.A(G311), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n752), .A2(new_n761), .ZN(new_n767));
  INV_X1    g0567(.A(G303), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n765), .A2(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n760), .A2(new_n748), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n764), .B(new_n769), .C1(G329), .C2(new_n771), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n751), .A2(new_n755), .A3(new_n759), .A4(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n289), .B1(new_n762), .B2(new_n502), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n770), .A2(new_n396), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT32), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n775), .A2(new_n776), .B1(new_n202), .B2(new_n743), .ZN(new_n777));
  INV_X1    g0577(.A(new_n767), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n774), .B(new_n777), .C1(G87), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n754), .A2(G58), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n775), .A2(new_n776), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(new_n215), .B2(new_n749), .ZN(new_n782));
  INV_X1    g0582(.A(new_n756), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n782), .B1(G50), .B2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n765), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n785), .A2(KEYINPUT95), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(KEYINPUT95), .ZN(new_n787));
  AND2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G77), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n779), .A2(new_n780), .A3(new_n784), .A4(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n741), .B1(new_n773), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G13), .A2(G33), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT93), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(new_n220), .ZN(new_n794));
  XOR2_X1   g0594(.A(new_n794), .B(KEYINPUT94), .Z(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n740), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n445), .A2(new_n229), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n799), .B1(new_n244), .B2(G45), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(G45), .B2(new_n224), .ZN(new_n801));
  INV_X1    g0601(.A(new_n229), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n802), .A2(G355), .A3(new_n289), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n801), .B(new_n803), .C1(G116), .C2(new_n802), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n791), .B1(new_n797), .B2(new_n804), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n739), .B(new_n805), .C1(new_n692), .C2(new_n795), .ZN(new_n806));
  INV_X1    g0606(.A(new_n739), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n693), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n692), .A2(G330), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n806), .B1(new_n808), .B2(new_n809), .ZN(G396));
  NAND2_X1  g0610(.A1(new_n662), .A2(new_n688), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n334), .A2(new_n678), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n352), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n340), .B2(new_n812), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n811), .B(new_n814), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(new_n731), .Z(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n807), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n788), .A2(G116), .B1(G303), .B2(new_n783), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n763), .B2(new_n743), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT98), .ZN(new_n820));
  INV_X1    g0620(.A(G294), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n753), .A2(new_n821), .B1(new_n749), .B2(new_n215), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT99), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n822), .A2(new_n823), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n312), .B1(new_n770), .B2(new_n766), .C1(new_n502), .C2(new_n767), .ZN(new_n826));
  NOR3_X1   g0626(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n820), .B(new_n827), .C1(new_n560), .C2(new_n762), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n788), .A2(G159), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n754), .A2(G143), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n744), .A2(G150), .B1(new_n783), .B2(G137), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT34), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n771), .A2(G132), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n832), .A2(new_n833), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n767), .A2(new_n205), .B1(new_n762), .B2(new_n202), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT100), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n427), .B(new_n838), .C1(G58), .C2(new_n750), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n834), .A2(new_n835), .A3(new_n836), .A4(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n741), .B1(new_n828), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n740), .A2(new_n792), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n841), .B1(new_n290), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n793), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n843), .B(new_n739), .C1(new_n844), .C2(new_n814), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n817), .A2(new_n845), .ZN(G384));
  NOR2_X1   g0646(.A1(new_n382), .A2(new_n678), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  AND3_X1   g0648(.A1(new_n460), .A2(new_n461), .A3(new_n464), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n461), .B1(new_n460), .B2(new_n464), .ZN(new_n850));
  AND3_X1   g0650(.A1(new_n468), .A2(new_n469), .A3(KEYINPUT18), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT18), .B1(new_n468), .B2(new_n469), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n849), .A2(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n676), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n469), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n469), .B1(new_n468), .B2(new_n854), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT37), .ZN(new_n859));
  AND3_X1   g0659(.A1(new_n858), .A2(new_n859), .A3(new_n458), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n859), .B1(new_n858), .B2(new_n458), .ZN(new_n861));
  OAI21_X1  g0661(.A(KEYINPUT102), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n458), .A2(new_n470), .A3(new_n855), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(KEYINPUT37), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT102), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n858), .A2(new_n859), .A3(new_n458), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n857), .A2(new_n862), .A3(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT38), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT39), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n412), .A2(new_n266), .A3(new_n432), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT16), .B1(new_n431), .B2(new_n399), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n439), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n853), .A2(new_n854), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n854), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n874), .A2(new_n468), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n876), .A2(new_n877), .A3(new_n458), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT37), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n866), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n875), .A2(KEYINPUT38), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n870), .A2(new_n871), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n860), .B1(KEYINPUT37), .B2(new_n878), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n876), .B1(new_n664), .B2(new_n667), .ZN(new_n884));
  NOR3_X1   g0684(.A1(new_n883), .A2(new_n884), .A3(new_n869), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT38), .B1(new_n875), .B2(new_n880), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT39), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n848), .B1(new_n882), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n381), .A2(new_n678), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n386), .B(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n662), .A2(new_n688), .A3(new_n814), .ZN(new_n891));
  OR2_X1    g0691(.A1(new_n340), .A2(new_n678), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n892), .B(KEYINPUT101), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n890), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n869), .B1(new_n883), .B2(new_n884), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n881), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n667), .A2(new_n854), .ZN(new_n898));
  NOR3_X1   g0698(.A1(new_n888), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n669), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n718), .B2(new_n479), .ZN(new_n901));
  XOR2_X1   g0701(.A(new_n899), .B(new_n901), .Z(new_n902));
  INV_X1    g0702(.A(new_n890), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n729), .A2(new_n903), .A3(new_n730), .A4(new_n814), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n881), .B2(new_n870), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT40), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n896), .A2(new_n906), .ZN(new_n907));
  OAI22_X1  g0707(.A1(new_n905), .A2(new_n906), .B1(new_n907), .B2(new_n904), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n729), .A2(new_n730), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n479), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n908), .B(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(G330), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n902), .B(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n219), .B2(new_n736), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT35), .ZN(new_n915));
  AOI211_X1 g0715(.A(new_n220), .B(new_n225), .C1(new_n507), .C2(new_n915), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n916), .B(G116), .C1(new_n915), .C2(new_n507), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT36), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n391), .A2(G77), .ZN(new_n919));
  OAI22_X1  g0719(.A1(new_n224), .A2(new_n919), .B1(G50), .B2(new_n202), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n920), .A2(G1), .A3(new_n228), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n914), .A2(new_n918), .A3(new_n921), .ZN(G367));
  NAND2_X1  g0722(.A1(new_n521), .A2(new_n678), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n525), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n644), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n678), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n685), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT42), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n639), .B1(new_n515), .B2(new_n520), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n688), .B1(new_n931), .B2(new_n925), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n928), .A2(new_n929), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n930), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n645), .A2(new_n647), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n678), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n655), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n650), .B2(new_n936), .ZN(new_n938));
  OR3_X1    g0738(.A1(new_n934), .A2(KEYINPUT43), .A3(new_n938), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n938), .B(KEYINPUT43), .Z(new_n940));
  NAND2_X1  g0740(.A1(new_n934), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(KEYINPUT103), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT103), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n934), .A2(new_n943), .A3(new_n940), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n939), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n927), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n945), .B1(new_n695), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n695), .A2(new_n946), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n939), .A2(new_n942), .A3(new_n948), .A4(new_n944), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n697), .B(KEYINPUT41), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n686), .A2(new_n927), .ZN(new_n952));
  XOR2_X1   g0752(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n953));
  XNOR2_X1  g0753(.A(new_n952), .B(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n946), .B1(new_n685), .B2(new_n680), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT44), .Z(new_n956));
  OAI211_X1 g0756(.A(new_n954), .B(new_n956), .C1(KEYINPUT105), .C2(new_n695), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n695), .A2(KEYINPUT105), .ZN(new_n958));
  INV_X1    g0758(.A(new_n953), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n952), .B(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n955), .B(KEYINPUT44), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n683), .B(new_n684), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(new_n694), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n957), .A2(new_n962), .A3(new_n733), .A4(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n951), .B1(new_n965), .B2(new_n733), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n947), .B(new_n949), .C1(new_n966), .C2(new_n738), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n445), .B1(new_n788), .B2(G283), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n771), .A2(G317), .ZN(new_n969));
  AOI21_X1  g0769(.A(KEYINPUT106), .B1(new_n778), .B2(G116), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT46), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n743), .A2(new_n821), .B1(new_n749), .B2(new_n502), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n753), .A2(new_n768), .B1(new_n762), .B2(new_n215), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n972), .B(new_n973), .C1(new_n757), .C2(G311), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n968), .A2(new_n969), .A3(new_n971), .A4(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(G137), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n767), .A2(new_n201), .B1(new_n770), .B2(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT107), .Z(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(G143), .B2(new_n757), .ZN(new_n979));
  INV_X1    g0779(.A(new_n762), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(G77), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n749), .A2(new_n202), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(G159), .B2(new_n744), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n259), .B2(new_n753), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(G50), .B2(new_n788), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n979), .A2(new_n981), .A3(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n975), .B1(new_n986), .B2(new_n312), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT47), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n807), .B1(new_n988), .B2(new_n740), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n797), .B1(new_n802), .B2(new_n326), .C1(new_n240), .C2(new_n799), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n989), .B(new_n990), .C1(new_n795), .C2(new_n938), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n967), .A2(new_n991), .ZN(G387));
  NOR2_X1   g0792(.A1(new_n683), .A2(new_n795), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n778), .A2(G294), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n788), .A2(G303), .B1(G317), .B2(new_n754), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n757), .A2(G322), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n995), .B(new_n996), .C1(new_n766), .C2(new_n743), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT48), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n994), .B1(new_n763), .B2(new_n749), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT109), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n997), .A2(new_n998), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT110), .Z(new_n1003));
  OR2_X1    g0803(.A1(new_n1003), .A2(KEYINPUT49), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(KEYINPUT49), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n980), .A2(G116), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n445), .B1(new_n771), .B2(new_n758), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n767), .A2(new_n290), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(G50), .A2(new_n754), .B1(new_n785), .B2(G68), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n259), .B2(new_n770), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n1009), .B(new_n1011), .C1(G97), .C2(new_n980), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n783), .A2(G159), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT108), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n750), .A2(new_n564), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n427), .B1(new_n436), .B2(new_n744), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1012), .A2(new_n1014), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n741), .B1(new_n1008), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n799), .B1(new_n237), .B2(G45), .ZN(new_n1019));
  NOR3_X1   g0819(.A1(new_n229), .A2(new_n699), .A3(new_n312), .ZN(new_n1020));
  INV_X1    g0820(.A(G45), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n330), .A2(G50), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1021), .B1(new_n1023), .B2(KEYINPUT50), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT50), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n699), .B1(new_n202), .B2(new_n290), .C1(new_n1022), .C2(new_n1025), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n1019), .A2(new_n1020), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n229), .A2(new_n502), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n993), .B(new_n1018), .C1(new_n797), .C2(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n1030), .A2(new_n739), .B1(new_n738), .B2(new_n964), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n964), .A2(new_n733), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n964), .A2(new_n733), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1032), .A2(new_n697), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1031), .A2(new_n1034), .ZN(G393));
  AND3_X1   g0835(.A1(new_n954), .A2(new_n956), .A3(new_n695), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n695), .B1(new_n954), .B2(new_n956), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1033), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1038), .A2(new_n965), .A3(new_n697), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n330), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n788), .A2(new_n1040), .B1(G50), .B2(new_n744), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT113), .Z(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n290), .B2(new_n749), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT114), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n753), .A2(new_n396), .B1(new_n756), .B2(new_n259), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT51), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n427), .B(new_n1048), .C1(G143), .C2(new_n771), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n767), .A2(new_n202), .B1(new_n762), .B2(new_n560), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1045), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n754), .A2(G311), .B1(new_n783), .B2(G317), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT52), .Z(new_n1054));
  NAND2_X1  g0854(.A1(new_n785), .A2(G294), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(G283), .A2(new_n778), .B1(new_n771), .B2(G322), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n743), .A2(new_n768), .B1(new_n762), .B2(new_n502), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n289), .B(new_n1057), .C1(G116), .C2(new_n750), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .A4(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n741), .B1(new_n1052), .B2(new_n1059), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n797), .B1(new_n215), .B2(new_n802), .C1(new_n247), .C2(new_n799), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n739), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT112), .Z(new_n1063));
  OR2_X1    g0863(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT115), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n927), .A2(new_n795), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1069), .A2(KEYINPUT111), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n1069), .A2(KEYINPUT111), .ZN(new_n1071));
  NOR4_X1   g0871(.A1(new_n1066), .A2(new_n1067), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1072), .B1(new_n1073), .B2(new_n738), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1039), .A2(new_n1074), .ZN(G390));
  INV_X1    g0875(.A(KEYINPUT119), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n729), .A2(new_n730), .A3(G330), .A4(new_n814), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1077), .A2(new_n890), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n882), .B(new_n887), .C1(new_n847), .C2(new_n894), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n870), .A2(new_n881), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n892), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n717), .B2(new_n814), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n848), .B(new_n1080), .C1(new_n1082), .C2(new_n890), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1078), .B1(new_n1079), .B2(new_n1083), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1079), .A2(new_n1083), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n731), .A2(KEYINPUT116), .A3(new_n814), .A4(new_n903), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT116), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n1077), .B2(new_n890), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1084), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n718), .A2(new_n479), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n479), .A2(G330), .A3(new_n909), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1091), .A2(new_n669), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(KEYINPUT117), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT117), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n901), .A2(new_n1095), .A3(new_n1092), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT118), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1077), .A2(new_n1097), .A3(new_n890), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n891), .A2(new_n893), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1078), .A2(new_n1097), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1077), .A2(new_n890), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1100), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1082), .A2(new_n1102), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n1088), .B2(new_n1086), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1094), .B(new_n1096), .C1(new_n1103), .C2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1076), .B1(new_n1090), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1089), .A2(new_n1079), .A3(new_n1083), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n1085), .B2(new_n1078), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1096), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1095), .B1(new_n901), .B2(new_n1092), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AND2_X1   g0912(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n1113), .A2(new_n1100), .B1(new_n1089), .B2(new_n1104), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1109), .A2(new_n1112), .A3(KEYINPUT119), .A4(new_n1114), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1107), .A2(new_n1115), .B1(new_n1090), .B2(new_n1106), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n697), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n882), .A2(new_n887), .A3(new_n793), .ZN(new_n1118));
  XOR2_X1   g0918(.A(KEYINPUT54), .B(G143), .Z(new_n1119));
  AOI22_X1  g0919(.A1(new_n788), .A2(new_n1119), .B1(G137), .B2(new_n744), .ZN(new_n1120));
  OR2_X1    g0920(.A1(new_n1120), .A2(KEYINPUT120), .ZN(new_n1121));
  INV_X1    g0921(.A(G125), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n289), .B1(new_n770), .B2(new_n1122), .C1(new_n205), .C2(new_n762), .ZN(new_n1123));
  OR3_X1    g0923(.A1(new_n767), .A2(KEYINPUT53), .A3(new_n259), .ZN(new_n1124));
  INV_X1    g0924(.A(G128), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n1124), .B1(new_n1125), .B2(new_n756), .C1(new_n396), .C2(new_n749), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n1123), .B(new_n1126), .C1(G132), .C2(new_n754), .ZN(new_n1127));
  OAI21_X1  g0927(.A(KEYINPUT53), .B1(new_n767), .B2(new_n259), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1120), .A2(KEYINPUT120), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1121), .A2(new_n1127), .A3(new_n1128), .A4(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n770), .A2(new_n821), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n289), .B1(new_n778), .B2(G87), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n788), .A2(G97), .B1(new_n1133), .B2(KEYINPUT121), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n743), .A2(new_n502), .B1(new_n749), .B2(new_n290), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(G283), .B2(new_n783), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n753), .A2(new_n210), .B1(new_n762), .B2(new_n202), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT121), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1137), .B1(new_n1132), .B2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1134), .A2(new_n1136), .A3(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1130), .B1(new_n1131), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n436), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n1141), .A2(new_n740), .B1(new_n1142), .B2(new_n842), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n1118), .A2(new_n1143), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1109), .A2(new_n738), .B1(new_n739), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1117), .A2(new_n1145), .ZN(G378));
  NAND2_X1  g0946(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(new_n1107), .B2(new_n1115), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n277), .A2(new_n854), .ZN(new_n1149));
  XOR2_X1   g0949(.A(new_n354), .B(new_n1149), .Z(new_n1150));
  XNOR2_X1  g0950(.A(new_n1150), .B(KEYINPUT55), .ZN(new_n1151));
  XOR2_X1   g0951(.A(new_n1151), .B(KEYINPUT56), .Z(new_n1152));
  NAND3_X1  g0952(.A1(new_n908), .A2(G330), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1152), .B1(new_n908), .B2(G330), .ZN(new_n1155));
  NOR3_X1   g0955(.A1(new_n1154), .A2(new_n899), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n899), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n908), .A2(G330), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1152), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1157), .B1(new_n1160), .B2(new_n1153), .ZN(new_n1161));
  OAI21_X1  g0961(.A(KEYINPUT57), .B1(new_n1156), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n697), .B1(new_n1148), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT124), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT57), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n899), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT123), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1160), .A2(new_n1157), .A3(new_n1153), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1156), .A2(KEYINPUT123), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1166), .B1(new_n1172), .B2(new_n1148), .ZN(new_n1173));
  OAI211_X1 g0973(.A(KEYINPUT124), .B(new_n697), .C1(new_n1148), .C2(new_n1162), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1165), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1170), .A2(new_n1171), .A3(new_n738), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n807), .B1(new_n205), .B2(new_n842), .ZN(new_n1177));
  XOR2_X1   g0977(.A(new_n1177), .B(KEYINPUT122), .Z(new_n1178));
  OAI22_X1  g0978(.A1(new_n756), .A2(new_n1122), .B1(new_n749), .B2(new_n259), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n754), .A2(G128), .B1(new_n778), .B2(new_n1119), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n976), .B2(new_n765), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1179), .B(new_n1181), .C1(G132), .C2(new_n744), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT59), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n257), .B1(new_n396), .B2(new_n762), .C1(new_n1182), .C2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1185));
  AOI21_X1  g0985(.A(G41), .B1(new_n771), .B2(G124), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(G41), .B1(new_n445), .B2(G33), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n1184), .A2(new_n1187), .B1(G50), .B2(new_n1188), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n762), .A2(new_n201), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n564), .B2(new_n785), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n754), .A2(G107), .B1(new_n771), .B2(G283), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1191), .A2(new_n1192), .A3(new_n295), .A4(new_n427), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n743), .A2(new_n215), .B1(new_n756), .B2(new_n210), .ZN(new_n1194));
  NOR4_X1   g0994(.A1(new_n1193), .A2(new_n982), .A3(new_n1009), .A4(new_n1194), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT58), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n740), .B1(new_n1189), .B2(new_n1196), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1178), .B(new_n1197), .C1(new_n1159), .C2(new_n844), .ZN(new_n1198));
  AND2_X1   g0998(.A1(new_n1176), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1175), .A2(new_n1199), .ZN(G375));
  NOR2_X1   g1000(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1147), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1202), .A2(new_n950), .A3(new_n1106), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n890), .A2(new_n792), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n744), .A2(G116), .B1(new_n783), .B2(G294), .ZN(new_n1205));
  AND4_X1   g1005(.A1(new_n312), .A2(new_n1205), .A3(new_n981), .A4(new_n1015), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n788), .A2(G107), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n754), .A2(G283), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(G97), .A2(new_n778), .B1(new_n771), .B2(G303), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n753), .A2(new_n976), .B1(new_n767), .B2(new_n396), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1211), .A2(new_n427), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1190), .B1(G132), .B2(new_n783), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n785), .A2(G150), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n744), .A2(new_n1119), .B1(new_n750), .B2(G50), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n770), .A2(new_n1125), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1210), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1218), .A2(new_n740), .B1(new_n202), .B2(new_n842), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1204), .A2(new_n739), .A3(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n1114), .B2(new_n738), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1203), .A2(new_n1221), .ZN(G381));
  NOR2_X1   g1022(.A1(G375), .A2(G378), .ZN(new_n1223));
  NOR3_X1   g1023(.A1(G393), .A2(G396), .A3(G381), .ZN(new_n1224));
  NOR3_X1   g1024(.A1(G387), .A2(G384), .A3(G390), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .ZN(G407));
  NAND2_X1  g1026(.A1(new_n677), .A2(G213), .ZN(new_n1227));
  XOR2_X1   g1027(.A(new_n1227), .B(KEYINPUT125), .Z(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1223), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(G407), .A2(G213), .A3(new_n1230), .ZN(G409));
  AOI21_X1  g1031(.A(G390), .B1(new_n967), .B2(new_n991), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  XOR2_X1   g1033(.A(G393), .B(G396), .Z(new_n1234));
  NAND3_X1  g1034(.A1(new_n967), .A2(new_n991), .A3(G390), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(G393), .B(G396), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1235), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1237), .B1(new_n1238), .B2(new_n1232), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1236), .A2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1175), .A2(G378), .A3(new_n1199), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n738), .B1(new_n1156), .B2(new_n1161), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n1172), .A2(new_n1148), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1198), .B(new_n1242), .C1(new_n1243), .C2(new_n951), .ZN(new_n1244));
  INV_X1    g1044(.A(G378), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1241), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1227), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT60), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n698), .B1(new_n1202), .B2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1147), .A2(new_n1201), .A3(KEYINPUT60), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1250), .A2(new_n1106), .A3(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1252), .A2(G384), .A3(new_n1221), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(G384), .B1(new_n1252), .B2(new_n1221), .ZN(new_n1255));
  OAI211_X1 g1055(.A(G2897), .B(new_n1229), .C1(new_n1254), .C2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1255), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n677), .A2(G213), .A3(G2897), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1257), .A2(new_n1253), .A3(new_n1258), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1256), .A2(new_n1259), .A3(KEYINPUT127), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT127), .B1(new_n1256), .B2(new_n1259), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1240), .B1(new_n1248), .B2(new_n1262), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1247), .A2(new_n1227), .A3(new_n1264), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT61), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1229), .B1(new_n1241), .B2(new_n1246), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1269), .A2(KEYINPUT63), .A3(new_n1264), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1263), .A2(new_n1267), .A3(new_n1268), .A4(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1256), .A2(new_n1259), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1268), .B1(new_n1269), .B2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT62), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1265), .A2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1269), .A2(KEYINPUT62), .A3(new_n1264), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1273), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1240), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1271), .B1(new_n1277), .B2(new_n1278), .ZN(G405));
  NAND2_X1  g1079(.A1(G375), .A2(new_n1245), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n1241), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1264), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1281), .A2(new_n1264), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1240), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1284), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1286), .A2(new_n1278), .A3(new_n1282), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1285), .A2(new_n1287), .ZN(G402));
endmodule


