

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U320 ( .A(n291), .B(n290), .ZN(n350) );
  INV_X1 U321 ( .A(KEYINPUT108), .ZN(n455) );
  XOR2_X1 U322 ( .A(KEYINPUT89), .B(n350), .Z(n352) );
  AND2_X1 U323 ( .A1(n464), .A2(n463), .ZN(n465) );
  XNOR2_X1 U324 ( .A(n359), .B(n289), .ZN(n360) );
  XNOR2_X1 U325 ( .A(n446), .B(KEYINPUT104), .ZN(n527) );
  XOR2_X1 U326 ( .A(n439), .B(n438), .Z(n288) );
  XOR2_X1 U327 ( .A(n358), .B(n357), .Z(n289) );
  INV_X1 U328 ( .A(KEYINPUT64), .ZN(n450) );
  XNOR2_X1 U329 ( .A(n450), .B(KEYINPUT45), .ZN(n451) );
  XNOR2_X1 U330 ( .A(n293), .B(n292), .ZN(n294) );
  XNOR2_X1 U331 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U332 ( .A(n350), .B(n294), .ZN(n297) );
  NOR2_X1 U333 ( .A1(n461), .A2(n541), .ZN(n462) );
  XNOR2_X1 U334 ( .A(n303), .B(n302), .ZN(n304) );
  NOR2_X1 U335 ( .A1(n577), .A2(n444), .ZN(n445) );
  XNOR2_X1 U336 ( .A(n440), .B(n288), .ZN(n441) );
  XNOR2_X1 U337 ( .A(n305), .B(n304), .ZN(n310) );
  XNOR2_X1 U338 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U339 ( .A(n442), .B(n441), .ZN(n460) );
  INV_X1 U340 ( .A(G106GAT), .ZN(n447) );
  XOR2_X1 U341 ( .A(KEYINPUT28), .B(n469), .Z(n520) );
  XNOR2_X1 U342 ( .A(n485), .B(KEYINPUT120), .ZN(n486) );
  XNOR2_X1 U343 ( .A(n447), .B(KEYINPUT44), .ZN(n448) );
  XNOR2_X1 U344 ( .A(n487), .B(n486), .ZN(G1351GAT) );
  XOR2_X1 U345 ( .A(G78GAT), .B(G148GAT), .Z(n291) );
  XNOR2_X1 U346 ( .A(G106GAT), .B(G204GAT), .ZN(n290) );
  NAND2_X1 U347 ( .A1(G230GAT), .A2(G233GAT), .ZN(n293) );
  INV_X1 U348 ( .A(KEYINPUT31), .ZN(n292) );
  INV_X1 U349 ( .A(n297), .ZN(n295) );
  NAND2_X1 U350 ( .A1(n295), .A2(KEYINPUT76), .ZN(n299) );
  INV_X1 U351 ( .A(KEYINPUT76), .ZN(n296) );
  NAND2_X1 U352 ( .A1(n297), .A2(n296), .ZN(n298) );
  NAND2_X1 U353 ( .A1(n299), .A2(n298), .ZN(n305) );
  XOR2_X1 U354 ( .A(G99GAT), .B(G85GAT), .Z(n428) );
  XNOR2_X1 U355 ( .A(G120GAT), .B(n428), .ZN(n303) );
  XOR2_X1 U356 ( .A(KEYINPUT33), .B(KEYINPUT75), .Z(n301) );
  XNOR2_X1 U357 ( .A(KEYINPUT74), .B(KEYINPUT32), .ZN(n300) );
  XNOR2_X1 U358 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U359 ( .A(G176GAT), .B(G92GAT), .ZN(n306) );
  XNOR2_X1 U360 ( .A(n306), .B(G64GAT), .ZN(n389) );
  XOR2_X1 U361 ( .A(KEYINPUT73), .B(KEYINPUT13), .Z(n308) );
  XNOR2_X1 U362 ( .A(G71GAT), .B(G57GAT), .ZN(n307) );
  XNOR2_X1 U363 ( .A(n308), .B(n307), .ZN(n330) );
  XNOR2_X1 U364 ( .A(n389), .B(n330), .ZN(n309) );
  XNOR2_X1 U365 ( .A(n310), .B(n309), .ZN(n573) );
  XOR2_X1 U366 ( .A(KEYINPUT41), .B(n573), .Z(n536) );
  INV_X1 U367 ( .A(n536), .ZN(n552) );
  XOR2_X1 U368 ( .A(KEYINPUT70), .B(KEYINPUT29), .Z(n312) );
  XNOR2_X1 U369 ( .A(KEYINPUT30), .B(KEYINPUT68), .ZN(n311) );
  XNOR2_X1 U370 ( .A(n312), .B(n311), .ZN(n329) );
  XOR2_X1 U371 ( .A(KEYINPUT66), .B(KEYINPUT67), .Z(n314) );
  XNOR2_X1 U372 ( .A(G113GAT), .B(G8GAT), .ZN(n313) );
  XNOR2_X1 U373 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U374 ( .A(n315), .B(G197GAT), .Z(n317) );
  XOR2_X1 U375 ( .A(G15GAT), .B(G1GAT), .Z(n331) );
  XNOR2_X1 U376 ( .A(G169GAT), .B(n331), .ZN(n316) );
  XNOR2_X1 U377 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U378 ( .A(KEYINPUT71), .B(KEYINPUT69), .Z(n319) );
  NAND2_X1 U379 ( .A1(G229GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U380 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U381 ( .A(n321), .B(n320), .Z(n327) );
  XNOR2_X1 U382 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n322) );
  XNOR2_X1 U383 ( .A(n322), .B(G29GAT), .ZN(n323) );
  XOR2_X1 U384 ( .A(n323), .B(KEYINPUT8), .Z(n325) );
  XNOR2_X1 U385 ( .A(G43GAT), .B(G50GAT), .ZN(n324) );
  XNOR2_X1 U386 ( .A(n325), .B(n324), .ZN(n440) );
  XOR2_X1 U387 ( .A(G141GAT), .B(G22GAT), .Z(n358) );
  XNOR2_X1 U388 ( .A(n440), .B(n358), .ZN(n326) );
  XNOR2_X1 U389 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U390 ( .A(n329), .B(n328), .Z(n550) );
  INV_X1 U391 ( .A(n550), .ZN(n568) );
  NOR2_X1 U392 ( .A1(n552), .A2(n568), .ZN(n514) );
  XOR2_X1 U393 ( .A(n330), .B(G155GAT), .Z(n333) );
  XNOR2_X1 U394 ( .A(G22GAT), .B(n331), .ZN(n332) );
  XNOR2_X1 U395 ( .A(n333), .B(n332), .ZN(n338) );
  XNOR2_X1 U396 ( .A(G8GAT), .B(G183GAT), .ZN(n334) );
  XNOR2_X1 U397 ( .A(n334), .B(G211GAT), .ZN(n387) );
  XOR2_X1 U398 ( .A(n387), .B(KEYINPUT14), .Z(n336) );
  NAND2_X1 U399 ( .A1(G231GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U400 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U401 ( .A(n338), .B(n337), .Z(n346) );
  XOR2_X1 U402 ( .A(KEYINPUT81), .B(G64GAT), .Z(n340) );
  XNOR2_X1 U403 ( .A(G127GAT), .B(G78GAT), .ZN(n339) );
  XNOR2_X1 U404 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U405 ( .A(KEYINPUT80), .B(KEYINPUT15), .Z(n342) );
  XNOR2_X1 U406 ( .A(KEYINPUT82), .B(KEYINPUT12), .ZN(n341) );
  XNOR2_X1 U407 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U408 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U409 ( .A(n346), .B(n345), .Z(n556) );
  INV_X1 U410 ( .A(n556), .ZN(n577) );
  XOR2_X1 U411 ( .A(KEYINPUT88), .B(KEYINPUT2), .Z(n348) );
  XNOR2_X1 U412 ( .A(KEYINPUT87), .B(G155GAT), .ZN(n347) );
  XNOR2_X1 U413 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U414 ( .A(KEYINPUT3), .B(n349), .Z(n411) );
  NAND2_X1 U415 ( .A1(G228GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U416 ( .A(n352), .B(n351), .ZN(n361) );
  XOR2_X1 U417 ( .A(G197GAT), .B(KEYINPUT21), .Z(n384) );
  XOR2_X1 U418 ( .A(G211GAT), .B(n384), .Z(n354) );
  XOR2_X1 U419 ( .A(G218GAT), .B(G162GAT), .Z(n429) );
  XNOR2_X1 U420 ( .A(G50GAT), .B(n429), .ZN(n353) );
  XNOR2_X1 U421 ( .A(n354), .B(n353), .ZN(n359) );
  XOR2_X1 U422 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n356) );
  XNOR2_X1 U423 ( .A(KEYINPUT90), .B(KEYINPUT24), .ZN(n355) );
  XNOR2_X1 U424 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U425 ( .A(n411), .B(n362), .ZN(n469) );
  XOR2_X1 U426 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n364) );
  XNOR2_X1 U427 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n363) );
  XNOR2_X1 U428 ( .A(n364), .B(n363), .ZN(n390) );
  XOR2_X1 U429 ( .A(G190GAT), .B(G134GAT), .Z(n439) );
  XOR2_X1 U430 ( .A(n390), .B(n439), .Z(n366) );
  NAND2_X1 U431 ( .A1(G227GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U432 ( .A(n366), .B(n365), .ZN(n370) );
  XOR2_X1 U433 ( .A(G71GAT), .B(KEYINPUT20), .Z(n368) );
  XNOR2_X1 U434 ( .A(G15GAT), .B(KEYINPUT86), .ZN(n367) );
  XNOR2_X1 U435 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U436 ( .A(n370), .B(n369), .Z(n379) );
  XNOR2_X1 U437 ( .A(G127GAT), .B(KEYINPUT85), .ZN(n371) );
  XNOR2_X1 U438 ( .A(n371), .B(KEYINPUT84), .ZN(n372) );
  XOR2_X1 U439 ( .A(n372), .B(KEYINPUT0), .Z(n374) );
  XNOR2_X1 U440 ( .A(G113GAT), .B(G120GAT), .ZN(n373) );
  XOR2_X1 U441 ( .A(n374), .B(n373), .Z(n419) );
  XOR2_X1 U442 ( .A(G183GAT), .B(G176GAT), .Z(n376) );
  XNOR2_X1 U443 ( .A(G43GAT), .B(G99GAT), .ZN(n375) );
  XNOR2_X1 U444 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U445 ( .A(n419), .B(n377), .Z(n378) );
  XOR2_X1 U446 ( .A(n379), .B(n378), .Z(n530) );
  INV_X1 U447 ( .A(n530), .ZN(n528) );
  NAND2_X1 U448 ( .A1(n469), .A2(n528), .ZN(n380) );
  XNOR2_X1 U449 ( .A(n380), .B(KEYINPUT26), .ZN(n566) );
  XOR2_X1 U450 ( .A(G218GAT), .B(G204GAT), .Z(n382) );
  XNOR2_X1 U451 ( .A(G36GAT), .B(G190GAT), .ZN(n381) );
  XNOR2_X1 U452 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U453 ( .A(n384), .B(n383), .Z(n386) );
  NAND2_X1 U454 ( .A1(G226GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U455 ( .A(n386), .B(n385), .ZN(n388) );
  XOR2_X1 U456 ( .A(n388), .B(n387), .Z(n392) );
  XNOR2_X1 U457 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U458 ( .A(n392), .B(n391), .ZN(n525) );
  XNOR2_X1 U459 ( .A(n525), .B(KEYINPUT27), .ZN(n423) );
  NOR2_X1 U460 ( .A1(n566), .A2(n423), .ZN(n549) );
  XOR2_X1 U461 ( .A(n549), .B(KEYINPUT98), .Z(n397) );
  NOR2_X1 U462 ( .A1(n528), .A2(n525), .ZN(n393) );
  XOR2_X1 U463 ( .A(KEYINPUT99), .B(n393), .Z(n394) );
  NOR2_X1 U464 ( .A1(n469), .A2(n394), .ZN(n395) );
  XNOR2_X1 U465 ( .A(KEYINPUT25), .B(n395), .ZN(n396) );
  NAND2_X1 U466 ( .A1(n397), .A2(n396), .ZN(n420) );
  XOR2_X1 U467 ( .A(G162GAT), .B(G148GAT), .Z(n399) );
  XNOR2_X1 U468 ( .A(G141GAT), .B(G134GAT), .ZN(n398) );
  XNOR2_X1 U469 ( .A(n399), .B(n398), .ZN(n401) );
  XOR2_X1 U470 ( .A(G29GAT), .B(G85GAT), .Z(n400) );
  XNOR2_X1 U471 ( .A(n401), .B(n400), .ZN(n415) );
  XOR2_X1 U472 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n403) );
  XNOR2_X1 U473 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n402) );
  XNOR2_X1 U474 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U475 ( .A(KEYINPUT96), .B(KEYINPUT5), .Z(n405) );
  XNOR2_X1 U476 ( .A(G1GAT), .B(G57GAT), .ZN(n404) );
  XNOR2_X1 U477 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U478 ( .A(n407), .B(n406), .Z(n413) );
  XOR2_X1 U479 ( .A(KEYINPUT94), .B(KEYINPUT91), .Z(n409) );
  XNOR2_X1 U480 ( .A(KEYINPUT95), .B(KEYINPUT4), .ZN(n408) );
  XNOR2_X1 U481 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U482 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U483 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U484 ( .A(n415), .B(n414), .ZN(n417) );
  NAND2_X1 U485 ( .A1(G225GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U486 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U487 ( .A(n419), .B(n418), .ZN(n547) );
  NAND2_X1 U488 ( .A1(n420), .A2(n547), .ZN(n426) );
  INV_X1 U489 ( .A(n547), .ZN(n421) );
  NAND2_X1 U490 ( .A1(n421), .A2(n520), .ZN(n422) );
  NOR2_X1 U491 ( .A1(n423), .A2(n422), .ZN(n531) );
  XOR2_X1 U492 ( .A(KEYINPUT97), .B(n531), .Z(n424) );
  NAND2_X1 U493 ( .A1(n424), .A2(n528), .ZN(n425) );
  NAND2_X1 U494 ( .A1(n426), .A2(n425), .ZN(n427) );
  XNOR2_X1 U495 ( .A(n427), .B(KEYINPUT100), .ZN(n492) );
  XNOR2_X1 U496 ( .A(KEYINPUT36), .B(KEYINPUT102), .ZN(n443) );
  XOR2_X1 U497 ( .A(n429), .B(n428), .Z(n431) );
  NAND2_X1 U498 ( .A1(G232GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U499 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U500 ( .A(KEYINPUT10), .B(KEYINPUT65), .Z(n433) );
  XNOR2_X1 U501 ( .A(G106GAT), .B(G92GAT), .ZN(n432) );
  XNOR2_X1 U502 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U503 ( .A(n435), .B(n434), .Z(n442) );
  XOR2_X1 U504 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n437) );
  XNOR2_X1 U505 ( .A(KEYINPUT9), .B(KEYINPUT11), .ZN(n436) );
  XNOR2_X1 U506 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U507 ( .A(n443), .B(n460), .Z(n579) );
  NAND2_X1 U508 ( .A1(n492), .A2(n579), .ZN(n444) );
  XOR2_X1 U509 ( .A(KEYINPUT37), .B(n445), .Z(n501) );
  NAND2_X1 U510 ( .A1(n514), .A2(n501), .ZN(n446) );
  NOR2_X1 U511 ( .A1(n527), .A2(n520), .ZN(n449) );
  XNOR2_X1 U512 ( .A(n449), .B(n448), .ZN(G1339GAT) );
  INV_X1 U513 ( .A(KEYINPUT113), .ZN(n473) );
  XOR2_X1 U514 ( .A(KEYINPUT72), .B(n550), .Z(n533) );
  NAND2_X1 U515 ( .A1(n579), .A2(n577), .ZN(n452) );
  INV_X1 U516 ( .A(n573), .ZN(n488) );
  NAND2_X1 U517 ( .A1(n453), .A2(n488), .ZN(n454) );
  NOR2_X1 U518 ( .A1(n533), .A2(n454), .ZN(n456) );
  XNOR2_X1 U519 ( .A(n456), .B(n455), .ZN(n464) );
  AND2_X1 U520 ( .A1(n536), .A2(n568), .ZN(n457) );
  XNOR2_X1 U521 ( .A(n457), .B(KEYINPUT46), .ZN(n458) );
  XOR2_X1 U522 ( .A(KEYINPUT106), .B(n556), .Z(n561) );
  NOR2_X1 U523 ( .A1(n458), .A2(n561), .ZN(n459) );
  XNOR2_X1 U524 ( .A(n459), .B(KEYINPUT107), .ZN(n461) );
  INV_X1 U525 ( .A(n460), .ZN(n541) );
  XNOR2_X1 U526 ( .A(n462), .B(KEYINPUT47), .ZN(n463) );
  XNOR2_X1 U527 ( .A(n465), .B(KEYINPUT48), .ZN(n546) );
  NOR2_X1 U528 ( .A1(n546), .A2(n525), .ZN(n467) );
  XNOR2_X1 U529 ( .A(KEYINPUT54), .B(KEYINPUT112), .ZN(n466) );
  XNOR2_X1 U530 ( .A(n467), .B(n466), .ZN(n468) );
  NAND2_X1 U531 ( .A1(n468), .A2(n547), .ZN(n565) );
  NOR2_X1 U532 ( .A1(n469), .A2(n565), .ZN(n470) );
  XNOR2_X1 U533 ( .A(n470), .B(KEYINPUT55), .ZN(n471) );
  NOR2_X1 U534 ( .A1(n528), .A2(n471), .ZN(n472) );
  XNOR2_X1 U535 ( .A(n473), .B(n472), .ZN(n562) );
  NAND2_X1 U536 ( .A1(n562), .A2(n536), .ZN(n479) );
  XOR2_X1 U537 ( .A(KEYINPUT118), .B(KEYINPUT117), .Z(n475) );
  XNOR2_X1 U538 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n474) );
  XNOR2_X1 U539 ( .A(n475), .B(n474), .ZN(n477) );
  XOR2_X1 U540 ( .A(G176GAT), .B(KEYINPUT116), .Z(n476) );
  XNOR2_X1 U541 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U542 ( .A(n479), .B(n478), .ZN(G1349GAT) );
  NAND2_X1 U543 ( .A1(n562), .A2(n533), .ZN(n482) );
  XOR2_X1 U544 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n480) );
  XNOR2_X1 U545 ( .A(n480), .B(G169GAT), .ZN(n481) );
  XNOR2_X1 U546 ( .A(n482), .B(n481), .ZN(G1348GAT) );
  NAND2_X1 U547 ( .A1(n541), .A2(n562), .ZN(n487) );
  XOR2_X1 U548 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n484) );
  XNOR2_X1 U549 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n483) );
  XNOR2_X1 U550 ( .A(n484), .B(n483), .ZN(n485) );
  NAND2_X1 U551 ( .A1(n488), .A2(n533), .ZN(n489) );
  XNOR2_X1 U552 ( .A(n489), .B(KEYINPUT77), .ZN(n502) );
  NAND2_X1 U553 ( .A1(n577), .A2(n460), .ZN(n490) );
  XNOR2_X1 U554 ( .A(n490), .B(KEYINPUT16), .ZN(n491) );
  XNOR2_X1 U555 ( .A(KEYINPUT83), .B(n491), .ZN(n493) );
  AND2_X1 U556 ( .A1(n493), .A2(n492), .ZN(n513) );
  NAND2_X1 U557 ( .A1(n502), .A2(n513), .ZN(n499) );
  NOR2_X1 U558 ( .A1(n547), .A2(n499), .ZN(n494) );
  XOR2_X1 U559 ( .A(G1GAT), .B(n494), .Z(n495) );
  XNOR2_X1 U560 ( .A(KEYINPUT34), .B(n495), .ZN(G1324GAT) );
  NOR2_X1 U561 ( .A1(n525), .A2(n499), .ZN(n496) );
  XOR2_X1 U562 ( .A(G8GAT), .B(n496), .Z(G1325GAT) );
  NOR2_X1 U563 ( .A1(n528), .A2(n499), .ZN(n498) );
  XNOR2_X1 U564 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n497) );
  XNOR2_X1 U565 ( .A(n498), .B(n497), .ZN(G1326GAT) );
  NOR2_X1 U566 ( .A1(n520), .A2(n499), .ZN(n500) );
  XOR2_X1 U567 ( .A(G22GAT), .B(n500), .Z(G1327GAT) );
  NAND2_X1 U568 ( .A1(n502), .A2(n501), .ZN(n503) );
  XNOR2_X1 U569 ( .A(n503), .B(KEYINPUT38), .ZN(n511) );
  NOR2_X1 U570 ( .A1(n547), .A2(n511), .ZN(n506) );
  XOR2_X1 U571 ( .A(G29GAT), .B(KEYINPUT101), .Z(n504) );
  XNOR2_X1 U572 ( .A(KEYINPUT39), .B(n504), .ZN(n505) );
  XNOR2_X1 U573 ( .A(n506), .B(n505), .ZN(G1328GAT) );
  NOR2_X1 U574 ( .A1(n525), .A2(n511), .ZN(n507) );
  XOR2_X1 U575 ( .A(G36GAT), .B(n507), .Z(G1329GAT) );
  XNOR2_X1 U576 ( .A(KEYINPUT40), .B(KEYINPUT103), .ZN(n509) );
  NOR2_X1 U577 ( .A1(n528), .A2(n511), .ZN(n508) );
  XNOR2_X1 U578 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U579 ( .A(G43GAT), .B(n510), .ZN(G1330GAT) );
  NOR2_X1 U580 ( .A1(n511), .A2(n520), .ZN(n512) );
  XOR2_X1 U581 ( .A(G50GAT), .B(n512), .Z(G1331GAT) );
  NAND2_X1 U582 ( .A1(n514), .A2(n513), .ZN(n519) );
  NOR2_X1 U583 ( .A1(n547), .A2(n519), .ZN(n515) );
  XOR2_X1 U584 ( .A(G57GAT), .B(n515), .Z(n516) );
  XNOR2_X1 U585 ( .A(KEYINPUT42), .B(n516), .ZN(G1332GAT) );
  NOR2_X1 U586 ( .A1(n525), .A2(n519), .ZN(n517) );
  XOR2_X1 U587 ( .A(G64GAT), .B(n517), .Z(G1333GAT) );
  NOR2_X1 U588 ( .A1(n528), .A2(n519), .ZN(n518) );
  XOR2_X1 U589 ( .A(G71GAT), .B(n518), .Z(G1334GAT) );
  NOR2_X1 U590 ( .A1(n520), .A2(n519), .ZN(n522) );
  XNOR2_X1 U591 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n521) );
  XNOR2_X1 U592 ( .A(n522), .B(n521), .ZN(G1335GAT) );
  NOR2_X1 U593 ( .A1(n547), .A2(n527), .ZN(n523) );
  XNOR2_X1 U594 ( .A(G85GAT), .B(n523), .ZN(n524) );
  XNOR2_X1 U595 ( .A(n524), .B(KEYINPUT105), .ZN(G1336GAT) );
  NOR2_X1 U596 ( .A1(n525), .A2(n527), .ZN(n526) );
  XOR2_X1 U597 ( .A(G92GAT), .B(n526), .Z(G1337GAT) );
  NOR2_X1 U598 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U599 ( .A(G99GAT), .B(n529), .Z(G1338GAT) );
  XOR2_X1 U600 ( .A(G113GAT), .B(KEYINPUT109), .Z(n535) );
  NAND2_X1 U601 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U602 ( .A1(n546), .A2(n532), .ZN(n542) );
  NAND2_X1 U603 ( .A1(n542), .A2(n533), .ZN(n534) );
  XNOR2_X1 U604 ( .A(n535), .B(n534), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .Z(n538) );
  NAND2_X1 U606 ( .A1(n542), .A2(n536), .ZN(n537) );
  XNOR2_X1 U607 ( .A(n538), .B(n537), .ZN(G1341GAT) );
  NAND2_X1 U608 ( .A1(n561), .A2(n542), .ZN(n539) );
  XNOR2_X1 U609 ( .A(n539), .B(KEYINPUT50), .ZN(n540) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(n540), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT110), .B(KEYINPUT51), .Z(n544) );
  NAND2_X1 U612 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U613 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U614 ( .A(G134GAT), .B(n545), .ZN(G1343GAT) );
  NOR2_X1 U615 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U616 ( .A1(n549), .A2(n548), .ZN(n559) );
  NOR2_X1 U617 ( .A1(n550), .A2(n559), .ZN(n551) );
  XOR2_X1 U618 ( .A(G141GAT), .B(n551), .Z(G1344GAT) );
  NOR2_X1 U619 ( .A1(n552), .A2(n559), .ZN(n554) );
  XNOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(n555), .ZN(G1345GAT) );
  NOR2_X1 U623 ( .A1(n556), .A2(n559), .ZN(n558) );
  XNOR2_X1 U624 ( .A(G155GAT), .B(KEYINPUT111), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(G1346GAT) );
  NOR2_X1 U626 ( .A1(n460), .A2(n559), .ZN(n560) );
  XOR2_X1 U627 ( .A(G162GAT), .B(n560), .Z(G1347GAT) );
  XOR2_X1 U628 ( .A(G183GAT), .B(KEYINPUT119), .Z(n564) );
  NAND2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1350GAT) );
  NOR2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U632 ( .A(KEYINPUT123), .B(n567), .Z(n580) );
  NAND2_X1 U633 ( .A1(n568), .A2(n580), .ZN(n572) );
  XOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n570) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1352GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n575) );
  NAND2_X1 U639 ( .A1(n580), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XOR2_X1 U641 ( .A(G204GAT), .B(n576), .Z(G1353GAT) );
  NAND2_X1 U642 ( .A1(n580), .A2(n577), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n582) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XOR2_X1 U647 ( .A(G218GAT), .B(n583), .Z(G1355GAT) );
endmodule

