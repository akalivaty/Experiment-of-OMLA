

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U552 ( .A1(n715), .A2(G2084), .ZN(n736) );
  NAND2_X1 U553 ( .A1(n769), .A2(n682), .ZN(n715) );
  INV_X1 U554 ( .A(KEYINPUT103), .ZN(n729) );
  NOR2_X2 U555 ( .A1(G2105), .A2(G2104), .ZN(n536) );
  AND2_X1 U556 ( .A1(n769), .A2(n682), .ZN(n707) );
  NOR2_X1 U557 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U558 ( .A(n730), .B(n729), .ZN(n731) );
  INV_X1 U559 ( .A(KEYINPUT101), .ZN(n740) );
  XNOR2_X1 U560 ( .A(n741), .B(n740), .ZN(n791) );
  NOR2_X1 U561 ( .A1(G651), .A2(n629), .ZN(n647) );
  AND2_X1 U562 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X1 U563 ( .A1(G651), .A2(G543), .ZN(n639) );
  NAND2_X1 U564 ( .A1(G89), .A2(n639), .ZN(n517) );
  XNOR2_X1 U565 ( .A(n517), .B(KEYINPUT4), .ZN(n518) );
  XNOR2_X1 U566 ( .A(n518), .B(KEYINPUT76), .ZN(n520) );
  XOR2_X1 U567 ( .A(KEYINPUT0), .B(G543), .Z(n629) );
  INV_X1 U568 ( .A(G651), .ZN(n522) );
  NOR2_X1 U569 ( .A1(n629), .A2(n522), .ZN(n643) );
  NAND2_X1 U570 ( .A1(G76), .A2(n643), .ZN(n519) );
  NAND2_X1 U571 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U572 ( .A(n521), .B(KEYINPUT5), .ZN(n529) );
  NOR2_X1 U573 ( .A1(G543), .A2(n522), .ZN(n523) );
  XOR2_X1 U574 ( .A(KEYINPUT1), .B(n523), .Z(n640) );
  NAND2_X1 U575 ( .A1(n640), .A2(G63), .ZN(n524) );
  XOR2_X1 U576 ( .A(KEYINPUT77), .B(n524), .Z(n526) );
  NAND2_X1 U577 ( .A1(n647), .A2(G51), .ZN(n525) );
  NAND2_X1 U578 ( .A1(n526), .A2(n525), .ZN(n527) );
  XOR2_X1 U579 ( .A(KEYINPUT6), .B(n527), .Z(n528) );
  NAND2_X1 U580 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U581 ( .A(n530), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U582 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U583 ( .A(KEYINPUT23), .B(KEYINPUT65), .Z(n532) );
  INV_X1 U584 ( .A(G2104), .ZN(n533) );
  NOR2_X2 U585 ( .A1(G2105), .A2(n533), .ZN(n880) );
  NAND2_X1 U586 ( .A1(G101), .A2(n880), .ZN(n531) );
  XNOR2_X1 U587 ( .A(n532), .B(n531), .ZN(n535) );
  AND2_X1 U588 ( .A1(n533), .A2(G2105), .ZN(n884) );
  AND2_X1 U589 ( .A1(G125), .A2(n884), .ZN(n534) );
  NOR2_X1 U590 ( .A1(n535), .A2(n534), .ZN(n542) );
  XOR2_X2 U591 ( .A(KEYINPUT17), .B(n536), .Z(n881) );
  NAND2_X1 U592 ( .A1(G137), .A2(n881), .ZN(n539) );
  NAND2_X1 U593 ( .A1(G2104), .A2(G2105), .ZN(n537) );
  XOR2_X2 U594 ( .A(KEYINPUT66), .B(n537), .Z(n885) );
  NAND2_X1 U595 ( .A1(G113), .A2(n885), .ZN(n538) );
  NAND2_X1 U596 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U597 ( .A(n540), .B(KEYINPUT67), .ZN(n541) );
  XNOR2_X1 U598 ( .A(n543), .B(KEYINPUT64), .ZN(n677) );
  BUF_X1 U599 ( .A(n677), .Z(G160) );
  AND2_X1 U600 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U601 ( .A(G108), .ZN(G238) );
  INV_X1 U602 ( .A(G132), .ZN(G219) );
  INV_X1 U603 ( .A(G82), .ZN(G220) );
  NAND2_X1 U604 ( .A1(G64), .A2(n640), .ZN(n545) );
  NAND2_X1 U605 ( .A1(G52), .A2(n647), .ZN(n544) );
  NAND2_X1 U606 ( .A1(n545), .A2(n544), .ZN(n550) );
  NAND2_X1 U607 ( .A1(G90), .A2(n639), .ZN(n547) );
  NAND2_X1 U608 ( .A1(G77), .A2(n643), .ZN(n546) );
  NAND2_X1 U609 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U610 ( .A(KEYINPUT9), .B(n548), .Z(n549) );
  NOR2_X1 U611 ( .A1(n550), .A2(n549), .ZN(G171) );
  NAND2_X1 U612 ( .A1(G62), .A2(n640), .ZN(n552) );
  NAND2_X1 U613 ( .A1(G75), .A2(n643), .ZN(n551) );
  NAND2_X1 U614 ( .A1(n552), .A2(n551), .ZN(n555) );
  NAND2_X1 U615 ( .A1(n639), .A2(G88), .ZN(n553) );
  XOR2_X1 U616 ( .A(KEYINPUT82), .B(n553), .Z(n554) );
  NOR2_X1 U617 ( .A1(n555), .A2(n554), .ZN(n557) );
  NAND2_X1 U618 ( .A1(n647), .A2(G50), .ZN(n556) );
  NAND2_X1 U619 ( .A1(n557), .A2(n556), .ZN(G303) );
  NAND2_X1 U620 ( .A1(G102), .A2(n880), .ZN(n559) );
  NAND2_X1 U621 ( .A1(G138), .A2(n881), .ZN(n558) );
  NAND2_X1 U622 ( .A1(n559), .A2(n558), .ZN(n563) );
  NAND2_X1 U623 ( .A1(n884), .A2(G126), .ZN(n561) );
  NAND2_X1 U624 ( .A1(G114), .A2(n885), .ZN(n560) );
  NAND2_X1 U625 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U626 ( .A1(n563), .A2(n562), .ZN(G164) );
  XOR2_X1 U627 ( .A(KEYINPUT71), .B(KEYINPUT10), .Z(n565) );
  NAND2_X1 U628 ( .A1(G7), .A2(G661), .ZN(n564) );
  XNOR2_X1 U629 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U630 ( .A(KEYINPUT70), .B(n566), .ZN(G223) );
  INV_X1 U631 ( .A(G223), .ZN(n827) );
  NAND2_X1 U632 ( .A1(n827), .A2(G567), .ZN(n567) );
  XOR2_X1 U633 ( .A(KEYINPUT11), .B(n567), .Z(G234) );
  NAND2_X1 U634 ( .A1(n640), .A2(G56), .ZN(n568) );
  XOR2_X1 U635 ( .A(KEYINPUT14), .B(n568), .Z(n576) );
  NAND2_X1 U636 ( .A1(n639), .A2(G81), .ZN(n569) );
  XOR2_X1 U637 ( .A(KEYINPUT12), .B(n569), .Z(n572) );
  NAND2_X1 U638 ( .A1(n643), .A2(G68), .ZN(n570) );
  XOR2_X1 U639 ( .A(n570), .B(KEYINPUT72), .Z(n571) );
  NOR2_X1 U640 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U641 ( .A(KEYINPUT13), .B(n573), .Z(n574) );
  XNOR2_X1 U642 ( .A(n574), .B(KEYINPUT73), .ZN(n575) );
  NOR2_X1 U643 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U644 ( .A1(n647), .A2(G43), .ZN(n577) );
  NAND2_X1 U645 ( .A1(n578), .A2(n577), .ZN(n970) );
  INV_X1 U646 ( .A(G860), .ZN(n616) );
  OR2_X1 U647 ( .A1(n970), .A2(n616), .ZN(G153) );
  NAND2_X1 U648 ( .A1(G868), .A2(G171), .ZN(n588) );
  NAND2_X1 U649 ( .A1(G79), .A2(n643), .ZN(n580) );
  NAND2_X1 U650 ( .A1(G54), .A2(n647), .ZN(n579) );
  NAND2_X1 U651 ( .A1(n580), .A2(n579), .ZN(n585) );
  NAND2_X1 U652 ( .A1(G92), .A2(n639), .ZN(n582) );
  NAND2_X1 U653 ( .A1(G66), .A2(n640), .ZN(n581) );
  NAND2_X1 U654 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U655 ( .A(KEYINPUT74), .B(n583), .ZN(n584) );
  NOR2_X1 U656 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U657 ( .A(n586), .B(KEYINPUT15), .ZN(n969) );
  INV_X1 U658 ( .A(n969), .ZN(n614) );
  INV_X1 U659 ( .A(G868), .ZN(n596) );
  NAND2_X1 U660 ( .A1(n614), .A2(n596), .ZN(n587) );
  NAND2_X1 U661 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U662 ( .A(n589), .B(KEYINPUT75), .ZN(G284) );
  NAND2_X1 U663 ( .A1(G65), .A2(n640), .ZN(n591) );
  NAND2_X1 U664 ( .A1(G53), .A2(n647), .ZN(n590) );
  NAND2_X1 U665 ( .A1(n591), .A2(n590), .ZN(n595) );
  NAND2_X1 U666 ( .A1(G91), .A2(n639), .ZN(n593) );
  NAND2_X1 U667 ( .A1(G78), .A2(n643), .ZN(n592) );
  NAND2_X1 U668 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U669 ( .A1(n595), .A2(n594), .ZN(n973) );
  XNOR2_X1 U670 ( .A(n973), .B(KEYINPUT69), .ZN(G299) );
  NAND2_X1 U671 ( .A1(G286), .A2(G868), .ZN(n598) );
  NAND2_X1 U672 ( .A1(G299), .A2(n596), .ZN(n597) );
  NAND2_X1 U673 ( .A1(n598), .A2(n597), .ZN(G297) );
  NAND2_X1 U674 ( .A1(n616), .A2(G559), .ZN(n599) );
  NAND2_X1 U675 ( .A1(n599), .A2(n614), .ZN(n600) );
  XNOR2_X1 U676 ( .A(n600), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U677 ( .A1(G868), .A2(n970), .ZN(n603) );
  NAND2_X1 U678 ( .A1(G868), .A2(n614), .ZN(n601) );
  NOR2_X1 U679 ( .A1(G559), .A2(n601), .ZN(n602) );
  NOR2_X1 U680 ( .A1(n603), .A2(n602), .ZN(G282) );
  NAND2_X1 U681 ( .A1(n885), .A2(G111), .ZN(n604) );
  XNOR2_X1 U682 ( .A(n604), .B(KEYINPUT78), .ZN(n611) );
  NAND2_X1 U683 ( .A1(G99), .A2(n880), .ZN(n606) );
  NAND2_X1 U684 ( .A1(G135), .A2(n881), .ZN(n605) );
  NAND2_X1 U685 ( .A1(n606), .A2(n605), .ZN(n609) );
  NAND2_X1 U686 ( .A1(n884), .A2(G123), .ZN(n607) );
  XOR2_X1 U687 ( .A(KEYINPUT18), .B(n607), .Z(n608) );
  NOR2_X1 U688 ( .A1(n609), .A2(n608), .ZN(n610) );
  NAND2_X1 U689 ( .A1(n611), .A2(n610), .ZN(n923) );
  XNOR2_X1 U690 ( .A(G2096), .B(n923), .ZN(n612) );
  NOR2_X1 U691 ( .A1(G2100), .A2(n612), .ZN(n613) );
  XNOR2_X1 U692 ( .A(KEYINPUT79), .B(n613), .ZN(G156) );
  NAND2_X1 U693 ( .A1(G559), .A2(n614), .ZN(n615) );
  XOR2_X1 U694 ( .A(n970), .B(n615), .Z(n655) );
  NAND2_X1 U695 ( .A1(n616), .A2(n655), .ZN(n624) );
  NAND2_X1 U696 ( .A1(G80), .A2(n643), .ZN(n617) );
  XNOR2_X1 U697 ( .A(n617), .B(KEYINPUT80), .ZN(n619) );
  NAND2_X1 U698 ( .A1(n640), .A2(G67), .ZN(n618) );
  NAND2_X1 U699 ( .A1(n619), .A2(n618), .ZN(n623) );
  NAND2_X1 U700 ( .A1(G93), .A2(n639), .ZN(n621) );
  NAND2_X1 U701 ( .A1(G55), .A2(n647), .ZN(n620) );
  NAND2_X1 U702 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U703 ( .A1(n623), .A2(n622), .ZN(n657) );
  XOR2_X1 U704 ( .A(n624), .B(n657), .Z(G145) );
  INV_X1 U705 ( .A(G303), .ZN(G166) );
  NAND2_X1 U706 ( .A1(G49), .A2(n647), .ZN(n626) );
  NAND2_X1 U707 ( .A1(G74), .A2(G651), .ZN(n625) );
  NAND2_X1 U708 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U709 ( .A1(n640), .A2(n627), .ZN(n628) );
  XOR2_X1 U710 ( .A(KEYINPUT81), .B(n628), .Z(n631) );
  NAND2_X1 U711 ( .A1(n629), .A2(G87), .ZN(n630) );
  NAND2_X1 U712 ( .A1(n631), .A2(n630), .ZN(G288) );
  NAND2_X1 U713 ( .A1(G60), .A2(n640), .ZN(n633) );
  NAND2_X1 U714 ( .A1(G47), .A2(n647), .ZN(n632) );
  NAND2_X1 U715 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U716 ( .A1(G85), .A2(n639), .ZN(n634) );
  XOR2_X1 U717 ( .A(KEYINPUT68), .B(n634), .Z(n635) );
  NOR2_X1 U718 ( .A1(n636), .A2(n635), .ZN(n638) );
  NAND2_X1 U719 ( .A1(n643), .A2(G72), .ZN(n637) );
  NAND2_X1 U720 ( .A1(n638), .A2(n637), .ZN(G290) );
  NAND2_X1 U721 ( .A1(G86), .A2(n639), .ZN(n642) );
  NAND2_X1 U722 ( .A1(G61), .A2(n640), .ZN(n641) );
  NAND2_X1 U723 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U724 ( .A1(n643), .A2(G73), .ZN(n644) );
  XOR2_X1 U725 ( .A(KEYINPUT2), .B(n644), .Z(n645) );
  NOR2_X1 U726 ( .A1(n646), .A2(n645), .ZN(n649) );
  NAND2_X1 U727 ( .A1(n647), .A2(G48), .ZN(n648) );
  NAND2_X1 U728 ( .A1(n649), .A2(n648), .ZN(G305) );
  XNOR2_X1 U729 ( .A(G166), .B(KEYINPUT19), .ZN(n654) );
  XNOR2_X1 U730 ( .A(n657), .B(G288), .ZN(n650) );
  XNOR2_X1 U731 ( .A(n650), .B(G299), .ZN(n651) );
  XNOR2_X1 U732 ( .A(n651), .B(G290), .ZN(n652) );
  XNOR2_X1 U733 ( .A(n652), .B(G305), .ZN(n653) );
  XNOR2_X1 U734 ( .A(n654), .B(n653), .ZN(n853) );
  XNOR2_X1 U735 ( .A(n655), .B(n853), .ZN(n656) );
  NAND2_X1 U736 ( .A1(n656), .A2(G868), .ZN(n659) );
  OR2_X1 U737 ( .A1(G868), .A2(n657), .ZN(n658) );
  NAND2_X1 U738 ( .A1(n659), .A2(n658), .ZN(G295) );
  NAND2_X1 U739 ( .A1(G2084), .A2(G2078), .ZN(n660) );
  XNOR2_X1 U740 ( .A(n660), .B(KEYINPUT20), .ZN(n661) );
  XNOR2_X1 U741 ( .A(n661), .B(KEYINPUT83), .ZN(n662) );
  NAND2_X1 U742 ( .A1(n662), .A2(G2090), .ZN(n663) );
  XNOR2_X1 U743 ( .A(KEYINPUT21), .B(n663), .ZN(n664) );
  NAND2_X1 U744 ( .A1(n664), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U745 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U746 ( .A1(G220), .A2(G219), .ZN(n665) );
  XOR2_X1 U747 ( .A(KEYINPUT22), .B(n665), .Z(n666) );
  NOR2_X1 U748 ( .A1(G218), .A2(n666), .ZN(n667) );
  NAND2_X1 U749 ( .A1(G96), .A2(n667), .ZN(n915) );
  NAND2_X1 U750 ( .A1(G2106), .A2(n915), .ZN(n673) );
  NAND2_X1 U751 ( .A1(G120), .A2(G69), .ZN(n668) );
  XOR2_X1 U752 ( .A(KEYINPUT84), .B(n668), .Z(n669) );
  NAND2_X1 U753 ( .A1(G57), .A2(n669), .ZN(n670) );
  NOR2_X1 U754 ( .A1(G238), .A2(n670), .ZN(n671) );
  XNOR2_X1 U755 ( .A(KEYINPUT85), .B(n671), .ZN(n916) );
  NAND2_X1 U756 ( .A1(G567), .A2(n916), .ZN(n672) );
  NAND2_X1 U757 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U758 ( .A(KEYINPUT86), .B(n674), .Z(G319) );
  INV_X1 U759 ( .A(G319), .ZN(n676) );
  NAND2_X1 U760 ( .A1(G661), .A2(G483), .ZN(n675) );
  NOR2_X1 U761 ( .A1(n676), .A2(n675), .ZN(n831) );
  NAND2_X1 U762 ( .A1(n831), .A2(G36), .ZN(G176) );
  INV_X1 U763 ( .A(G171), .ZN(G301) );
  NOR2_X1 U764 ( .A1(G164), .A2(G1384), .ZN(n769) );
  NAND2_X1 U765 ( .A1(n677), .A2(G40), .ZN(n768) );
  XOR2_X1 U766 ( .A(KEYINPUT94), .B(n768), .Z(n682) );
  NAND2_X1 U767 ( .A1(G8), .A2(n715), .ZN(n797) );
  NOR2_X1 U768 ( .A1(G1971), .A2(n797), .ZN(n679) );
  NOR2_X1 U769 ( .A1(G2090), .A2(n715), .ZN(n678) );
  NOR2_X1 U770 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U771 ( .A(KEYINPUT102), .B(n680), .ZN(n681) );
  NAND2_X1 U772 ( .A1(n681), .A2(G303), .ZN(n728) );
  NAND2_X1 U773 ( .A1(G2072), .A2(n707), .ZN(n684) );
  XOR2_X1 U774 ( .A(KEYINPUT98), .B(KEYINPUT27), .Z(n683) );
  XNOR2_X1 U775 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U776 ( .A(n685), .B(KEYINPUT97), .ZN(n687) );
  AND2_X1 U777 ( .A1(G1956), .A2(n715), .ZN(n686) );
  NOR2_X1 U778 ( .A1(n687), .A2(n686), .ZN(n690) );
  NOR2_X1 U779 ( .A1(n973), .A2(n690), .ZN(n689) );
  XNOR2_X1 U780 ( .A(KEYINPUT99), .B(KEYINPUT28), .ZN(n688) );
  XNOR2_X1 U781 ( .A(n689), .B(n688), .ZN(n705) );
  NAND2_X1 U782 ( .A1(n973), .A2(n690), .ZN(n703) );
  NAND2_X1 U783 ( .A1(G1348), .A2(n715), .ZN(n692) );
  NAND2_X1 U784 ( .A1(n707), .A2(G2067), .ZN(n691) );
  NAND2_X1 U785 ( .A1(n692), .A2(n691), .ZN(n697) );
  NAND2_X1 U786 ( .A1(n969), .A2(n697), .ZN(n701) );
  AND2_X1 U787 ( .A1(n707), .A2(G1996), .ZN(n693) );
  XOR2_X1 U788 ( .A(n693), .B(KEYINPUT26), .Z(n695) );
  NAND2_X1 U789 ( .A1(n715), .A2(G1341), .ZN(n694) );
  NAND2_X1 U790 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U791 ( .A1(n970), .A2(n696), .ZN(n699) );
  NOR2_X1 U792 ( .A1(n969), .A2(n697), .ZN(n698) );
  OR2_X1 U793 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U794 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U795 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U796 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U797 ( .A(n706), .B(KEYINPUT29), .ZN(n712) );
  NOR2_X1 U798 ( .A1(n707), .A2(G1961), .ZN(n708) );
  XNOR2_X1 U799 ( .A(n708), .B(KEYINPUT96), .ZN(n710) );
  XOR2_X1 U800 ( .A(G2078), .B(KEYINPUT25), .Z(n948) );
  NOR2_X1 U801 ( .A1(n715), .A2(n948), .ZN(n709) );
  NOR2_X1 U802 ( .A1(n710), .A2(n709), .ZN(n720) );
  NOR2_X1 U803 ( .A1(G301), .A2(n720), .ZN(n711) );
  NOR2_X1 U804 ( .A1(n712), .A2(n711), .ZN(n725) );
  INV_X1 U805 ( .A(G8), .ZN(n713) );
  NOR2_X1 U806 ( .A1(n713), .A2(G1966), .ZN(n714) );
  AND2_X1 U807 ( .A1(n715), .A2(n714), .ZN(n734) );
  XNOR2_X1 U808 ( .A(n736), .B(KEYINPUT95), .ZN(n716) );
  NAND2_X1 U809 ( .A1(G8), .A2(n716), .ZN(n717) );
  NOR2_X1 U810 ( .A1(n734), .A2(n717), .ZN(n718) );
  XOR2_X1 U811 ( .A(KEYINPUT30), .B(n718), .Z(n719) );
  NOR2_X1 U812 ( .A1(G168), .A2(n719), .ZN(n722) );
  AND2_X1 U813 ( .A1(G301), .A2(n720), .ZN(n721) );
  NOR2_X1 U814 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U815 ( .A(n723), .B(KEYINPUT31), .ZN(n724) );
  NOR2_X1 U816 ( .A1(n725), .A2(n724), .ZN(n733) );
  INV_X1 U817 ( .A(G286), .ZN(n726) );
  OR2_X1 U818 ( .A1(n733), .A2(n726), .ZN(n727) );
  NAND2_X1 U819 ( .A1(n728), .A2(n727), .ZN(n730) );
  NAND2_X1 U820 ( .A1(n731), .A2(G8), .ZN(n732) );
  XNOR2_X1 U821 ( .A(n732), .B(KEYINPUT32), .ZN(n792) );
  XNOR2_X1 U822 ( .A(n735), .B(KEYINPUT100), .ZN(n739) );
  XOR2_X1 U823 ( .A(KEYINPUT95), .B(n736), .Z(n737) );
  NAND2_X1 U824 ( .A1(G8), .A2(n737), .ZN(n738) );
  NAND2_X1 U825 ( .A1(n739), .A2(n738), .ZN(n741) );
  XOR2_X1 U826 ( .A(G1981), .B(G305), .Z(n987) );
  NOR2_X1 U827 ( .A1(G1976), .A2(G288), .ZN(n742) );
  XOR2_X1 U828 ( .A(KEYINPUT104), .B(n742), .Z(n984) );
  NOR2_X1 U829 ( .A1(n797), .A2(n984), .ZN(n743) );
  NAND2_X1 U830 ( .A1(KEYINPUT33), .A2(n743), .ZN(n744) );
  AND2_X1 U831 ( .A1(n987), .A2(n744), .ZN(n802) );
  NAND2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n978) );
  AND2_X1 U833 ( .A1(n802), .A2(n978), .ZN(n746) );
  AND2_X1 U834 ( .A1(n791), .A2(n746), .ZN(n745) );
  NAND2_X1 U835 ( .A1(n792), .A2(n745), .ZN(n751) );
  INV_X1 U836 ( .A(n746), .ZN(n749) );
  OR2_X1 U837 ( .A1(G1971), .A2(G303), .ZN(n747) );
  AND2_X1 U838 ( .A1(n747), .A2(n984), .ZN(n748) );
  OR2_X1 U839 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U840 ( .A1(n751), .A2(n750), .ZN(n754) );
  NOR2_X1 U841 ( .A1(G1981), .A2(G305), .ZN(n752) );
  XNOR2_X1 U842 ( .A(KEYINPUT24), .B(n752), .ZN(n753) );
  NOR2_X1 U843 ( .A1(n754), .A2(n753), .ZN(n790) );
  XOR2_X1 U844 ( .A(G2067), .B(KEYINPUT37), .Z(n755) );
  XNOR2_X1 U845 ( .A(KEYINPUT87), .B(n755), .ZN(n811) );
  NAND2_X1 U846 ( .A1(n884), .A2(G128), .ZN(n756) );
  XNOR2_X1 U847 ( .A(n756), .B(KEYINPUT90), .ZN(n758) );
  NAND2_X1 U848 ( .A1(G116), .A2(n885), .ZN(n757) );
  NAND2_X1 U849 ( .A1(n758), .A2(n757), .ZN(n759) );
  XOR2_X1 U850 ( .A(KEYINPUT35), .B(n759), .Z(n766) );
  XNOR2_X1 U851 ( .A(KEYINPUT88), .B(KEYINPUT89), .ZN(n760) );
  XNOR2_X1 U852 ( .A(n760), .B(KEYINPUT34), .ZN(n764) );
  NAND2_X1 U853 ( .A1(G104), .A2(n880), .ZN(n762) );
  NAND2_X1 U854 ( .A1(G140), .A2(n881), .ZN(n761) );
  NAND2_X1 U855 ( .A1(n762), .A2(n761), .ZN(n763) );
  XOR2_X1 U856 ( .A(n764), .B(n763), .Z(n765) );
  NOR2_X1 U857 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U858 ( .A(KEYINPUT36), .B(n767), .ZN(n896) );
  NOR2_X1 U859 ( .A1(n811), .A2(n896), .ZN(n919) );
  NOR2_X1 U860 ( .A1(n769), .A2(n768), .ZN(n821) );
  NAND2_X1 U861 ( .A1(n919), .A2(n821), .ZN(n770) );
  XOR2_X1 U862 ( .A(KEYINPUT91), .B(n770), .Z(n818) );
  NAND2_X1 U863 ( .A1(G95), .A2(n880), .ZN(n772) );
  NAND2_X1 U864 ( .A1(G107), .A2(n885), .ZN(n771) );
  NAND2_X1 U865 ( .A1(n772), .A2(n771), .ZN(n776) );
  NAND2_X1 U866 ( .A1(G131), .A2(n881), .ZN(n774) );
  NAND2_X1 U867 ( .A1(G119), .A2(n884), .ZN(n773) );
  NAND2_X1 U868 ( .A1(n774), .A2(n773), .ZN(n775) );
  OR2_X1 U869 ( .A1(n776), .A2(n775), .ZN(n873) );
  NAND2_X1 U870 ( .A1(G1991), .A2(n873), .ZN(n786) );
  XOR2_X1 U871 ( .A(KEYINPUT38), .B(KEYINPUT92), .Z(n778) );
  NAND2_X1 U872 ( .A1(G105), .A2(n880), .ZN(n777) );
  XNOR2_X1 U873 ( .A(n778), .B(n777), .ZN(n782) );
  NAND2_X1 U874 ( .A1(G141), .A2(n881), .ZN(n780) );
  NAND2_X1 U875 ( .A1(G117), .A2(n885), .ZN(n779) );
  NAND2_X1 U876 ( .A1(n780), .A2(n779), .ZN(n781) );
  NOR2_X1 U877 ( .A1(n782), .A2(n781), .ZN(n784) );
  NAND2_X1 U878 ( .A1(n884), .A2(G129), .ZN(n783) );
  NAND2_X1 U879 ( .A1(n784), .A2(n783), .ZN(n892) );
  NAND2_X1 U880 ( .A1(G1996), .A2(n892), .ZN(n785) );
  NAND2_X1 U881 ( .A1(n786), .A2(n785), .ZN(n921) );
  NAND2_X1 U882 ( .A1(n821), .A2(n921), .ZN(n814) );
  XOR2_X1 U883 ( .A(KEYINPUT93), .B(n814), .Z(n787) );
  NAND2_X1 U884 ( .A1(n818), .A2(n787), .ZN(n804) );
  OR2_X1 U885 ( .A1(n797), .A2(n804), .ZN(n788) );
  XNOR2_X1 U886 ( .A(G1986), .B(G290), .ZN(n975) );
  NAND2_X1 U887 ( .A1(n975), .A2(n821), .ZN(n798) );
  INV_X1 U888 ( .A(n798), .ZN(n806) );
  OR2_X1 U889 ( .A1(n788), .A2(n806), .ZN(n789) );
  NOR2_X1 U890 ( .A1(n790), .A2(n789), .ZN(n810) );
  NAND2_X1 U891 ( .A1(n792), .A2(n791), .ZN(n795) );
  NOR2_X1 U892 ( .A1(G2090), .A2(G303), .ZN(n793) );
  NAND2_X1 U893 ( .A1(G8), .A2(n793), .ZN(n794) );
  NAND2_X1 U894 ( .A1(n795), .A2(n794), .ZN(n801) );
  INV_X1 U895 ( .A(n804), .ZN(n796) );
  AND2_X1 U896 ( .A1(n797), .A2(n796), .ZN(n799) );
  AND2_X1 U897 ( .A1(n799), .A2(n798), .ZN(n800) );
  NAND2_X1 U898 ( .A1(n801), .A2(n800), .ZN(n808) );
  NAND2_X1 U899 ( .A1(n802), .A2(KEYINPUT33), .ZN(n803) );
  OR2_X1 U900 ( .A1(n804), .A2(n803), .ZN(n805) );
  OR2_X1 U901 ( .A1(n806), .A2(n805), .ZN(n807) );
  NAND2_X1 U902 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U903 ( .A1(n810), .A2(n809), .ZN(n824) );
  NAND2_X1 U904 ( .A1(n811), .A2(n896), .ZN(n918) );
  NOR2_X1 U905 ( .A1(G1991), .A2(n873), .ZN(n922) );
  NOR2_X1 U906 ( .A1(G1986), .A2(G290), .ZN(n812) );
  NOR2_X1 U907 ( .A1(n922), .A2(n812), .ZN(n813) );
  XNOR2_X1 U908 ( .A(n813), .B(KEYINPUT105), .ZN(n815) );
  NAND2_X1 U909 ( .A1(n815), .A2(n814), .ZN(n816) );
  OR2_X1 U910 ( .A1(n892), .A2(G1996), .ZN(n927) );
  NAND2_X1 U911 ( .A1(n816), .A2(n927), .ZN(n817) );
  XOR2_X1 U912 ( .A(KEYINPUT39), .B(n817), .Z(n819) );
  NAND2_X1 U913 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U914 ( .A1(n918), .A2(n820), .ZN(n822) );
  NAND2_X1 U915 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U916 ( .A1(n824), .A2(n823), .ZN(n826) );
  XNOR2_X1 U917 ( .A(KEYINPUT40), .B(KEYINPUT106), .ZN(n825) );
  XNOR2_X1 U918 ( .A(n826), .B(n825), .ZN(G329) );
  NAND2_X1 U919 ( .A1(n827), .A2(G2106), .ZN(n828) );
  XNOR2_X1 U920 ( .A(n828), .B(KEYINPUT108), .ZN(G217) );
  AND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n829) );
  NAND2_X1 U922 ( .A1(G661), .A2(n829), .ZN(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n830) );
  NAND2_X1 U924 ( .A1(n831), .A2(n830), .ZN(G188) );
  XNOR2_X1 U925 ( .A(G69), .B(KEYINPUT109), .ZN(G235) );
  XOR2_X1 U926 ( .A(KEYINPUT112), .B(G1981), .Z(n833) );
  XNOR2_X1 U927 ( .A(G1986), .B(G1961), .ZN(n832) );
  XNOR2_X1 U928 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U929 ( .A(n834), .B(KEYINPUT41), .Z(n836) );
  XNOR2_X1 U930 ( .A(G1996), .B(G1991), .ZN(n835) );
  XNOR2_X1 U931 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U932 ( .A(G1976), .B(G1971), .Z(n838) );
  XNOR2_X1 U933 ( .A(G1966), .B(G1956), .ZN(n837) );
  XNOR2_X1 U934 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U935 ( .A(n840), .B(n839), .Z(n842) );
  XNOR2_X1 U936 ( .A(KEYINPUT111), .B(G2474), .ZN(n841) );
  XNOR2_X1 U937 ( .A(n842), .B(n841), .ZN(G229) );
  XOR2_X1 U938 ( .A(G2096), .B(KEYINPUT43), .Z(n844) );
  XNOR2_X1 U939 ( .A(G2090), .B(KEYINPUT42), .ZN(n843) );
  XNOR2_X1 U940 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U941 ( .A(n845), .B(G2678), .Z(n847) );
  XNOR2_X1 U942 ( .A(G2067), .B(G2072), .ZN(n846) );
  XNOR2_X1 U943 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U944 ( .A(KEYINPUT110), .B(G2100), .Z(n849) );
  XNOR2_X1 U945 ( .A(G2084), .B(G2078), .ZN(n848) );
  XNOR2_X1 U946 ( .A(n849), .B(n848), .ZN(n850) );
  XNOR2_X1 U947 ( .A(n851), .B(n850), .ZN(G227) );
  XNOR2_X1 U948 ( .A(G286), .B(G301), .ZN(n852) );
  XNOR2_X1 U949 ( .A(n852), .B(n970), .ZN(n855) );
  XNOR2_X1 U950 ( .A(n969), .B(n853), .ZN(n854) );
  XNOR2_X1 U951 ( .A(n855), .B(n854), .ZN(n856) );
  NOR2_X1 U952 ( .A1(G37), .A2(n856), .ZN(G397) );
  NAND2_X1 U953 ( .A1(G124), .A2(n884), .ZN(n857) );
  XNOR2_X1 U954 ( .A(n857), .B(KEYINPUT44), .ZN(n860) );
  NAND2_X1 U955 ( .A1(G100), .A2(n880), .ZN(n858) );
  XOR2_X1 U956 ( .A(KEYINPUT113), .B(n858), .Z(n859) );
  NAND2_X1 U957 ( .A1(n860), .A2(n859), .ZN(n864) );
  NAND2_X1 U958 ( .A1(G136), .A2(n881), .ZN(n862) );
  NAND2_X1 U959 ( .A1(G112), .A2(n885), .ZN(n861) );
  NAND2_X1 U960 ( .A1(n862), .A2(n861), .ZN(n863) );
  NOR2_X1 U961 ( .A1(n864), .A2(n863), .ZN(G162) );
  NAND2_X1 U962 ( .A1(n884), .A2(G130), .ZN(n866) );
  NAND2_X1 U963 ( .A1(G118), .A2(n885), .ZN(n865) );
  NAND2_X1 U964 ( .A1(n866), .A2(n865), .ZN(n872) );
  NAND2_X1 U965 ( .A1(G106), .A2(n880), .ZN(n868) );
  NAND2_X1 U966 ( .A1(G142), .A2(n881), .ZN(n867) );
  NAND2_X1 U967 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U968 ( .A(KEYINPUT45), .B(n869), .Z(n870) );
  XNOR2_X1 U969 ( .A(KEYINPUT114), .B(n870), .ZN(n871) );
  NOR2_X1 U970 ( .A1(n872), .A2(n871), .ZN(n877) );
  XNOR2_X1 U971 ( .A(KEYINPUT115), .B(KEYINPUT48), .ZN(n875) );
  XNOR2_X1 U972 ( .A(n873), .B(KEYINPUT46), .ZN(n874) );
  XNOR2_X1 U973 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U974 ( .A(n877), .B(n876), .ZN(n879) );
  XNOR2_X1 U975 ( .A(n923), .B(G162), .ZN(n878) );
  XNOR2_X1 U976 ( .A(n879), .B(n878), .ZN(n891) );
  NAND2_X1 U977 ( .A1(G103), .A2(n880), .ZN(n883) );
  NAND2_X1 U978 ( .A1(G139), .A2(n881), .ZN(n882) );
  NAND2_X1 U979 ( .A1(n883), .A2(n882), .ZN(n890) );
  NAND2_X1 U980 ( .A1(n884), .A2(G127), .ZN(n887) );
  NAND2_X1 U981 ( .A1(G115), .A2(n885), .ZN(n886) );
  NAND2_X1 U982 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U983 ( .A(KEYINPUT47), .B(n888), .Z(n889) );
  NOR2_X1 U984 ( .A1(n890), .A2(n889), .ZN(n934) );
  XOR2_X1 U985 ( .A(n891), .B(n934), .Z(n894) );
  XOR2_X1 U986 ( .A(G164), .B(n892), .Z(n893) );
  XNOR2_X1 U987 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U988 ( .A(n895), .B(G160), .ZN(n897) );
  XNOR2_X1 U989 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U990 ( .A1(n898), .A2(G37), .ZN(n899) );
  XNOR2_X1 U991 ( .A(n899), .B(KEYINPUT116), .ZN(G395) );
  XOR2_X1 U992 ( .A(G2454), .B(G2430), .Z(n901) );
  XNOR2_X1 U993 ( .A(G2451), .B(G2446), .ZN(n900) );
  XNOR2_X1 U994 ( .A(n901), .B(n900), .ZN(n908) );
  XOR2_X1 U995 ( .A(G2443), .B(G2427), .Z(n903) );
  XNOR2_X1 U996 ( .A(G2438), .B(KEYINPUT107), .ZN(n902) );
  XNOR2_X1 U997 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U998 ( .A(n904), .B(G2435), .Z(n906) );
  XNOR2_X1 U999 ( .A(G1348), .B(G1341), .ZN(n905) );
  XNOR2_X1 U1000 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1001 ( .A(n908), .B(n907), .ZN(n909) );
  NAND2_X1 U1002 ( .A1(n909), .A2(G14), .ZN(n917) );
  NAND2_X1 U1003 ( .A1(n917), .A2(G319), .ZN(n912) );
  NOR2_X1 U1004 ( .A1(G229), .A2(G227), .ZN(n910) );
  XNOR2_X1 U1005 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NOR2_X1 U1006 ( .A1(n912), .A2(n911), .ZN(n914) );
  NOR2_X1 U1007 ( .A1(G397), .A2(G395), .ZN(n913) );
  NAND2_X1 U1008 ( .A1(n914), .A2(n913), .ZN(G225) );
  XNOR2_X1 U1009 ( .A(KEYINPUT117), .B(G225), .ZN(G308) );
  INV_X1 U1011 ( .A(G120), .ZN(G236) );
  INV_X1 U1012 ( .A(G96), .ZN(G221) );
  INV_X1 U1013 ( .A(G57), .ZN(G237) );
  NOR2_X1 U1014 ( .A1(n916), .A2(n915), .ZN(G325) );
  INV_X1 U1015 ( .A(G325), .ZN(G261) );
  INV_X1 U1016 ( .A(n917), .ZN(G401) );
  INV_X1 U1017 ( .A(n918), .ZN(n920) );
  NOR2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(n933) );
  NOR2_X1 U1019 ( .A1(n922), .A2(n921), .ZN(n924) );
  NAND2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(n931) );
  XOR2_X1 U1021 ( .A(KEYINPUT51), .B(KEYINPUT119), .Z(n929) );
  XNOR2_X1 U1022 ( .A(G2090), .B(G162), .ZN(n925) );
  XNOR2_X1 U1023 ( .A(n925), .B(KEYINPUT118), .ZN(n926) );
  NAND2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1025 ( .A(n929), .B(n928), .Z(n930) );
  NOR2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1027 ( .A1(n933), .A2(n932), .ZN(n941) );
  XOR2_X1 U1028 ( .A(G2072), .B(n934), .Z(n936) );
  XOR2_X1 U1029 ( .A(G164), .B(G2078), .Z(n935) );
  NOR2_X1 U1030 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1031 ( .A(KEYINPUT50), .B(n937), .ZN(n939) );
  XNOR2_X1 U1032 ( .A(G160), .B(G2084), .ZN(n938) );
  NAND2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1034 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1035 ( .A(KEYINPUT52), .B(n942), .ZN(n944) );
  INV_X1 U1036 ( .A(KEYINPUT55), .ZN(n943) );
  NAND2_X1 U1037 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1038 ( .A1(n945), .A2(G29), .ZN(n1025) );
  XNOR2_X1 U1039 ( .A(KEYINPUT121), .B(G1996), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(n946), .B(G32), .ZN(n957) );
  XOR2_X1 U1041 ( .A(G1991), .B(G25), .Z(n947) );
  NAND2_X1 U1042 ( .A1(n947), .A2(G28), .ZN(n955) );
  XOR2_X1 U1043 ( .A(n948), .B(G27), .Z(n953) );
  XNOR2_X1 U1044 ( .A(G2067), .B(G26), .ZN(n950) );
  XNOR2_X1 U1045 ( .A(G2072), .B(G33), .ZN(n949) );
  NOR2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1047 ( .A(n951), .B(KEYINPUT120), .ZN(n952) );
  NAND2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1050 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1051 ( .A(n958), .B(KEYINPUT53), .ZN(n961) );
  XOR2_X1 U1052 ( .A(G2084), .B(G34), .Z(n959) );
  XNOR2_X1 U1053 ( .A(KEYINPUT54), .B(n959), .ZN(n960) );
  NAND2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n963) );
  XNOR2_X1 U1055 ( .A(G35), .B(G2090), .ZN(n962) );
  NOR2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(KEYINPUT55), .B(n964), .ZN(n966) );
  INV_X1 U1058 ( .A(G29), .ZN(n965) );
  NAND2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1060 ( .A1(n967), .A2(G11), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(KEYINPUT122), .B(n968), .ZN(n1022) );
  XNOR2_X1 U1062 ( .A(G16), .B(KEYINPUT56), .ZN(n995) );
  XNOR2_X1 U1063 ( .A(n969), .B(G1348), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(n970), .B(G1341), .ZN(n971) );
  NOR2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n983) );
  XNOR2_X1 U1066 ( .A(G166), .B(G1971), .ZN(n977) );
  XOR2_X1 U1067 ( .A(n973), .B(G1956), .Z(n974) );
  NOR2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n981) );
  XNOR2_X1 U1070 ( .A(G171), .B(G1961), .ZN(n979) );
  NAND2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1073 ( .A1(n983), .A2(n982), .ZN(n986) );
  XNOR2_X1 U1074 ( .A(KEYINPUT125), .B(n984), .ZN(n985) );
  NOR2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n993) );
  XNOR2_X1 U1076 ( .A(G1966), .B(G168), .ZN(n988) );
  NAND2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1078 ( .A(n989), .B(KEYINPUT57), .ZN(n991) );
  XOR2_X1 U1079 ( .A(KEYINPUT124), .B(KEYINPUT123), .Z(n990) );
  XNOR2_X1 U1080 ( .A(n991), .B(n990), .ZN(n992) );
  NAND2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1082 ( .A1(n995), .A2(n994), .ZN(n1020) );
  INV_X1 U1083 ( .A(G16), .ZN(n1018) );
  XNOR2_X1 U1084 ( .A(G1348), .B(KEYINPUT59), .ZN(n996) );
  XNOR2_X1 U1085 ( .A(n996), .B(G4), .ZN(n1000) );
  XNOR2_X1 U1086 ( .A(G1956), .B(G20), .ZN(n998) );
  XNOR2_X1 U1087 ( .A(G6), .B(G1981), .ZN(n997) );
  NOR2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1003) );
  XNOR2_X1 U1090 ( .A(G19), .B(G1341), .ZN(n1001) );
  XNOR2_X1 U1091 ( .A(KEYINPUT126), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(KEYINPUT60), .B(n1004), .ZN(n1008) );
  XNOR2_X1 U1094 ( .A(G1966), .B(G21), .ZN(n1006) );
  XNOR2_X1 U1095 ( .A(G5), .B(G1961), .ZN(n1005) );
  NOR2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1015) );
  XNOR2_X1 U1098 ( .A(G1971), .B(G22), .ZN(n1010) );
  XNOR2_X1 U1099 ( .A(G23), .B(G1976), .ZN(n1009) );
  NOR2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XOR2_X1 U1101 ( .A(G1986), .B(G24), .Z(n1011) );
  NAND2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1103 ( .A(KEYINPUT58), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1105 ( .A(KEYINPUT61), .B(n1016), .ZN(n1017) );
  NAND2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1109 ( .A(KEYINPUT127), .B(n1023), .Z(n1024) );
  NAND2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1111 ( .A(KEYINPUT62), .B(n1026), .Z(G311) );
  INV_X1 U1112 ( .A(G311), .ZN(G150) );
endmodule

