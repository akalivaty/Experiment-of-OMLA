//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 1 0 0 0 0 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 0 0 0 0 1 1 1 1 1 1 0 1 0 0 0 0 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936;
  XNOR2_X1  g000(.A(G116), .B(G119), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT2), .B(G113), .ZN(new_n189));
  OR2_X1    g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n189), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G101), .ZN(new_n193));
  OR2_X1    g007(.A1(KEYINPUT3), .A2(G107), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT78), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G104), .ZN(new_n196));
  INV_X1    g010(.A(G104), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(KEYINPUT78), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n194), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(KEYINPUT3), .A2(G107), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  NOR2_X1   g015(.A1(KEYINPUT3), .A2(G107), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n201), .B1(G104), .B2(new_n202), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n193), .B1(new_n199), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT4), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n192), .A2(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n199), .A2(new_n203), .A3(new_n193), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT79), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n208), .B1(new_n204), .B2(new_n209), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n200), .B1(new_n194), .B2(new_n197), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n197), .A2(KEYINPUT78), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n195), .A2(G104), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n202), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n209), .B(G101), .C1(new_n211), .C2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT4), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT80), .B1(new_n210), .B2(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n205), .B1(new_n204), .B2(new_n209), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT80), .ZN(new_n219));
  OAI21_X1  g033(.A(G101), .B1(new_n211), .B2(new_n214), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT79), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n218), .A2(new_n219), .A3(new_n208), .A4(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n207), .B1(new_n217), .B2(new_n222), .ZN(new_n223));
  XOR2_X1   g037(.A(G110), .B(G122), .Z(new_n224));
  NAND2_X1  g038(.A1(G104), .A2(G107), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT78), .B(G104), .ZN(new_n226));
  OAI211_X1 g040(.A(G101), .B(new_n225), .C1(new_n226), .C2(G107), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT81), .ZN(new_n228));
  INV_X1    g042(.A(G107), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n229), .B1(new_n196), .B2(new_n198), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT81), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n230), .A2(new_n231), .A3(G101), .A4(new_n225), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n228), .A2(new_n208), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT5), .ZN(new_n234));
  INV_X1    g048(.A(G119), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(new_n235), .A3(G116), .ZN(new_n236));
  OAI211_X1 g050(.A(G113), .B(new_n236), .C1(new_n188), .C2(new_n234), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(new_n190), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n233), .A2(new_n238), .ZN(new_n239));
  OR3_X1    g053(.A1(new_n223), .A2(new_n224), .A3(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n224), .B1(new_n223), .B2(new_n239), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n240), .A2(KEYINPUT6), .A3(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(G143), .B(G146), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT0), .ZN(new_n244));
  INV_X1    g058(.A(G128), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  XOR2_X1   g060(.A(KEYINPUT0), .B(G128), .Z(new_n247));
  OAI21_X1  g061(.A(new_n246), .B1(new_n243), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G125), .ZN(new_n249));
  OR3_X1    g063(.A1(new_n248), .A2(KEYINPUT88), .A3(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G146), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G143), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(G128), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n245), .A2(KEYINPUT1), .ZN(new_n254));
  INV_X1    g068(.A(G143), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G146), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n254), .A2(new_n252), .A3(new_n256), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT66), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n254), .A2(new_n252), .A3(new_n256), .A4(KEYINPUT66), .ZN(new_n261));
  AOI211_X1 g075(.A(new_n253), .B(new_n257), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n249), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT88), .B1(new_n248), .B2(new_n249), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n250), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT90), .ZN(new_n266));
  INV_X1    g080(.A(G953), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G224), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n268), .B(KEYINPUT89), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT90), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n250), .A2(new_n263), .A3(new_n270), .A4(new_n264), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n266), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n269), .B1(new_n266), .B2(new_n271), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n275), .B(new_n224), .C1(new_n223), .C2(new_n239), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n242), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G902), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n269), .A2(KEYINPUT7), .ZN(new_n279));
  XOR2_X1   g093(.A(new_n265), .B(new_n279), .Z(new_n280));
  XOR2_X1   g094(.A(new_n233), .B(new_n238), .Z(new_n281));
  XNOR2_X1  g095(.A(new_n224), .B(KEYINPUT8), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n280), .B(new_n240), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n277), .A2(new_n278), .A3(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(G210), .B1(G237), .B2(G902), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n277), .A2(new_n278), .A3(new_n285), .A4(new_n283), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(G214), .B1(G237), .B2(G902), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  XOR2_X1   g105(.A(KEYINPUT9), .B(G234), .Z(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(G221), .B1(new_n293), .B2(G902), .ZN(new_n294));
  XOR2_X1   g108(.A(new_n294), .B(KEYINPUT77), .Z(new_n295));
  OAI21_X1  g109(.A(KEYINPUT82), .B1(new_n233), .B2(new_n262), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT10), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT10), .ZN(new_n298));
  OAI211_X1 g112(.A(KEYINPUT82), .B(new_n298), .C1(new_n233), .C2(new_n262), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n206), .A2(new_n248), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n301), .B1(new_n217), .B2(new_n222), .ZN(new_n302));
  INV_X1    g116(.A(G131), .ZN(new_n303));
  INV_X1    g117(.A(G137), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT64), .ZN(new_n305));
  INV_X1    g119(.A(G134), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(KEYINPUT64), .A2(G134), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n304), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT11), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n307), .A2(new_n304), .A3(new_n308), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(KEYINPUT11), .A2(G134), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT65), .B1(new_n313), .B2(G137), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT65), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n315), .A2(new_n304), .A3(KEYINPUT11), .A4(G134), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n303), .B1(new_n312), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n311), .A2(new_n310), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n307), .A2(new_n308), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G137), .ZN(new_n321));
  AND4_X1   g135(.A1(new_n303), .A2(new_n317), .A3(new_n319), .A4(new_n321), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NOR3_X1   g138(.A1(new_n300), .A2(new_n302), .A3(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(G110), .B(G140), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n267), .A2(G227), .ZN(new_n327));
  XOR2_X1   g141(.A(new_n326), .B(new_n327), .Z(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT85), .B1(new_n325), .B2(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n233), .B(new_n262), .ZN(new_n331));
  AND3_X1   g145(.A1(new_n331), .A2(KEYINPUT12), .A3(new_n324), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT12), .B1(new_n331), .B2(new_n324), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n301), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n211), .A2(new_n214), .A3(G101), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n337), .B1(KEYINPUT79), .B2(new_n220), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n219), .B1(new_n338), .B2(new_n218), .ZN(new_n339));
  NOR3_X1   g153(.A1(new_n210), .A2(new_n216), .A3(KEYINPUT80), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n336), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n341), .A2(new_n323), .A3(new_n297), .A4(new_n299), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT85), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n342), .A2(new_n343), .A3(new_n328), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n330), .A2(new_n335), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT86), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n324), .B1(new_n300), .B2(new_n302), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n342), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n346), .B1(new_n348), .B2(new_n329), .ZN(new_n349));
  AOI211_X1 g163(.A(KEYINPUT86), .B(new_n328), .C1(new_n347), .C2(new_n342), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n345), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G469), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(new_n352), .A3(new_n278), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT83), .B1(new_n325), .B2(new_n329), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT83), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n342), .A2(new_n355), .A3(new_n328), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n354), .A2(new_n347), .A3(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n329), .B1(new_n334), .B2(new_n325), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(G469), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(G469), .A2(G902), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(KEYINPUT84), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n353), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(KEYINPUT84), .B1(new_n359), .B2(new_n360), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n295), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT87), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI211_X1 g180(.A(KEYINPUT87), .B(new_n295), .C1(new_n362), .C2(new_n363), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n291), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G140), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G125), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT75), .B1(new_n370), .B2(KEYINPUT16), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT75), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT16), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n372), .A2(new_n373), .A3(new_n369), .A4(G125), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n249), .A2(G140), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n371), .B(new_n374), .C1(new_n376), .C2(new_n373), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n377), .A2(new_n251), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT76), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n377), .A2(new_n251), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  XOR2_X1   g196(.A(KEYINPUT24), .B(G110), .Z(new_n383));
  XNOR2_X1  g197(.A(G119), .B(G128), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NOR3_X1   g199(.A1(new_n235), .A2(KEYINPUT23), .A3(G128), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n386), .B1(new_n384), .B2(KEYINPUT23), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G110), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n377), .A2(new_n379), .A3(new_n251), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n382), .A2(new_n385), .A3(new_n388), .A4(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n376), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n378), .B1(new_n251), .B2(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n387), .A2(G110), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n383), .A2(new_n384), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n267), .A2(G221), .A3(G234), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n397), .B(KEYINPUT22), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n398), .B(G137), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n396), .B(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n278), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT25), .ZN(new_n402));
  INV_X1    g216(.A(G217), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n403), .B1(G234), .B2(new_n278), .ZN(new_n404));
  XOR2_X1   g218(.A(new_n404), .B(KEYINPUT74), .Z(new_n405));
  INV_X1    g219(.A(KEYINPUT25), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n400), .A2(new_n406), .A3(new_n278), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n402), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  OR2_X1    g222(.A1(new_n401), .A2(new_n404), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(G472), .A2(G902), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n248), .B1(new_n318), .B2(new_n322), .ZN(new_n412));
  INV_X1    g226(.A(new_n192), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n260), .A2(new_n261), .ZN(new_n414));
  INV_X1    g228(.A(new_n253), .ZN(new_n415));
  INV_X1    g229(.A(new_n257), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n312), .A2(new_n303), .A3(new_n317), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n311), .B1(G134), .B2(new_n304), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G131), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n417), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n412), .A2(new_n413), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT70), .ZN(new_n423));
  XNOR2_X1  g237(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(G237), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n426), .A2(new_n267), .A3(G210), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n427), .B(KEYINPUT69), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT26), .B(G101), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n428), .A2(new_n429), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n425), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n432), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(new_n424), .A3(new_n430), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n422), .A2(new_n423), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n423), .B1(new_n422), .B2(new_n436), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n421), .ZN(new_n440));
  INV_X1    g254(.A(new_n248), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n317), .A2(new_n319), .A3(new_n321), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G131), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n441), .B1(new_n443), .B2(new_n418), .ZN(new_n444));
  OAI211_X1 g258(.A(KEYINPUT67), .B(KEYINPUT30), .C1(new_n440), .C2(new_n444), .ZN(new_n445));
  OR2_X1    g259(.A1(KEYINPUT67), .A2(KEYINPUT30), .ZN(new_n446));
  NAND2_X1  g260(.A1(KEYINPUT67), .A2(KEYINPUT30), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n412), .A2(new_n446), .A3(new_n421), .A4(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n413), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  NOR3_X1   g263(.A1(new_n439), .A2(KEYINPUT71), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT71), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n422), .A2(new_n436), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT70), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n422), .A2(new_n423), .A3(new_n436), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n445), .A2(new_n448), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n192), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n451), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(KEYINPUT31), .B1(new_n450), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n439), .A2(new_n449), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT31), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT28), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n192), .B1(new_n440), .B2(new_n444), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n462), .B1(new_n463), .B2(new_n422), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n422), .A2(new_n462), .ZN(new_n465));
  OR2_X1    g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n436), .ZN(new_n467));
  AOI22_X1  g281(.A1(new_n460), .A2(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(KEYINPUT72), .B1(new_n459), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(KEYINPUT71), .B1(new_n439), .B2(new_n449), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n455), .A2(new_n457), .A3(new_n451), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n461), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT72), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n467), .B1(new_n464), .B2(new_n465), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n455), .A2(new_n457), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n474), .B1(new_n475), .B2(KEYINPUT31), .ZN(new_n476));
  NOR3_X1   g290(.A1(new_n472), .A2(new_n473), .A3(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n411), .B1(new_n469), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(KEYINPUT32), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n473), .B1(new_n472), .B2(new_n476), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n459), .A2(KEYINPUT72), .A3(new_n468), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT32), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n483), .A3(new_n411), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n479), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n457), .A2(new_n422), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n467), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(KEYINPUT73), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT29), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n489), .B1(new_n466), .B2(new_n467), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n278), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  NOR3_X1   g305(.A1(new_n466), .A2(new_n489), .A3(new_n467), .ZN(new_n492));
  OAI21_X1  g306(.A(G472), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n410), .B1(new_n485), .B2(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(G113), .B(G122), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(new_n197), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n426), .A2(new_n267), .A3(G214), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(G143), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n498), .A2(new_n303), .ZN(new_n499));
  AOI22_X1  g313(.A1(new_n382), .A2(new_n389), .B1(KEYINPUT17), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n303), .ZN(new_n501));
  OR2_X1    g315(.A1(new_n501), .A2(KEYINPUT91), .ZN(new_n502));
  OR2_X1    g316(.A1(new_n498), .A2(new_n303), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(KEYINPUT91), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n500), .B1(KEYINPUT17), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT18), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n498), .B1(new_n507), .B2(new_n303), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n376), .B(G146), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n508), .B(new_n509), .C1(new_n503), .C2(new_n507), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n496), .B1(new_n506), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT94), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n506), .A2(new_n496), .A3(new_n510), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT94), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n512), .B(new_n278), .C1(new_n515), .C2(new_n511), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(G475), .ZN(new_n517));
  XOR2_X1   g331(.A(new_n376), .B(KEYINPUT19), .Z(new_n518));
  AOI21_X1  g332(.A(new_n378), .B1(new_n251), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n505), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n496), .B1(new_n520), .B2(new_n510), .ZN(new_n521));
  OR2_X1    g335(.A1(new_n521), .A2(KEYINPUT92), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(KEYINPUT92), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n522), .A2(new_n513), .A3(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(G475), .A2(G902), .ZN(new_n525));
  XOR2_X1   g339(.A(new_n525), .B(KEYINPUT93), .Z(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT20), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n524), .A2(KEYINPUT20), .A3(new_n526), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n517), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(G128), .B(G143), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n306), .B1(new_n533), .B2(KEYINPUT13), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n255), .A2(G128), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n534), .B1(KEYINPUT13), .B2(new_n535), .ZN(new_n536));
  OR2_X1    g350(.A1(new_n536), .A2(KEYINPUT95), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n320), .A2(new_n533), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  XOR2_X1   g353(.A(G116), .B(G122), .Z(new_n540));
  OR2_X1    g354(.A1(new_n540), .A2(G107), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(G107), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n539), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n536), .A2(KEYINPUT95), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n537), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(G116), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(KEYINPUT14), .A3(G122), .ZN(new_n547));
  OAI211_X1 g361(.A(G107), .B(new_n547), .C1(new_n540), .C2(KEYINPUT14), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n320), .A2(new_n533), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n548), .B(new_n541), .C1(new_n539), .C2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n293), .A2(new_n403), .A3(G953), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n552), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n545), .A2(new_n550), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n553), .A2(new_n278), .A3(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(G478), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n557), .A2(KEYINPUT15), .ZN(new_n558));
  XOR2_X1   g372(.A(new_n556), .B(new_n558), .Z(new_n559));
  NAND2_X1  g373(.A1(new_n532), .A2(new_n559), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n267), .A2(G952), .ZN(new_n561));
  NAND2_X1  g375(.A1(G234), .A2(G237), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  XOR2_X1   g378(.A(KEYINPUT21), .B(G898), .Z(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n562), .A2(G902), .A3(G953), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n564), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n560), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n368), .A2(new_n494), .A3(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(G101), .ZN(G3));
  NAND2_X1  g386(.A1(new_n366), .A2(new_n367), .ZN(new_n573));
  INV_X1    g387(.A(new_n410), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n278), .B1(new_n469), .B2(new_n477), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(G472), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n576), .A2(new_n478), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n573), .A2(new_n574), .A3(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT96), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n551), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n552), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n551), .A2(new_n579), .A3(new_n554), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n581), .A2(KEYINPUT33), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT97), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT97), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n553), .A2(new_n555), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n585), .B1(new_n586), .B2(KEYINPUT33), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n584), .B1(new_n583), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n588), .A2(G478), .A3(new_n278), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n556), .A2(new_n557), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n531), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n592), .A2(new_n291), .A3(new_n569), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n578), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT34), .B(G104), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(G6));
  OR2_X1    g411(.A1(new_n531), .A2(new_n559), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n598), .A2(new_n291), .A3(new_n569), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n578), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT35), .B(G107), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G9));
  INV_X1    g417(.A(new_n399), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n604), .A2(KEYINPUT36), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n396), .B(new_n605), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n606), .B(new_n278), .C1(new_n403), .C2(G234), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n408), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n368), .A2(new_n570), .A3(new_n577), .A4(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(KEYINPUT37), .ZN(new_n610));
  XOR2_X1   g424(.A(new_n610), .B(G110), .Z(G12));
  INV_X1    g425(.A(new_n608), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n612), .B1(new_n485), .B2(new_n493), .ZN(new_n613));
  INV_X1    g427(.A(new_n291), .ZN(new_n614));
  OR2_X1    g428(.A1(new_n567), .A2(G900), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n563), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n598), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n613), .A2(new_n573), .A3(new_n614), .A4(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G128), .ZN(G30));
  XNOR2_X1  g434(.A(new_n616), .B(KEYINPUT39), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n573), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT98), .B(KEYINPUT40), .Z(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n289), .B(KEYINPUT38), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n450), .A2(new_n458), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n436), .B1(new_n463), .B2(new_n422), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n278), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(G472), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n485), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n633), .A2(new_n608), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n532), .A2(new_n559), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n636), .B1(new_n622), .B2(new_n623), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n627), .A2(new_n290), .A3(new_n634), .A4(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G143), .ZN(G45));
  AOI21_X1  g453(.A(new_n483), .B1(new_n482), .B2(new_n411), .ZN(new_n640));
  INV_X1    g454(.A(new_n411), .ZN(new_n641));
  AOI211_X1 g455(.A(KEYINPUT32), .B(new_n641), .C1(new_n480), .C2(new_n481), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n493), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n591), .A2(new_n531), .A3(new_n616), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n644), .A2(new_n291), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n573), .A2(new_n643), .A3(new_n608), .A4(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT99), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G146), .ZN(G48));
  INV_X1    g462(.A(new_n294), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n351), .A2(new_n278), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(G469), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n651), .A2(KEYINPUT100), .A3(new_n353), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT100), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n650), .A2(new_n653), .A3(G469), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n649), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n643), .A2(new_n574), .A3(new_n593), .A4(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT41), .B(G113), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G15));
  NAND4_X1  g472(.A1(new_n643), .A2(new_n599), .A3(new_n574), .A4(new_n655), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G116), .ZN(G18));
  NAND3_X1  g474(.A1(new_n643), .A2(new_n570), .A3(new_n608), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n655), .A2(new_n614), .ZN(new_n662));
  OAI21_X1  g476(.A(KEYINPUT101), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT101), .ZN(new_n664));
  AOI211_X1 g478(.A(new_n649), .B(new_n291), .C1(new_n652), .C2(new_n654), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n613), .A2(new_n664), .A3(new_n570), .A4(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G119), .ZN(G21));
  AOI21_X1  g482(.A(new_n641), .B1(new_n459), .B2(new_n468), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(G902), .B1(new_n480), .B2(new_n481), .ZN(new_n671));
  INV_X1    g485(.A(G472), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n574), .B(new_n670), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n291), .A2(new_n569), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n674), .A2(new_n655), .A3(new_n675), .A4(new_n635), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G122), .ZN(G24));
  INV_X1    g491(.A(new_n644), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n669), .B1(new_n575), .B2(G472), .ZN(new_n679));
  AOI21_X1  g493(.A(KEYINPUT102), .B1(new_n679), .B2(new_n608), .ZN(new_n680));
  OAI211_X1 g494(.A(new_n608), .B(new_n670), .C1(new_n671), .C2(new_n672), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT102), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n678), .B(new_n665), .C1(new_n680), .C2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G125), .ZN(G27));
  NAND2_X1  g499(.A1(new_n494), .A2(KEYINPUT106), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n643), .A2(new_n574), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT105), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n287), .A2(new_n290), .A3(new_n288), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n360), .B(KEYINPUT103), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n359), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n649), .B1(new_n694), .B2(new_n353), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n692), .B1(new_n695), .B2(KEYINPUT104), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT104), .ZN(new_n697));
  AOI211_X1 g511(.A(new_n697), .B(new_n649), .C1(new_n694), .C2(new_n353), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n690), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  AND3_X1   g513(.A1(new_n351), .A2(new_n352), .A3(new_n278), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n359), .A2(new_n693), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n294), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n697), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n695), .A2(KEYINPUT104), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n703), .A2(KEYINPUT105), .A3(new_n704), .A4(new_n692), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n699), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n686), .A2(new_n689), .A3(new_n706), .A4(new_n678), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n687), .B1(new_n699), .B2(new_n705), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n644), .A2(KEYINPUT42), .ZN(new_n709));
  AOI22_X1  g523(.A1(new_n707), .A2(KEYINPUT42), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G131), .ZN(G33));
  AOI21_X1  g525(.A(new_n691), .B1(new_n702), .B2(new_n697), .ZN(new_n712));
  AOI21_X1  g526(.A(KEYINPUT105), .B1(new_n712), .B2(new_n704), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n696), .A2(new_n690), .A3(new_n698), .ZN(new_n714));
  OAI211_X1 g528(.A(new_n494), .B(new_n618), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G134), .ZN(G36));
  NOR2_X1   g530(.A1(new_n577), .A2(new_n612), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n532), .A2(new_n718), .A3(new_n591), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n531), .B(KEYINPUT108), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n720), .A2(new_n591), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n717), .B(new_n719), .C1(new_n718), .C2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n692), .B1(new_n723), .B2(KEYINPUT44), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n357), .A2(new_n358), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(KEYINPUT45), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(G469), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(KEYINPUT46), .A3(new_n693), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n353), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT107), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n728), .A2(KEYINPUT107), .A3(new_n353), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n727), .A2(new_n693), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n731), .B(new_n732), .C1(KEYINPUT46), .C2(new_n733), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n734), .A2(new_n294), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n621), .ZN(new_n736));
  AOI211_X1 g550(.A(new_n724), .B(new_n736), .C1(KEYINPUT44), .C2(new_n723), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(new_n304), .ZN(G39));
  NAND2_X1  g552(.A1(new_n692), .A2(new_n616), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n734), .A2(new_n294), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT47), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n734), .A2(KEYINPUT47), .A3(new_n294), .ZN(new_n743));
  AOI211_X1 g557(.A(new_n643), .B(new_n739), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n592), .A2(new_n574), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G140), .ZN(G42));
  AND2_X1   g561(.A1(new_n655), .A2(new_n692), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n633), .A2(new_n748), .A3(new_n574), .A4(new_n564), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n561), .B1(new_n749), .B2(new_n592), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n564), .B(new_n719), .C1(new_n721), .C2(new_n718), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n751), .A2(new_n673), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n750), .B1(new_n665), .B2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(KEYINPUT120), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n652), .A2(new_n654), .ZN(new_n755));
  INV_X1    g569(.A(new_n295), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n742), .A2(new_n743), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT119), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n751), .A2(new_n673), .A3(new_n691), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT119), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n742), .A2(new_n761), .A3(new_n743), .A4(new_n757), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n759), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n290), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n655), .A2(KEYINPUT116), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(KEYINPUT116), .B1(new_n655), .B2(new_n764), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n625), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n752), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT50), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n749), .A2(new_n531), .A3(new_n591), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT117), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  INV_X1    g588(.A(new_n748), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n681), .A2(new_n682), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n576), .A2(KEYINPUT102), .A3(new_n608), .A4(new_n670), .ZN(new_n777));
  AOI211_X1 g591(.A(new_n775), .B(new_n751), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n773), .A2(new_n774), .A3(new_n778), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n763), .B(new_n770), .C1(KEYINPUT118), .C2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT51), .ZN(new_n781));
  XOR2_X1   g595(.A(new_n757), .B(KEYINPUT115), .Z(new_n782));
  NAND3_X1  g596(.A1(new_n742), .A2(new_n743), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(KEYINPUT51), .B1(new_n783), .B2(new_n760), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n784), .A2(new_n770), .ZN(new_n785));
  AND2_X1   g599(.A1(KEYINPUT118), .A2(KEYINPUT51), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n779), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n754), .B1(new_n781), .B2(new_n787), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n684), .A2(new_n646), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n616), .A2(KEYINPUT111), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n616), .A2(KEYINPUT111), .ZN(new_n791));
  AND4_X1   g605(.A1(new_n614), .A2(new_n635), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n792), .A2(new_n632), .A3(new_n612), .A4(new_n695), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n789), .A2(KEYINPUT52), .A3(new_n619), .A4(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n619), .A2(new_n684), .A3(new_n793), .A4(new_n646), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n644), .B1(new_n777), .B2(new_n776), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n706), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n739), .A2(new_n560), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n613), .A2(new_n573), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n715), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT110), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n715), .A2(new_n800), .A3(KEYINPUT110), .A4(new_n802), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n798), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n531), .A2(new_n559), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n675), .A2(KEYINPUT109), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT109), .B1(new_n675), .B2(new_n809), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n594), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n812), .A2(new_n574), .A3(new_n573), .A4(new_n577), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n813), .A2(new_n571), .A3(new_n609), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n659), .A2(new_n656), .A3(new_n676), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n667), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n814), .A2(new_n816), .A3(new_n710), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n818));
  OR3_X1    g632(.A1(new_n808), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT112), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n818), .B1(new_n808), .B2(new_n817), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  OAI211_X1 g636(.A(KEYINPUT112), .B(new_n818), .C1(new_n808), .C2(new_n817), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n822), .A2(KEYINPUT54), .A3(new_n823), .ZN(new_n824));
  AND4_X1   g638(.A1(KEYINPUT53), .A2(new_n813), .A3(new_n571), .A4(new_n609), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n798), .A2(new_n807), .A3(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n667), .A2(KEYINPUT113), .A3(new_n815), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT113), .B1(new_n667), .B2(new_n815), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n710), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI211_X1 g645(.A(KEYINPUT114), .B(new_n710), .C1(new_n827), .C2(new_n828), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n826), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n833), .A2(new_n834), .A3(new_n821), .ZN(new_n835));
  INV_X1    g649(.A(new_n751), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n836), .A2(new_n689), .A3(new_n686), .A4(new_n748), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(KEYINPUT48), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n788), .A2(new_n824), .A3(new_n835), .A4(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n839), .B1(G952), .B2(G953), .ZN(new_n840));
  XOR2_X1   g654(.A(new_n755), .B(KEYINPUT49), .Z(new_n841));
  NOR4_X1   g655(.A1(new_n841), .A2(new_n410), .A3(new_n756), .A4(new_n764), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n842), .A2(new_n633), .A3(new_n626), .A4(new_n721), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n840), .A2(new_n843), .ZN(G75));
  XNOR2_X1  g658(.A(new_n274), .B(KEYINPUT55), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n242), .A2(new_n276), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(KEYINPUT121), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n278), .B1(new_n833), .B2(new_n821), .ZN(new_n848));
  AOI211_X1 g662(.A(KEYINPUT56), .B(new_n847), .C1(new_n848), .C2(G210), .ZN(new_n849));
  INV_X1    g663(.A(new_n847), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n833), .A2(new_n821), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n851), .A2(G210), .A3(G902), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT56), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n850), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n845), .B1(new_n849), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n267), .A2(G952), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(G210), .ZN(new_n858));
  AOI211_X1 g672(.A(new_n858), .B(new_n278), .C1(new_n833), .C2(new_n821), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n847), .B1(new_n859), .B2(KEYINPUT56), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n852), .A2(new_n853), .A3(new_n850), .ZN(new_n861));
  INV_X1    g675(.A(new_n845), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n855), .A2(new_n857), .A3(new_n863), .ZN(G51));
  NAND2_X1  g678(.A1(new_n851), .A2(KEYINPUT54), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n865), .A2(KEYINPUT122), .A3(new_n835), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT122), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n851), .A2(new_n867), .A3(KEYINPUT54), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n693), .B(KEYINPUT57), .Z(new_n869));
  NAND3_X1  g683(.A1(new_n866), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n351), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n848), .A2(G469), .A3(new_n726), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n856), .B1(new_n871), .B2(new_n872), .ZN(G54));
  INV_X1    g687(.A(new_n848), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT123), .B1(KEYINPUT58), .B2(G475), .ZN(new_n875));
  AND3_X1   g689(.A1(KEYINPUT123), .A2(KEYINPUT58), .A3(G475), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n877), .A2(new_n524), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n877), .A2(new_n524), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n878), .A2(new_n879), .A3(new_n856), .ZN(G60));
  NAND2_X1  g694(.A1(G478), .A2(G902), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(KEYINPUT59), .Z(new_n882));
  AOI21_X1  g696(.A(new_n882), .B1(new_n824), .B2(new_n835), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n857), .B1(new_n883), .B2(new_n588), .ZN(new_n884));
  INV_X1    g698(.A(new_n882), .ZN(new_n885));
  AND4_X1   g699(.A1(new_n588), .A2(new_n866), .A3(new_n868), .A4(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n884), .A2(new_n886), .ZN(G63));
  NAND2_X1  g701(.A1(G217), .A2(G902), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n888), .B(KEYINPUT60), .Z(new_n889));
  XOR2_X1   g703(.A(new_n606), .B(KEYINPUT124), .Z(new_n890));
  NAND3_X1  g704(.A1(new_n851), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n851), .A2(new_n889), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n857), .B(new_n891), .C1(new_n892), .C2(new_n400), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT61), .B1(new_n891), .B2(KEYINPUT125), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n893), .B(new_n894), .ZN(G66));
  AOI21_X1  g709(.A(new_n267), .B1(new_n565), .B2(G224), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n814), .A2(new_n816), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT126), .Z(new_n898));
  AOI21_X1  g712(.A(new_n896), .B1(new_n898), .B2(new_n267), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n850), .B1(G898), .B2(new_n267), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n899), .B(new_n900), .Z(G69));
  XNOR2_X1  g715(.A(new_n456), .B(new_n518), .ZN(new_n902));
  NAND2_X1  g716(.A1(G900), .A2(G953), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n737), .B1(new_n744), .B2(new_n745), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n789), .A2(new_n619), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  AND4_X1   g720(.A1(new_n621), .A2(new_n735), .A3(new_n689), .A4(new_n686), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n636), .A2(new_n291), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n710), .A2(new_n715), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n904), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n902), .B(new_n903), .C1(new_n911), .C2(G953), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n638), .A2(new_n905), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(KEYINPUT62), .Z(new_n914));
  NAND2_X1  g728(.A1(new_n598), .A2(new_n592), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n622), .A2(new_n494), .A3(new_n692), .A4(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n914), .A2(new_n904), .A3(new_n916), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n917), .A2(new_n267), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n912), .B1(new_n918), .B2(new_n902), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n267), .B1(G227), .B2(G900), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n920), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n922), .B(new_n912), .C1(new_n918), .C2(new_n902), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n921), .A2(new_n923), .ZN(G72));
  XOR2_X1   g738(.A(KEYINPUT127), .B(KEYINPUT63), .Z(new_n925));
  NOR2_X1   g739(.A1(new_n672), .A2(new_n278), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n928), .B1(new_n917), .B2(new_n898), .ZN(new_n929));
  INV_X1    g743(.A(new_n486), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n930), .A2(new_n467), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n856), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n928), .B1(new_n911), .B2(new_n898), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n933), .A2(new_n467), .A3(new_n930), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n488), .A2(new_n628), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n822), .A2(new_n823), .A3(new_n928), .A4(new_n935), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n932), .A2(new_n934), .A3(new_n936), .ZN(G57));
endmodule


