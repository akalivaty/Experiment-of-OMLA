//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 0 0 1 1 0 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1218,
    new_n1219, new_n1220, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(new_n203), .A2(G50), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT65), .Z(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G1), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n211), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G58), .A2(G232), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n219));
  AND4_X1   g0019(.A1(new_n216), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(KEYINPUT66), .B(G244), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(G77), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n215), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT1), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n213), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(new_n215), .ZN(new_n226));
  OR3_X1    g0026(.A1(new_n226), .A2(KEYINPUT64), .A3(G13), .ZN(new_n227));
  OAI21_X1  g0027(.A(KEYINPUT64), .B1(new_n226), .B2(G13), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n229), .B(G250), .C1(G257), .C2(G264), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT0), .Z(new_n231));
  AOI211_X1 g0031(.A(new_n225), .B(new_n231), .C1(new_n224), .C2(new_n223), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  INV_X1    g0043(.A(G50), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(G68), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n202), .A2(G50), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n243), .B(new_n249), .ZN(G351));
  NAND3_X1  g0050(.A1(new_n214), .A2(G13), .A3(G20), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT68), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g0053(.A1(new_n214), .A2(KEYINPUT68), .A3(G13), .A4(G20), .ZN(new_n254));
  AND2_X1   g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G116), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n253), .A2(new_n254), .ZN(new_n258));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n210), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n214), .A2(G33), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n258), .A2(new_n261), .A3(G116), .A4(new_n262), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n259), .A2(new_n210), .B1(G20), .B2(new_n256), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G283), .ZN(new_n265));
  INV_X1    g0065(.A(G97), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n265), .B(new_n211), .C1(G33), .C2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(KEYINPUT20), .B1(new_n264), .B2(new_n267), .ZN(new_n268));
  AND3_X1   g0068(.A1(new_n264), .A2(KEYINPUT20), .A3(new_n267), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n257), .B(new_n263), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT5), .B(G41), .ZN(new_n271));
  INV_X1    g0071(.A(G45), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G1), .ZN(new_n273));
  INV_X1    g0073(.A(new_n210), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n271), .A2(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n214), .A2(G45), .ZN(new_n277));
  NOR2_X1   g0077(.A1(KEYINPUT5), .A2(G41), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(KEYINPUT5), .A2(G41), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n277), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G274), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n282), .B1(new_n274), .B2(new_n275), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n276), .A2(G270), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT3), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(G33), .ZN(new_n286));
  INV_X1    g0086(.A(G33), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(KEYINPUT3), .ZN(new_n288));
  OAI21_X1  g0088(.A(G303), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(KEYINPUT3), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n285), .A2(G33), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n290), .A2(new_n291), .A3(G264), .A4(G1698), .ZN(new_n292));
  INV_X1    g0092(.A(G1698), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n290), .A2(new_n291), .A3(G257), .A4(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n289), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n210), .B1(G33), .B2(G41), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n284), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n270), .A2(new_n298), .A3(G169), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT21), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n298), .A2(G200), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n257), .A2(new_n263), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n269), .A2(new_n268), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G190), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n306), .A2(KEYINPUT80), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(KEYINPUT80), .ZN(new_n308));
  OR2_X1    g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n284), .A2(new_n297), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n302), .A2(new_n305), .A3(new_n310), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n270), .A2(new_n298), .A3(KEYINPUT21), .A4(G169), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n270), .A2(G179), .A3(new_n297), .A4(new_n284), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n301), .A2(new_n311), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT83), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n312), .A2(new_n313), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT83), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n316), .A2(new_n317), .A3(new_n301), .A4(new_n311), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g0119(.A(KEYINPUT3), .B(G33), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n320), .A2(G232), .A3(new_n293), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n320), .A2(G238), .A3(G1698), .ZN(new_n322));
  INV_X1    g0122(.A(G107), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n321), .B(new_n322), .C1(new_n323), .C2(new_n320), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n296), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n214), .B1(G41), .B2(G45), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n326), .A2(new_n282), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n275), .A2(G1), .A3(G13), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n328), .A2(new_n326), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n327), .B1(new_n329), .B2(new_n221), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G169), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  XOR2_X1   g0134(.A(KEYINPUT15), .B(G87), .Z(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT70), .ZN(new_n336));
  XNOR2_X1  g0136(.A(KEYINPUT15), .B(G87), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT70), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n211), .A2(G33), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  XOR2_X1   g0142(.A(KEYINPUT8), .B(G58), .Z(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(G20), .A2(G33), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G77), .ZN(new_n347));
  OAI22_X1  g0147(.A1(new_n344), .A2(new_n346), .B1(new_n211), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n260), .B1(new_n342), .B2(new_n348), .ZN(new_n349));
  OR3_X1    g0149(.A1(new_n258), .A2(KEYINPUT71), .A3(G77), .ZN(new_n350));
  OAI21_X1  g0150(.A(KEYINPUT71), .B1(new_n258), .B2(G77), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n260), .B1(new_n253), .B2(new_n254), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n347), .B1(new_n214), .B2(G20), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n350), .A2(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n349), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G179), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n331), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n334), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n296), .B1(new_n320), .B2(G77), .ZN(new_n360));
  XNOR2_X1  g0160(.A(KEYINPUT67), .B(G223), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(G1698), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(G222), .B2(G1698), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n360), .B1(new_n363), .B2(new_n320), .ZN(new_n364));
  AOI211_X1 g0164(.A(new_n327), .B(new_n364), .C1(G226), .C2(new_n329), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n365), .A2(G169), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n344), .A2(new_n341), .ZN(new_n367));
  OAI21_X1  g0167(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n368));
  INV_X1    g0168(.A(G150), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n368), .B1(new_n369), .B2(new_n346), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n260), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n214), .A2(G20), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n352), .A2(G50), .A3(new_n372), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n371), .B(new_n373), .C1(G50), .C2(new_n258), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n365), .A2(new_n356), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n366), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT69), .ZN(new_n377));
  OR2_X1    g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n376), .A2(new_n377), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n359), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(G200), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n331), .A2(new_n381), .ZN(new_n382));
  OR3_X1    g0182(.A1(new_n382), .A2(KEYINPUT72), .A3(new_n355), .ZN(new_n383));
  OAI21_X1  g0183(.A(KEYINPUT72), .B1(new_n382), .B2(new_n355), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n383), .B(new_n384), .C1(new_n306), .C2(new_n332), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n365), .A2(new_n381), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n386), .B1(G190), .B2(new_n365), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n374), .B(KEYINPUT9), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT10), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT10), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n387), .A2(new_n391), .A3(new_n388), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n380), .A2(new_n385), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n253), .A2(new_n202), .A3(new_n254), .ZN(new_n395));
  XNOR2_X1  g0195(.A(new_n395), .B(KEYINPUT12), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n352), .A2(G68), .A3(new_n372), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT11), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n211), .A2(G33), .A3(G77), .ZN(new_n399));
  OAI221_X1 g0199(.A(new_n399), .B1(new_n211), .B2(G68), .C1(new_n346), .C2(new_n244), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n398), .B1(new_n400), .B2(new_n260), .ZN(new_n401));
  AND3_X1   g0201(.A1(new_n400), .A2(new_n398), .A3(new_n260), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n396), .B(new_n397), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n290), .A2(new_n291), .A3(G232), .A4(G1698), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n290), .A2(new_n291), .A3(G226), .A4(new_n293), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G97), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n296), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n327), .B1(new_n329), .B2(G238), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT13), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT13), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n408), .A2(new_n412), .A3(new_n409), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(G169), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n415), .A2(KEYINPUT14), .ZN(new_n416));
  AND3_X1   g0216(.A1(new_n408), .A2(new_n412), .A3(new_n409), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n412), .B1(new_n408), .B2(new_n409), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(G179), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n415), .B2(KEYINPUT14), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n403), .B1(new_n416), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT74), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n403), .B1(new_n419), .B2(G190), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT73), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(new_n414), .B2(G200), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n425), .B(G200), .C1(new_n417), .C2(new_n418), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n423), .B(new_n424), .C1(new_n426), .C2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(G200), .B1(new_n417), .B2(new_n418), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT73), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n427), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n423), .B1(new_n433), .B2(new_n424), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n422), .B1(new_n430), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n328), .A2(G232), .A3(new_n326), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n436), .B(KEYINPUT78), .ZN(new_n437));
  INV_X1    g0237(.A(new_n327), .ZN(new_n438));
  INV_X1    g0238(.A(G87), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n287), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(G223), .A2(G1698), .ZN(new_n441));
  INV_X1    g0241(.A(G226), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n441), .B1(new_n442), .B2(G1698), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n440), .B1(new_n443), .B2(new_n320), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n438), .B1(new_n444), .B2(new_n328), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT79), .B1(new_n437), .B2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT78), .ZN(new_n447));
  XNOR2_X1  g0247(.A(new_n436), .B(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n442), .A2(G1698), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(G223), .B2(G1698), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n290), .A2(new_n291), .ZN(new_n451));
  OAI22_X1  g0251(.A1(new_n450), .A2(new_n451), .B1(new_n287), .B2(new_n439), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n327), .B1(new_n452), .B2(new_n296), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT79), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n448), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(G169), .B1(new_n446), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n448), .A2(new_n453), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(G179), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G58), .A2(G68), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n211), .B1(new_n203), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n461), .B1(G159), .B2(new_n345), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT7), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT76), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT76), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT7), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n451), .A2(new_n467), .A3(new_n211), .ZN(new_n468));
  OAI21_X1  g0268(.A(KEYINPUT75), .B1(new_n286), .B2(new_n288), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT75), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n290), .A2(new_n291), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n469), .A2(new_n211), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n468), .B1(new_n472), .B2(new_n463), .ZN(new_n473));
  OAI211_X1 g0273(.A(KEYINPUT16), .B(new_n462), .C1(new_n473), .C2(new_n202), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n467), .B1(new_n320), .B2(G20), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n451), .A2(new_n463), .A3(new_n211), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n475), .A2(new_n476), .A3(G68), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n462), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT16), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n474), .A2(new_n480), .A3(new_n260), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n343), .A2(new_n372), .ZN(new_n482));
  XOR2_X1   g0282(.A(new_n482), .B(KEYINPUT77), .Z(new_n483));
  AOI22_X1  g0283(.A1(new_n483), .A2(new_n352), .B1(new_n255), .B2(new_n344), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n459), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT18), .ZN(new_n487));
  INV_X1    g0287(.A(new_n485), .ZN(new_n488));
  AOI21_X1  g0288(.A(G200), .B1(new_n446), .B2(new_n455), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n457), .A2(new_n309), .ZN(new_n490));
  OR2_X1    g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n488), .A2(new_n491), .A3(KEYINPUT17), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n481), .B(new_n484), .C1(new_n489), .C2(new_n490), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT17), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT18), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n459), .A2(new_n485), .A3(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n487), .A2(new_n492), .A3(new_n495), .A4(new_n497), .ZN(new_n498));
  NOR3_X1   g0298(.A1(new_n394), .A2(new_n435), .A3(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n290), .A2(new_n291), .A3(new_n211), .A4(G87), .ZN(new_n500));
  NAND2_X1  g0300(.A1(KEYINPUT84), .A2(KEYINPUT22), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  XNOR2_X1  g0302(.A(new_n500), .B(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT87), .ZN(new_n504));
  OAI21_X1  g0304(.A(KEYINPUT23), .B1(new_n211), .B2(G107), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT23), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n506), .A2(new_n323), .A3(G20), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n211), .A2(G33), .A3(G116), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n505), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT86), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n505), .A2(new_n507), .A3(new_n508), .A4(KEYINPUT86), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  XOR2_X1   g0313(.A(KEYINPUT85), .B(KEYINPUT24), .Z(new_n514));
  NAND4_X1  g0314(.A1(new_n503), .A2(new_n504), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  AND2_X1   g0315(.A1(new_n515), .A2(new_n260), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n511), .A2(new_n512), .ZN(new_n517));
  XNOR2_X1  g0317(.A(new_n500), .B(new_n501), .ZN(new_n518));
  OAI21_X1  g0318(.A(KEYINPUT87), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n514), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n503), .A2(new_n504), .A3(new_n513), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n516), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n255), .A2(new_n323), .ZN(new_n524));
  XNOR2_X1  g0324(.A(new_n524), .B(KEYINPUT25), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n352), .A2(new_n262), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n525), .B1(G107), .B2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n290), .A2(new_n291), .A3(G257), .A4(G1698), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n290), .A2(new_n291), .A3(G250), .A4(new_n293), .ZN(new_n529));
  NAND2_X1  g0329(.A1(G33), .A2(G294), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n531), .A2(new_n296), .B1(new_n276), .B2(G264), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n283), .A2(new_n273), .A3(new_n271), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n381), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n532), .A2(new_n533), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n534), .B1(new_n536), .B2(G190), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n523), .A2(new_n527), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n535), .A2(new_n333), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(G179), .B2(new_n535), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n540), .B1(new_n523), .B2(new_n527), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n290), .A2(new_n291), .A3(G244), .A4(new_n293), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT4), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n320), .A2(KEYINPUT4), .A3(G244), .A4(new_n293), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n320), .A2(G250), .A3(G1698), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n545), .A2(new_n546), .A3(new_n265), .A4(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n296), .ZN(new_n549));
  INV_X1    g0349(.A(new_n280), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n273), .B1(new_n550), .B2(new_n278), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n328), .ZN(new_n552));
  INV_X1    g0352(.A(G257), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n533), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n549), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n333), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n475), .A2(new_n476), .A3(G107), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT6), .ZN(new_n560));
  NOR3_X1   g0360(.A1(new_n560), .A2(new_n266), .A3(G107), .ZN(new_n561));
  XNOR2_X1  g0361(.A(G97), .B(G107), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n561), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  OAI22_X1  g0363(.A1(new_n563), .A2(new_n211), .B1(new_n347), .B2(new_n346), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n260), .B1(new_n559), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n352), .A2(G97), .A3(new_n262), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n255), .A2(new_n266), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n554), .B1(new_n548), .B2(new_n296), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n356), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n557), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n277), .A2(G250), .ZN(new_n574));
  OAI22_X1  g0374(.A1(new_n296), .A2(new_n574), .B1(new_n282), .B2(new_n277), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n290), .A2(new_n291), .A3(G238), .A4(new_n293), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n290), .A2(new_n291), .A3(G244), .A4(G1698), .ZN(new_n577));
  NAND2_X1  g0377(.A1(G33), .A2(G116), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n575), .B1(new_n579), .B2(new_n296), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n356), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT81), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n579), .A2(new_n296), .ZN(new_n583));
  INV_X1    g0383(.A(new_n575), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n581), .A2(new_n582), .B1(new_n585), .B2(new_n333), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n580), .A2(KEYINPUT81), .A3(new_n356), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n340), .A2(new_n255), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT19), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n211), .B1(new_n406), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(G87), .B2(new_n206), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n290), .A2(new_n291), .A3(new_n211), .A4(G68), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n589), .B1(new_n341), .B2(new_n266), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n260), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n352), .A2(new_n336), .A3(new_n262), .A4(new_n339), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n588), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT82), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n588), .A2(new_n595), .A3(KEYINPUT82), .A4(new_n596), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n586), .A2(new_n587), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n571), .A2(G190), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n345), .A2(G77), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n558), .B(new_n603), .C1(new_n211), .C2(new_n563), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n568), .B1(new_n604), .B2(new_n260), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n602), .B(new_n605), .C1(new_n381), .C2(new_n571), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n352), .A2(G87), .A3(new_n262), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n588), .A2(new_n595), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n585), .A2(G200), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n608), .B(new_n609), .C1(new_n306), .C2(new_n585), .ZN(new_n610));
  AND4_X1   g0410(.A1(new_n573), .A2(new_n601), .A3(new_n606), .A4(new_n610), .ZN(new_n611));
  AND4_X1   g0411(.A1(new_n319), .A2(new_n499), .A3(new_n542), .A4(new_n611), .ZN(G372));
  OAI211_X1 g0412(.A(new_n597), .B(new_n581), .C1(G169), .C2(new_n580), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n523), .A2(new_n527), .A3(new_n537), .ZN(new_n615));
  AND4_X1   g0415(.A1(new_n615), .A2(new_n573), .A3(new_n606), .A4(new_n610), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n316), .A2(new_n301), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n523), .A2(new_n527), .ZN(new_n619));
  INV_X1    g0419(.A(new_n540), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n614), .B1(new_n616), .B2(new_n622), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n601), .A2(new_n610), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n557), .A2(new_n570), .A3(new_n572), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n624), .A2(KEYINPUT88), .A3(KEYINPUT26), .A4(new_n625), .ZN(new_n626));
  AND4_X1   g0426(.A1(KEYINPUT26), .A2(new_n625), .A3(new_n610), .A4(new_n601), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT88), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n333), .A2(new_n556), .B1(new_n565), .B2(new_n569), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n629), .A2(new_n610), .A3(new_n572), .A4(new_n613), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT26), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n628), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n626), .B1(new_n627), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n623), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n499), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n424), .B1(new_n426), .B2(new_n428), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT74), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n429), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n359), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n422), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n492), .A2(new_n495), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n487), .A2(new_n497), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n644), .A2(new_n393), .B1(new_n379), .B2(new_n378), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n635), .A2(new_n645), .ZN(G369));
  NAND3_X1  g0446(.A1(new_n214), .A2(new_n211), .A3(G13), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(G213), .A3(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(G343), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n270), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n654), .B1(new_n315), .B2(new_n318), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT89), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n617), .A2(new_n654), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n658), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT89), .B1(new_n655), .B2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n659), .A2(G330), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n619), .A2(new_n652), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n621), .A2(new_n663), .A3(new_n615), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n541), .A2(new_n652), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n652), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n542), .A2(new_n617), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n541), .A2(new_n667), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n666), .A2(new_n670), .ZN(G399));
  INV_X1    g0471(.A(G41), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n229), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT90), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n675), .A2(new_n214), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n208), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n678), .B1(new_n679), .B2(new_n675), .ZN(new_n680));
  XOR2_X1   g0480(.A(new_n680), .B(KEYINPUT28), .Z(new_n681));
  AOI211_X1 g0481(.A(KEYINPUT29), .B(new_n652), .C1(new_n623), .C2(new_n633), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT29), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n616), .A2(new_n622), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n630), .A2(KEYINPUT26), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n625), .A2(new_n631), .A3(new_n601), .A4(new_n610), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n684), .A2(new_n613), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n683), .B1(new_n688), .B2(new_n667), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n682), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n542), .A2(new_n319), .A3(new_n611), .A4(new_n667), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n532), .A2(new_n580), .ZN(new_n692));
  AND3_X1   g0492(.A1(new_n284), .A2(new_n297), .A3(G179), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(new_n693), .A3(new_n571), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT30), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n692), .A2(new_n693), .A3(KEYINPUT30), .A4(new_n571), .ZN(new_n697));
  AOI21_X1  g0497(.A(G179), .B1(new_n284), .B2(new_n297), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n556), .A2(new_n535), .A3(new_n698), .A4(new_n585), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n696), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n700), .A2(KEYINPUT31), .A3(new_n652), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT91), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  AOI22_X1  g0503(.A1(new_n549), .A2(new_n555), .B1(new_n532), .B2(new_n533), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n704), .A2(KEYINPUT91), .A3(new_n585), .A4(new_n698), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n703), .A2(new_n696), .A3(new_n705), .A4(new_n697), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n652), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT31), .ZN(new_n708));
  AOI21_X1  g0508(.A(KEYINPUT92), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT92), .ZN(new_n710));
  AOI211_X1 g0510(.A(new_n710), .B(KEYINPUT31), .C1(new_n706), .C2(new_n652), .ZN(new_n711));
  OAI211_X1 g0511(.A(new_n691), .B(new_n701), .C1(new_n709), .C2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G330), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT93), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n712), .A2(KEYINPUT93), .A3(G330), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n690), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n681), .B1(new_n718), .B2(G1), .ZN(G364));
  AND2_X1   g0519(.A1(new_n211), .A2(G13), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n214), .B1(new_n720), .B2(G45), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n675), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n210), .B1(G20), .B2(new_n333), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n211), .A2(G179), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n727), .A2(G190), .A3(G200), .ZN(new_n728));
  INV_X1    g0528(.A(G303), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n309), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n211), .A2(new_n356), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n731), .A2(G200), .A3(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(G322), .ZN(new_n736));
  INV_X1    g0536(.A(G294), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n306), .A2(G179), .A3(G200), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(new_n211), .ZN(new_n739));
  OAI22_X1  g0539(.A1(new_n735), .A2(new_n736), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n733), .A2(new_n381), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(new_n731), .ZN(new_n743));
  XNOR2_X1  g0543(.A(KEYINPUT98), .B(G326), .ZN(new_n744));
  AOI211_X1 g0544(.A(new_n730), .B(new_n740), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G190), .A2(G200), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n732), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(G311), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n451), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n727), .A2(new_n746), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n749), .B1(G329), .B2(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n727), .A2(new_n306), .A3(G200), .ZN(new_n753));
  XOR2_X1   g0553(.A(new_n753), .B(KEYINPUT96), .Z(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G283), .ZN(new_n755));
  OAI21_X1  g0555(.A(KEYINPUT97), .B1(new_n742), .B2(G190), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n742), .A2(KEYINPUT97), .A3(G190), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  XNOR2_X1  g0560(.A(KEYINPUT33), .B(G317), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n745), .A2(new_n752), .A3(new_n755), .A4(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n728), .A2(new_n439), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n451), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT95), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(new_n760), .B2(G68), .ZN(new_n768));
  INV_X1    g0568(.A(G159), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n750), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT32), .ZN(new_n771));
  INV_X1    g0571(.A(new_n743), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n735), .A2(new_n201), .B1(new_n772), .B2(new_n244), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n739), .A2(new_n266), .B1(new_n747), .B2(new_n347), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n754), .A2(G107), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n776), .B1(new_n766), .B2(new_n765), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n768), .A2(new_n771), .A3(new_n775), .A4(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n726), .B1(new_n763), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G13), .A2(G33), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(G20), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n725), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n229), .A2(G355), .A3(new_n320), .ZN(new_n784));
  INV_X1    g0584(.A(new_n229), .ZN(new_n785));
  AND3_X1   g0585(.A1(new_n290), .A2(new_n291), .A3(new_n470), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n470), .B1(new_n290), .B2(new_n291), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(new_n272), .B2(new_n249), .ZN(new_n791));
  AND2_X1   g0591(.A1(new_n209), .A2(new_n272), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n784), .B1(G116), .B2(new_n229), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n724), .B(new_n779), .C1(new_n783), .C2(new_n793), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n659), .A2(new_n661), .ZN(new_n795));
  INV_X1    g0595(.A(new_n782), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n795), .A2(G330), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n662), .B(new_n724), .C1(new_n798), .C2(KEYINPUT94), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n798), .A2(KEYINPUT94), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n797), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT99), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(G396));
  INV_X1    g0603(.A(new_n716), .ZN(new_n804));
  AOI21_X1  g0604(.A(KEYINPUT93), .B1(new_n712), .B2(G330), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n634), .A2(new_n667), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n358), .A2(new_n652), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n355), .A2(new_n652), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n385), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n808), .B1(new_n810), .B2(new_n358), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n807), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n634), .A2(new_n811), .A3(new_n667), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n723), .B1(new_n806), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n806), .B2(new_n815), .ZN(new_n817));
  INV_X1    g0617(.A(new_n747), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n734), .A2(G143), .B1(G159), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(G137), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n819), .B1(new_n820), .B2(new_n772), .C1(new_n759), .C2(new_n369), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT34), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n754), .A2(G68), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n788), .B1(G132), .B2(new_n751), .ZN(new_n824));
  INV_X1    g0624(.A(new_n739), .ZN(new_n825));
  INV_X1    g0625(.A(new_n728), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n825), .A2(G58), .B1(new_n826), .B2(G50), .ZN(new_n827));
  AND4_X1   g0627(.A1(new_n822), .A2(new_n823), .A3(new_n824), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n754), .A2(G87), .ZN(new_n829));
  XNOR2_X1  g0629(.A(KEYINPUT100), .B(G283), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n829), .B1(new_n759), .B2(new_n830), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n825), .A2(G97), .B1(new_n826), .B2(G107), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n832), .B1(new_n772), .B2(new_n729), .C1(new_n737), .C2(new_n735), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n451), .B1(new_n750), .B2(new_n748), .C1(new_n256), .C2(new_n747), .ZN(new_n834));
  NOR3_X1   g0634(.A1(new_n831), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n725), .B1(new_n828), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n726), .A2(new_n781), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n723), .B1(G77), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n836), .B(new_n839), .C1(new_n811), .C2(new_n781), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n817), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(G384));
  NAND2_X1  g0642(.A1(new_n562), .A2(new_n560), .ZN(new_n843));
  INV_X1    g0643(.A(new_n561), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OR2_X1    g0645(.A1(new_n845), .A2(KEYINPUT35), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(KEYINPUT35), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n846), .A2(G116), .A3(new_n212), .A4(new_n847), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n848), .B(KEYINPUT36), .Z(new_n849));
  NAND3_X1  g0649(.A1(new_n679), .A2(G77), .A3(new_n460), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n214), .B(G13), .C1(new_n850), .C2(new_n245), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT40), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT7), .B1(new_n788), .B2(new_n211), .ZN(new_n854));
  OAI21_X1  g0654(.A(G68), .B1(new_n854), .B2(new_n468), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT16), .B1(new_n855), .B2(new_n462), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n474), .A2(new_n260), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n484), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n650), .B1(new_n456), .B2(new_n458), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n488), .A2(new_n491), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT37), .ZN(new_n861));
  OAI21_X1  g0661(.A(KEYINPUT101), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n650), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n485), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n486), .A2(new_n864), .A3(new_n861), .A4(new_n493), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT101), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n858), .A2(new_n859), .ZN(new_n867));
  INV_X1    g0667(.A(new_n493), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n866), .B(KEYINPUT37), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n862), .A2(new_n865), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n498), .A2(new_n863), .A3(new_n858), .ZN(new_n871));
  AND3_X1   g0671(.A1(new_n870), .A2(KEYINPUT38), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT38), .B1(new_n870), .B2(new_n871), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n403), .A2(new_n652), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n435), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n638), .A2(new_n422), .A3(new_n875), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n707), .A2(new_n708), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n706), .A2(KEYINPUT31), .A3(new_n652), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n691), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n879), .A2(new_n811), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n853), .B1(new_n874), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT38), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n864), .B1(new_n643), .B2(new_n641), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n486), .A2(new_n864), .A3(new_n493), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n887), .B(new_n861), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n885), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n870), .A2(KEYINPUT38), .A3(new_n871), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n879), .A2(new_n811), .A3(new_n882), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n891), .A2(new_n892), .A3(KEYINPUT40), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n884), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n894), .A2(new_n499), .A3(new_n882), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(G330), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n894), .B1(new_n499), .B2(new_n882), .ZN(new_n897));
  OR2_X1    g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT39), .B1(new_n872), .B2(new_n873), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT39), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n889), .A2(new_n890), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n899), .A2(KEYINPUT102), .A3(new_n901), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n422), .A2(new_n652), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT102), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n905), .B(KEYINPUT39), .C1(new_n872), .C2(new_n873), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n902), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n643), .A2(new_n863), .ZN(new_n908));
  INV_X1    g0708(.A(new_n879), .ZN(new_n909));
  INV_X1    g0709(.A(new_n808), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n909), .B1(new_n814), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n870), .A2(new_n871), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n885), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n890), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n908), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n907), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n499), .B1(new_n689), .B2(new_n682), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n645), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n916), .B(new_n918), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n898), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT103), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI221_X1 g0722(.A(new_n922), .B1(new_n214), .B2(new_n720), .C1(new_n919), .C2(new_n898), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n920), .A2(new_n921), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n852), .B1(new_n923), .B2(new_n924), .ZN(G367));
  OAI211_X1 g0725(.A(new_n606), .B(new_n573), .C1(new_n605), .C2(new_n667), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n625), .A2(new_n652), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n668), .A2(new_n928), .ZN(new_n929));
  OR3_X1    g0729(.A1(new_n929), .A2(KEYINPUT104), .A3(KEYINPUT42), .ZN(new_n930));
  OAI21_X1  g0730(.A(KEYINPUT104), .B1(new_n929), .B2(KEYINPUT42), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n929), .A2(KEYINPUT42), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n573), .B1(new_n621), .B2(new_n926), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n667), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n930), .A2(new_n931), .A3(new_n932), .A4(new_n934), .ZN(new_n935));
  OR3_X1    g0735(.A1(new_n613), .A2(new_n608), .A3(new_n667), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n610), .B(new_n613), .C1(new_n608), .C2(new_n667), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(KEYINPUT43), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n935), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n938), .A2(KEYINPUT43), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n940), .A2(new_n941), .ZN(new_n944));
  INV_X1    g0744(.A(new_n666), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n943), .A2(new_n944), .B1(new_n945), .B2(new_n928), .ZN(new_n946));
  INV_X1    g0746(.A(new_n944), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n945), .A2(new_n928), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n947), .A2(new_n948), .A3(new_n942), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n675), .B(new_n952), .Z(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT108), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n617), .A2(new_n667), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n664), .A2(new_n665), .A3(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT107), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n664), .A2(KEYINPUT107), .A3(new_n665), .A4(new_n956), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n959), .A2(new_n668), .A3(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(new_n662), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n955), .B1(new_n717), .B2(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n795), .A2(new_n961), .A3(G330), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n662), .A2(new_n668), .A3(new_n959), .A4(new_n960), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n806), .A2(new_n966), .A3(KEYINPUT108), .A4(new_n690), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n963), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT109), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n963), .A2(new_n967), .A3(KEYINPUT109), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n670), .A2(new_n928), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT45), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n670), .A2(new_n928), .ZN(new_n974));
  XOR2_X1   g0774(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n975));
  XNOR2_X1  g0775(.A(new_n974), .B(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(new_n945), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n970), .A2(new_n971), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n954), .B1(new_n979), .B2(new_n718), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n951), .B1(new_n980), .B2(new_n722), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n320), .B1(new_n750), .B2(new_n820), .C1(new_n244), .C2(new_n747), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n201), .A2(new_n728), .B1(new_n753), .B2(new_n347), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n982), .B(new_n983), .C1(new_n760), .C2(G159), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n743), .A2(G143), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n985), .B1(new_n202), .B2(new_n739), .C1(new_n735), .C2(new_n369), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n986), .A2(KEYINPUT110), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(KEYINPUT110), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n984), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(KEYINPUT46), .B1(new_n728), .B2(new_n256), .ZN(new_n990));
  OR3_X1    g0790(.A1(new_n728), .A2(KEYINPUT46), .A3(new_n256), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n760), .A2(G294), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(G317), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n747), .A2(new_n830), .B1(new_n750), .B2(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n789), .A2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n753), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n825), .A2(G107), .B1(new_n996), .B2(G97), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n734), .A2(G303), .B1(new_n743), .B2(G311), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n992), .A2(new_n995), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n989), .A2(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(KEYINPUT111), .B(KEYINPUT47), .Z(new_n1001));
  XNOR2_X1  g0801(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n725), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n936), .A2(new_n937), .A3(new_n782), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n790), .A2(new_n239), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n783), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n340), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1006), .B1(new_n785), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n724), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1003), .A2(new_n1004), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n981), .A2(new_n1010), .ZN(G387));
  OAI21_X1  g0811(.A(new_n790), .B1(new_n236), .B2(new_n272), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n229), .A2(new_n677), .A3(new_n320), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OR3_X1    g0814(.A1(new_n344), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1015));
  OAI21_X1  g0815(.A(KEYINPUT50), .B1(new_n344), .B2(G50), .ZN(new_n1016));
  AOI21_X1  g0816(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1015), .A2(new_n676), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n1014), .A2(new_n1018), .B1(new_n323), .B2(new_n785), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n723), .B1(new_n1019), .B2(new_n1006), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n760), .A2(new_n343), .B1(G97), .B2(new_n754), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n735), .A2(new_n244), .B1(new_n772), .B2(new_n769), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(G77), .B2(new_n826), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1007), .A2(new_n825), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n747), .A2(new_n202), .B1(new_n750), .B2(new_n369), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n788), .A2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1021), .A2(new_n1023), .A3(new_n1024), .A4(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n789), .B1(new_n751), .B2(new_n744), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n739), .A2(new_n830), .B1(new_n728), .B2(new_n737), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT112), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n743), .A2(G322), .B1(G303), .B2(new_n818), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n993), .B2(new_n735), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(G311), .B2(new_n760), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1030), .B1(new_n1033), .B2(KEYINPUT48), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(KEYINPUT48), .B2(new_n1033), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT49), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1028), .B1(new_n256), .B2(new_n753), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  AND2_X1   g0837(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1027), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1020), .B1(new_n1039), .B2(new_n725), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n664), .A2(new_n665), .A3(new_n782), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n966), .A2(new_n722), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n968), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n675), .B(KEYINPUT113), .Z(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n718), .B2(new_n966), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1042), .B1(new_n1043), .B2(new_n1045), .ZN(G393));
  INV_X1    g0846(.A(new_n1044), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n977), .B(new_n666), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1047), .B1(new_n1048), .B2(new_n968), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n979), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n978), .A2(new_n722), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n343), .A2(new_n818), .B1(new_n751), .B2(G143), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n739), .A2(new_n347), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(G68), .B2(new_n826), .ZN(new_n1054));
  AND4_X1   g0854(.A1(new_n789), .A2(new_n829), .A3(new_n1052), .A4(new_n1054), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n734), .A2(G159), .B1(new_n743), .B2(G150), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT115), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n1058), .A2(KEYINPUT51), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1058), .A2(KEYINPUT51), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1055), .B1(new_n244), .B2(new_n759), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(KEYINPUT116), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n734), .A2(G311), .B1(new_n743), .B2(G317), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT52), .Z(new_n1064));
  OAI221_X1 g0864(.A(new_n451), .B1(new_n750), .B2(new_n736), .C1(new_n737), .C2(new_n747), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n739), .A2(new_n256), .B1(new_n728), .B2(new_n830), .ZN(new_n1066));
  NOR3_X1   g0866(.A1(new_n776), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1064), .B(new_n1067), .C1(new_n729), .C2(new_n759), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1062), .A2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1061), .A2(KEYINPUT116), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n725), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n928), .A2(new_n782), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT114), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n790), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n783), .B1(new_n266), .B2(new_n229), .C1(new_n1074), .C2(new_n243), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1071), .A2(new_n723), .A3(new_n1073), .A4(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1050), .A2(new_n1051), .A3(new_n1076), .ZN(G390));
  OAI21_X1  g0877(.A(new_n723), .B1(new_n343), .B2(new_n837), .ZN(new_n1078));
  INV_X1    g0878(.A(G283), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n735), .A2(new_n256), .B1(new_n772), .B2(new_n1079), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n451), .B1(new_n750), .B2(new_n737), .C1(new_n266), .C2(new_n747), .ZN(new_n1081));
  OR4_X1    g0881(.A1(new_n764), .A2(new_n1080), .A3(new_n1053), .A4(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n823), .B1(new_n759), .B2(new_n323), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n760), .A2(G137), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(KEYINPUT54), .B(G143), .ZN(new_n1085));
  INV_X1    g0885(.A(G125), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n747), .A2(new_n1085), .B1(new_n750), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(G159), .B2(new_n825), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n734), .A2(G132), .B1(new_n743), .B2(G128), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n728), .A2(new_n369), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT53), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1084), .A2(new_n1088), .A3(new_n1089), .A4(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n320), .B1(new_n753), .B2(new_n244), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n1093), .B(KEYINPUT118), .Z(new_n1094));
  OAI22_X1  g0894(.A1(new_n1082), .A2(new_n1083), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1078), .B1(new_n1095), .B2(new_n725), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n906), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n905), .B1(new_n914), .B2(KEYINPUT39), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1097), .B1(new_n1098), .B2(new_n901), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1096), .B1(new_n1099), .B2(new_n781), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n652), .B1(new_n623), .B2(new_n687), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n810), .A2(new_n358), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n808), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  OR2_X1    g0903(.A1(new_n1103), .A2(new_n909), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1104), .A2(new_n903), .A3(new_n891), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n812), .B1(new_n715), .B2(new_n716), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n879), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n911), .A2(new_n904), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1105), .B(new_n1107), .C1(new_n1099), .C2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n892), .A2(G330), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1108), .B1(new_n902), .B2(new_n906), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1105), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1109), .A2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1100), .B1(new_n1115), .B2(new_n721), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n882), .A2(G330), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n499), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n917), .A2(new_n1119), .A3(new_n645), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1110), .B1(new_n1106), .B2(new_n879), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n814), .A2(new_n910), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1118), .A2(KEYINPUT117), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT117), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n811), .B1(new_n1117), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n909), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1107), .A2(new_n1103), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1120), .B1(new_n1123), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1129), .A2(new_n1109), .A3(new_n1114), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1123), .A2(new_n1128), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1120), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1047), .B1(new_n1115), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1116), .B1(new_n1130), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(G378));
  NAND2_X1  g0936(.A1(new_n760), .A2(G132), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1085), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n826), .A2(new_n1138), .B1(new_n818), .B2(G137), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n734), .A2(G128), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n743), .A2(G125), .B1(G150), .B2(new_n825), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1137), .A2(new_n1139), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  OR2_X1    g0942(.A1(new_n1142), .A2(KEYINPUT59), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(KEYINPUT59), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n996), .A2(G159), .ZN(new_n1145));
  AOI211_X1 g0945(.A(G33), .B(G41), .C1(new_n751), .C2(G124), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1143), .A2(new_n1144), .A3(new_n1145), .A4(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n734), .A2(G107), .ZN(new_n1148));
  XOR2_X1   g0948(.A(new_n1148), .B(KEYINPUT120), .Z(new_n1149));
  NAND2_X1  g0949(.A1(new_n760), .A2(G97), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n743), .A2(G116), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n753), .A2(new_n201), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(G77), .B2(new_n826), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .A4(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n340), .A2(new_n747), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n788), .A2(new_n672), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n739), .A2(new_n202), .B1(new_n1079), .B2(new_n750), .ZN(new_n1157));
  NOR4_X1   g0957(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  OR2_X1    g0958(.A1(new_n1158), .A2(KEYINPUT58), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(KEYINPUT58), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1156), .B(new_n244), .C1(G33), .C2(G41), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT119), .ZN(new_n1162));
  AND4_X1   g0962(.A1(new_n1147), .A2(new_n1159), .A3(new_n1160), .A4(new_n1162), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n723), .B1(G50), .B2(new_n837), .C1(new_n1163), .C2(new_n726), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n374), .A2(new_n863), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n393), .A2(new_n376), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1167), .B1(new_n393), .B2(new_n376), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1166), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1170), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1172), .A2(new_n1168), .A3(new_n1165), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1164), .B1(new_n1175), .B2(new_n780), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n883), .B1(new_n913), .B2(new_n890), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n893), .B(G330), .C1(new_n1177), .C2(KEYINPUT40), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(new_n1175), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n884), .A2(new_n1174), .A3(G330), .A4(new_n893), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n916), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1179), .A2(new_n907), .A3(new_n1180), .A4(new_n915), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1176), .B1(new_n1184), .B2(new_n722), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n916), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT121), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1186), .A2(new_n1187), .A3(new_n1180), .A4(new_n1179), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1183), .A2(KEYINPUT121), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1188), .A2(new_n1189), .A3(new_n1182), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1190), .A2(new_n1191), .A3(KEYINPUT57), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(new_n1044), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1130), .A2(new_n1132), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1194), .A2(KEYINPUT57), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1185), .B1(new_n1193), .B2(new_n1195), .ZN(G375));
  NAND3_X1  g0996(.A1(new_n1123), .A2(new_n1128), .A3(new_n1120), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1133), .A2(new_n953), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n909), .A2(new_n780), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n723), .B1(G68), .B2(new_n837), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n760), .A2(G116), .B1(G77), .B2(new_n754), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n451), .B1(new_n750), .B2(new_n729), .C1(new_n323), .C2(new_n747), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n1007), .B2(new_n825), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n826), .A2(G97), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n734), .A2(G283), .B1(new_n743), .B2(G294), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1201), .A2(new_n1203), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  XOR2_X1   g1006(.A(new_n1206), .B(KEYINPUT122), .Z(new_n1207));
  OAI22_X1  g1007(.A1(new_n739), .A2(new_n244), .B1(new_n747), .B2(new_n369), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT123), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n735), .A2(new_n820), .B1(new_n769), .B2(new_n728), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1152), .B(new_n1210), .C1(G132), .C2(new_n743), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n788), .B1(G128), .B2(new_n751), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1211), .B(new_n1212), .C1(new_n759), .C2(new_n1085), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1207), .B1(new_n1209), .B2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1200), .B1(new_n1214), .B2(new_n725), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1131), .A2(new_n722), .B1(new_n1199), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1198), .A2(new_n1216), .ZN(G381));
  OAI211_X1 g1017(.A(new_n1192), .B(new_n1044), .C1(KEYINPUT57), .C2(new_n1194), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1218), .A2(new_n1135), .A3(new_n1185), .ZN(new_n1219));
  OR4_X1    g1019(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1220));
  OR4_X1    g1020(.A1(G387), .A2(new_n1219), .A3(new_n1220), .A4(G381), .ZN(G407));
  OAI211_X1 g1021(.A(G407), .B(G213), .C1(G343), .C2(new_n1219), .ZN(G409));
  INV_X1    g1022(.A(KEYINPUT60), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1197), .A2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1224), .A2(new_n1044), .A3(new_n1133), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT124), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n1197), .B2(new_n1223), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1197), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1228), .A2(KEYINPUT124), .A3(KEYINPUT60), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1225), .B1(new_n1227), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1216), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n841), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1225), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1229), .A2(new_n1227), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1235), .A2(G384), .A3(new_n1216), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n651), .A2(G213), .A3(G2897), .ZN(new_n1237));
  AND3_X1   g1037(.A1(new_n1232), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1237), .B1(new_n1232), .B2(new_n1236), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(G375), .A2(G378), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1194), .A2(new_n953), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1176), .B1(new_n1190), .B2(new_n722), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1135), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n651), .A2(G213), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1241), .A2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(KEYINPUT61), .B1(new_n1240), .B2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT63), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1232), .A2(new_n1236), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1250), .B1(new_n1248), .B2(new_n1251), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n981), .A2(new_n1010), .A3(G390), .ZN(new_n1253));
  AOI21_X1  g1053(.A(G390), .B1(new_n981), .B2(new_n1010), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(G393), .B(new_n802), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(new_n1253), .A2(new_n1254), .A3(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(G390), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n963), .A2(new_n967), .A3(KEYINPUT109), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT109), .B1(new_n963), .B2(new_n967), .ZN(new_n1260));
  NOR3_X1   g1060(.A1(new_n1259), .A2(new_n1260), .A3(new_n1048), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n953), .B1(new_n1261), .B2(new_n717), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n950), .B1(new_n1262), .B2(new_n721), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1010), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1258), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n981), .A2(new_n1010), .A3(G390), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1255), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1257), .A2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1135), .B1(new_n1218), .B2(new_n1185), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1269), .A2(new_n1246), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1251), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1270), .A2(KEYINPUT63), .A3(new_n1271), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1249), .A2(new_n1252), .A3(new_n1268), .A4(new_n1272), .ZN(new_n1273));
  OAI211_X1 g1073(.A(KEYINPUT125), .B(KEYINPUT62), .C1(new_n1248), .C2(new_n1251), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n1275));
  OR2_X1    g1075(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1270), .A2(new_n1275), .A3(new_n1276), .A4(new_n1271), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1274), .A2(new_n1249), .A3(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT126), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1279), .B1(new_n1257), .B2(new_n1267), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1256), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1265), .A2(new_n1255), .A3(new_n1266), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1281), .A2(new_n1282), .A3(KEYINPUT126), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1280), .A2(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1273), .B1(new_n1278), .B2(new_n1284), .ZN(G405));
  INV_X1    g1085(.A(KEYINPUT127), .ZN(new_n1286));
  AND3_X1   g1086(.A1(new_n1218), .A2(new_n1135), .A3(new_n1185), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1286), .B1(new_n1287), .B2(new_n1269), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1241), .A2(KEYINPUT127), .A3(new_n1219), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1288), .A2(new_n1251), .A3(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1251), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(new_n1290), .A2(new_n1291), .A3(new_n1284), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1281), .A2(KEYINPUT126), .A3(new_n1282), .ZN(new_n1293));
  AOI21_X1  g1093(.A(KEYINPUT126), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  NOR3_X1   g1095(.A1(new_n1287), .A2(new_n1269), .A3(new_n1286), .ZN(new_n1296));
  AOI21_X1  g1096(.A(KEYINPUT127), .B1(new_n1241), .B2(new_n1219), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1271), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1288), .A2(new_n1251), .A3(new_n1289), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1295), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1292), .A2(new_n1300), .ZN(G402));
endmodule


