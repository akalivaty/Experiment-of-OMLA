//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 0 0 1 0 0 1 0 0 0 1 1 1 1 0 1 0 0 0 1 0 0 1 1 0 1 0 0 0 1 1 1 0 0 0 1 0 1 1 0 0 1 0 1 0 0 1 1 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n842,
    new_n843, new_n844, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n202));
  INV_X1    g001(.A(G120gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G113gat), .ZN(new_n204));
  INV_X1    g003(.A(G113gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G120gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT1), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G134gat), .ZN(new_n210));
  AND2_X1   g009(.A1(new_n210), .A2(KEYINPUT67), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(KEYINPUT67), .ZN(new_n212));
  OAI21_X1  g011(.A(G127gat), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(G127gat), .A2(G134gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n209), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n207), .A2(KEYINPUT68), .ZN(new_n217));
  NAND2_X1  g016(.A1(G127gat), .A2(G134gat), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT1), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT68), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n206), .A3(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n217), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n216), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT25), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n225));
  INV_X1    g024(.A(G169gat), .ZN(new_n226));
  INV_X1    g025(.A(G176gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n226), .A2(new_n227), .A3(KEYINPUT64), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT64), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n229), .B1(G169gat), .B2(G176gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n230), .A3(KEYINPUT23), .ZN(new_n231));
  NAND2_X1  g030(.A1(G169gat), .A2(G176gat), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n225), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT23), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n234), .B1(G169gat), .B2(G176gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT24), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n236), .A2(G183gat), .A3(G190gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(G183gat), .B(G190gat), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n235), .B(new_n237), .C1(new_n238), .C2(new_n236), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n233), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n231), .A2(new_n225), .A3(new_n232), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n224), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(G183gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(KEYINPUT27), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT27), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(G183gat), .ZN(new_n246));
  INV_X1    g045(.A(G190gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n244), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT28), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n249), .A2(KEYINPUT66), .ZN(new_n250));
  AOI22_X1  g049(.A1(new_n248), .A2(new_n250), .B1(G183gat), .B2(G190gat), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT26), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n228), .A2(new_n230), .A3(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n254), .A2(new_n232), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT27), .B(G183gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n257), .A2(new_n258), .A3(new_n247), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n251), .A2(new_n256), .A3(new_n259), .ZN(new_n260));
  OR2_X1    g059(.A1(new_n238), .A2(new_n236), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n226), .A2(new_n227), .A3(KEYINPUT23), .ZN(new_n262));
  AND3_X1   g061(.A1(new_n235), .A2(new_n224), .A3(new_n232), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n261), .A2(new_n237), .A3(new_n262), .A4(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n260), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n223), .B1(new_n242), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n231), .A2(new_n232), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT65), .ZN(new_n268));
  INV_X1    g067(.A(new_n239), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n268), .A2(new_n269), .A3(new_n241), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT25), .ZN(new_n271));
  AND2_X1   g070(.A1(new_n260), .A2(new_n264), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n216), .A2(new_n222), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G227gat), .ZN(new_n275));
  INV_X1    g074(.A(G233gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n266), .A2(new_n274), .A3(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT33), .ZN(new_n279));
  XNOR2_X1  g078(.A(G15gat), .B(G43gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(KEYINPUT69), .ZN(new_n281));
  XNOR2_X1  g080(.A(G71gat), .B(G99gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n278), .B(KEYINPUT32), .C1(new_n279), .C2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n284), .B1(new_n278), .B2(KEYINPUT32), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n278), .A2(new_n279), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT70), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n287), .A2(KEYINPUT70), .A3(new_n288), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n286), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n266), .A2(new_n274), .ZN(new_n294));
  INV_X1    g093(.A(new_n277), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n296), .A2(KEYINPUT34), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n296), .A2(KEYINPUT34), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n202), .B1(new_n293), .B2(new_n299), .ZN(new_n300));
  AND3_X1   g099(.A1(new_n287), .A2(KEYINPUT70), .A3(new_n288), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT70), .B1(new_n287), .B2(new_n288), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n285), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n299), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n299), .B(new_n285), .C1(new_n301), .C2(new_n302), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n300), .B1(new_n307), .B2(new_n202), .ZN(new_n308));
  XOR2_X1   g107(.A(G78gat), .B(G106gat), .Z(new_n309));
  XNOR2_X1  g108(.A(new_n309), .B(KEYINPUT81), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT31), .B(G50gat), .ZN(new_n311));
  XOR2_X1   g110(.A(new_n310), .B(new_n311), .Z(new_n312));
  INV_X1    g111(.A(G228gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n313), .A2(new_n276), .ZN(new_n314));
  NAND2_X1  g113(.A1(G155gat), .A2(G162gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(G155gat), .A2(G162gat), .ZN(new_n317));
  OAI21_X1  g116(.A(KEYINPUT77), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(G155gat), .ZN(new_n319));
  INV_X1    g118(.A(G162gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT77), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n321), .A2(new_n322), .A3(new_n315), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n315), .A2(KEYINPUT2), .ZN(new_n325));
  INV_X1    g124(.A(G148gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n326), .A2(G141gat), .ZN(new_n327));
  INV_X1    g126(.A(G141gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n328), .A2(G148gat), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n325), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT78), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n331), .B1(new_n326), .B2(G141gat), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n328), .A2(KEYINPUT78), .A3(G148gat), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n332), .B(new_n333), .C1(new_n328), .C2(G148gat), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n315), .B1(new_n321), .B2(KEYINPUT2), .ZN(new_n335));
  AOI22_X1  g134(.A1(new_n324), .A2(new_n330), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  XOR2_X1   g135(.A(G211gat), .B(G218gat), .Z(new_n337));
  INV_X1    g136(.A(KEYINPUT22), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n338), .A2(KEYINPUT73), .B1(G211gat), .B2(G218gat), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT74), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT73), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT22), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n339), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(G197gat), .B(G204gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n340), .B1(new_n339), .B2(new_n342), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n337), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n346), .ZN(new_n348));
  INV_X1    g147(.A(new_n337), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n348), .A2(new_n349), .A3(new_n343), .A4(new_n344), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT29), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT3), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n336), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT79), .B1(new_n336), .B2(new_n354), .ZN(new_n356));
  NOR3_X1   g155(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT77), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n322), .B1(new_n321), .B2(new_n315), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n330), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n334), .A2(new_n335), .ZN(new_n360));
  AND4_X1   g159(.A1(KEYINPUT79), .A2(new_n359), .A3(new_n354), .A4(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n352), .B1(new_n356), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n351), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT82), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n355), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n362), .A2(KEYINPUT82), .A3(new_n363), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n314), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT3), .B1(new_n351), .B2(new_n352), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n314), .B1(new_n369), .B2(new_n336), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT83), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n351), .B1(new_n362), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT79), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n359), .A2(new_n360), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n373), .B1(new_n374), .B2(KEYINPUT3), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n336), .A2(KEYINPUT79), .A3(new_n354), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT29), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT83), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n370), .B1(new_n372), .B2(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n368), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(KEYINPUT85), .A2(G22gat), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n312), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI211_X1 g181(.A(KEYINPUT85), .B(G22gat), .C1(new_n368), .C2(new_n379), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT84), .ZN(new_n385));
  OAI21_X1  g184(.A(G22gat), .B1(new_n368), .B2(new_n379), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n365), .B1(new_n377), .B2(new_n351), .ZN(new_n387));
  INV_X1    g186(.A(new_n355), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(new_n388), .A3(new_n367), .ZN(new_n389));
  INV_X1    g188(.A(new_n314), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n379), .ZN(new_n392));
  INV_X1    g191(.A(G22gat), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n386), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n385), .B1(new_n395), .B2(new_n312), .ZN(new_n396));
  INV_X1    g195(.A(new_n312), .ZN(new_n397));
  AOI211_X1 g196(.A(KEYINPUT84), .B(new_n397), .C1(new_n386), .C2(new_n394), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n384), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n336), .A2(new_n216), .A3(new_n222), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT4), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n223), .A2(KEYINPUT4), .A3(new_n336), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(G225gat), .A2(G233gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n374), .A2(KEYINPUT3), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n273), .B(new_n406), .C1(new_n356), .C2(new_n361), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n404), .A2(KEYINPUT5), .A3(new_n405), .A4(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n273), .B1(new_n336), .B2(new_n354), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n409), .B1(new_n375), .B2(new_n376), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n402), .A2(new_n403), .ZN(new_n411));
  INV_X1    g210(.A(new_n405), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT5), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n273), .A2(new_n374), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n414), .B1(new_n416), .B2(new_n412), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n408), .B1(new_n413), .B2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(G1gat), .B(G29gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(KEYINPUT0), .ZN(new_n420));
  XNOR2_X1  g219(.A(G57gat), .B(G85gat), .ZN(new_n421));
  XOR2_X1   g220(.A(new_n420), .B(new_n421), .Z(new_n422));
  NAND2_X1  g221(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT6), .ZN(new_n424));
  INV_X1    g223(.A(new_n422), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n425), .B(new_n408), .C1(new_n413), .C2(new_n417), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n423), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n426), .A2(new_n424), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT75), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n352), .B1(new_n242), .B2(new_n265), .ZN(new_n432));
  NAND2_X1  g231(.A1(G226gat), .A2(G233gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  OAI211_X1 g233(.A(G226gat), .B(G233gat), .C1(new_n242), .C2(new_n265), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(new_n351), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n351), .B1(new_n434), .B2(new_n435), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n431), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(G8gat), .B(G36gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(G64gat), .B(G92gat), .ZN(new_n441));
  XOR2_X1   g240(.A(new_n440), .B(new_n441), .Z(new_n442));
  XNOR2_X1  g241(.A(new_n442), .B(KEYINPUT76), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n434), .A2(new_n435), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n363), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n445), .A2(KEYINPUT75), .A3(new_n436), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n439), .A2(new_n443), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n445), .A2(new_n442), .A3(new_n436), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT30), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n445), .A2(KEYINPUT30), .A3(new_n442), .A4(new_n436), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n447), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NOR3_X1   g251(.A1(new_n430), .A2(new_n452), .A3(KEYINPUT35), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n308), .A2(new_n399), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n307), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n428), .B1(new_n427), .B2(KEYINPUT80), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT80), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n423), .A2(new_n457), .A3(new_n424), .A4(new_n426), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n452), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n399), .A2(new_n455), .A3(new_n459), .ZN(new_n460));
  AOI22_X1  g259(.A1(KEYINPUT88), .A2(new_n454), .B1(new_n460), .B2(KEYINPUT35), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT88), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n308), .A2(new_n399), .A3(new_n462), .A4(new_n453), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n305), .A2(KEYINPUT36), .A3(new_n306), .ZN(new_n464));
  OR2_X1    g263(.A1(new_n464), .A2(KEYINPUT71), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(KEYINPUT71), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n465), .B(new_n466), .C1(new_n308), .C2(KEYINPUT36), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n459), .B(new_n384), .C1(new_n396), .C2(new_n398), .ZN(new_n468));
  XOR2_X1   g267(.A(KEYINPUT87), .B(KEYINPUT39), .Z(new_n469));
  INV_X1    g268(.A(KEYINPUT86), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n404), .A2(new_n407), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n470), .B1(new_n471), .B2(new_n412), .ZN(new_n472));
  AOI211_X1 g271(.A(KEYINPUT86), .B(new_n405), .C1(new_n404), .C2(new_n407), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n469), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n471), .A2(new_n470), .A3(new_n412), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n412), .B1(new_n410), .B2(new_n411), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT86), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n415), .A2(new_n400), .A3(new_n405), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n475), .A2(new_n477), .A3(KEYINPUT39), .A4(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n474), .A2(new_n422), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT40), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n474), .A2(new_n479), .A3(KEYINPUT40), .A4(new_n422), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n482), .A2(new_n426), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n439), .A2(KEYINPUT37), .A3(new_n446), .ZN(new_n485));
  INV_X1    g284(.A(new_n442), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT37), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n445), .A2(new_n487), .A3(new_n436), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n485), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT38), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT37), .B1(new_n437), .B2(new_n438), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT38), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n443), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n491), .A2(new_n488), .A3(new_n493), .ZN(new_n494));
  AND4_X1   g293(.A1(new_n427), .A2(new_n429), .A3(new_n494), .A4(new_n448), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n484), .A2(new_n452), .B1(new_n490), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n399), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n468), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n461), .A2(new_n463), .B1(new_n467), .B2(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(G113gat), .B(G141gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(G197gat), .ZN(new_n501));
  XOR2_X1   g300(.A(KEYINPUT11), .B(G169gat), .Z(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(KEYINPUT89), .B(KEYINPUT12), .ZN(new_n504));
  XOR2_X1   g303(.A(new_n503), .B(new_n504), .Z(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(G29gat), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n507), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n508));
  AND2_X1   g307(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n509));
  NOR2_X1   g308(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n508), .B1(new_n511), .B2(G36gat), .ZN(new_n512));
  OR2_X1    g311(.A1(new_n512), .A2(KEYINPUT15), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(KEYINPUT15), .ZN(new_n514));
  XNOR2_X1  g313(.A(G43gat), .B(G50gat), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  OR2_X1    g315(.A1(new_n514), .A2(new_n515), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G15gat), .B(G22gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT90), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(G1gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT16), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n519), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n519), .A2(new_n520), .A3(G1gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT91), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n528), .B1(new_n519), .B2(G1gat), .ZN(new_n529));
  INV_X1    g328(.A(G8gat), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OR2_X1    g330(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n527), .A2(new_n531), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n518), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n532), .A2(new_n533), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT92), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n518), .B(KEYINPUT17), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n535), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G229gat), .A2(G233gat), .ZN(new_n541));
  NOR2_X1   g340(.A1(KEYINPUT93), .A2(KEYINPUT18), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n540), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n518), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n536), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n546), .A2(KEYINPUT94), .A3(new_n534), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT94), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n545), .A2(new_n536), .A3(new_n548), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n541), .B(KEYINPUT13), .Z(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n544), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n543), .B1(new_n540), .B2(new_n541), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n506), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n539), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(new_n534), .ZN(new_n557));
  INV_X1    g356(.A(new_n541), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n542), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n559), .A2(new_n505), .A3(new_n552), .A4(new_n544), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G85gat), .A2(G92gat), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT101), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(KEYINPUT101), .A2(G85gat), .A3(G92gat), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n565), .A2(KEYINPUT7), .A3(new_n566), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n567), .A2(KEYINPUT102), .ZN(new_n568));
  XOR2_X1   g367(.A(KEYINPUT103), .B(G92gat), .Z(new_n569));
  INV_X1    g368(.A(G85gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(G99gat), .A2(G106gat), .ZN(new_n571));
  AOI22_X1  g370(.A1(new_n569), .A2(new_n570), .B1(KEYINPUT8), .B2(new_n571), .ZN(new_n572));
  OR2_X1    g371(.A1(new_n563), .A2(KEYINPUT7), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n567), .A2(KEYINPUT102), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n568), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G99gat), .B(G106gat), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n575), .A2(KEYINPUT104), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n575), .A2(new_n577), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT104), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n568), .A2(new_n572), .A3(new_n576), .A4(new_n574), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n539), .A2(new_n578), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n578), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(new_n518), .ZN(new_n585));
  XNOR2_X1  g384(.A(G190gat), .B(G218gat), .ZN(new_n586));
  AND2_X1   g385(.A1(G232gat), .A2(G233gat), .ZN(new_n587));
  AOI22_X1  g386(.A1(new_n586), .A2(KEYINPUT105), .B1(KEYINPUT41), .B2(new_n587), .ZN(new_n588));
  AND2_X1   g387(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n583), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n586), .A2(KEYINPUT105), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n590), .B(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n587), .A2(KEYINPUT41), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT100), .ZN(new_n595));
  XNOR2_X1  g394(.A(G134gat), .B(G162gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n593), .B(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(G71gat), .B(G78gat), .Z(new_n600));
  NOR2_X1   g399(.A1(new_n600), .A2(KEYINPUT95), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT9), .ZN(new_n602));
  INV_X1    g401(.A(G71gat), .ZN(new_n603));
  INV_X1    g402(.A(G78gat), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(G57gat), .B(G64gat), .Z(new_n606));
  AOI21_X1  g405(.A(new_n601), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n600), .A2(KEYINPUT95), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n600), .A2(new_n606), .A3(KEYINPUT95), .A4(new_n605), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT21), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(new_n536), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT99), .ZN(new_n614));
  XNOR2_X1  g413(.A(G127gat), .B(G155gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT20), .ZN(new_n616));
  NAND2_X1  g415(.A1(G231gat), .A2(G233gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT97), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n616), .B(new_n618), .Z(new_n619));
  XNOR2_X1  g418(.A(new_n614), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(KEYINPUT96), .B(KEYINPUT21), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n609), .A2(new_n621), .A3(new_n610), .ZN(new_n622));
  XOR2_X1   g421(.A(KEYINPUT98), .B(KEYINPUT19), .Z(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G183gat), .B(G211gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n620), .B(new_n626), .Z(new_n627));
  NAND2_X1  g426(.A1(G230gat), .A2(G233gat), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT10), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n611), .A2(new_n579), .A3(new_n581), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n630), .B(new_n631), .C1(new_n584), .C2(new_n611), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n584), .A2(KEYINPUT10), .A3(new_n611), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n629), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n631), .B1(new_n584), .B2(new_n611), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n635), .A2(new_n629), .ZN(new_n636));
  XNOR2_X1  g435(.A(G120gat), .B(G148gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(G176gat), .B(G204gat), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n637), .B(new_n638), .Z(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  OR3_X1    g439(.A1(new_n634), .A2(new_n636), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT106), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n640), .B1(new_n634), .B2(new_n636), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  OAI211_X1 g443(.A(KEYINPUT106), .B(new_n640), .C1(new_n634), .C2(new_n636), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n599), .A2(new_n627), .A3(new_n646), .ZN(new_n647));
  NOR3_X1   g446(.A1(new_n499), .A2(new_n562), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n456), .A2(new_n458), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(G1gat), .ZN(G1324gat));
  INV_X1    g451(.A(new_n648), .ZN(new_n653));
  INV_X1    g452(.A(new_n452), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g454(.A(KEYINPUT16), .B(G8gat), .Z(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n657), .B1(new_n530), .B2(new_n655), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(KEYINPUT42), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT42), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(G1325gat));
  OR2_X1    g461(.A1(new_n467), .A2(KEYINPUT107), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n467), .A2(KEYINPUT107), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(G15gat), .B1(new_n653), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(G15gat), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n648), .A2(new_n667), .A3(new_n308), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n666), .A2(new_n668), .ZN(G1326gat));
  NAND2_X1  g468(.A1(new_n648), .A2(new_n497), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT108), .ZN(new_n671));
  XOR2_X1   g470(.A(KEYINPUT43), .B(G22gat), .Z(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(G1327gat));
  INV_X1    g472(.A(new_n627), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n674), .A2(new_n561), .A3(new_n646), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n499), .A2(KEYINPUT110), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n454), .A2(KEYINPUT88), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n460), .A2(KEYINPUT35), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n677), .A2(new_n678), .A3(new_n463), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n498), .A2(new_n467), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT110), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n676), .A2(new_n683), .A3(new_n684), .A4(new_n598), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n599), .B1(new_n679), .B2(new_n680), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n686), .A2(new_n684), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n675), .B1(new_n685), .B2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(G29gat), .B1(new_n690), .B2(new_n649), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n674), .A2(new_n598), .A3(new_n646), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n499), .A2(new_n562), .A3(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT109), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n649), .A2(G29gat), .ZN(new_n695));
  AND3_X1   g494(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n694), .B1(new_n693), .B2(new_n695), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT45), .ZN(new_n698));
  OR3_X1    g497(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n698), .B1(new_n696), .B2(new_n697), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n691), .A2(new_n699), .A3(new_n700), .ZN(G1328gat));
  OAI21_X1  g500(.A(G36gat), .B1(new_n690), .B2(new_n654), .ZN(new_n702));
  AOI21_X1  g501(.A(G36gat), .B1(KEYINPUT111), .B2(KEYINPUT46), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n693), .A2(new_n452), .A3(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n702), .A2(new_n706), .ZN(G1329gat));
  INV_X1    g506(.A(G43gat), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n693), .A2(new_n708), .A3(new_n308), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(KEYINPUT112), .ZN(new_n710));
  INV_X1    g509(.A(new_n665), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n689), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n710), .B1(new_n712), .B2(G43gat), .ZN(new_n713));
  NAND2_X1  g512(.A1(KEYINPUT47), .A2(G43gat), .ZN(new_n714));
  INV_X1    g513(.A(new_n467), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n714), .B1(new_n689), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n709), .B1(KEYINPUT112), .B2(KEYINPUT47), .ZN(new_n717));
  OAI22_X1  g516(.A1(new_n713), .A2(KEYINPUT47), .B1(new_n716), .B2(new_n717), .ZN(G1330gat));
  AOI21_X1  g517(.A(G50gat), .B1(new_n693), .B2(new_n497), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n497), .A2(G50gat), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n719), .B1(new_n689), .B2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT48), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(G1331gat));
  AND3_X1   g522(.A1(new_n679), .A2(KEYINPUT110), .A3(new_n680), .ZN(new_n724));
  AOI21_X1  g523(.A(KEYINPUT110), .B1(new_n679), .B2(new_n680), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR4_X1   g525(.A1(new_n674), .A2(new_n598), .A3(new_n561), .A4(new_n646), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n650), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(G57gat), .ZN(G1332gat));
  NAND3_X1  g529(.A1(new_n726), .A2(new_n452), .A3(new_n727), .ZN(new_n731));
  XOR2_X1   g530(.A(KEYINPUT49), .B(G64gat), .Z(new_n732));
  OR2_X1    g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n731), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT113), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT113), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n733), .A2(new_n737), .A3(new_n734), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(G1333gat));
  NAND3_X1  g538(.A1(new_n728), .A2(new_n603), .A3(new_n308), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n726), .A2(new_n727), .ZN(new_n741));
  OAI21_X1  g540(.A(G71gat), .B1(new_n741), .B2(new_n665), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT50), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(G1334gat));
  NOR2_X1   g544(.A1(new_n741), .A2(new_n399), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(new_n604), .ZN(G1335gat));
  NAND2_X1  g546(.A1(new_n685), .A2(new_n688), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n627), .A2(new_n561), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n750), .A2(new_n646), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(KEYINPUT114), .B1(new_n752), .B2(new_n649), .ZN(new_n753));
  INV_X1    g552(.A(new_n751), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n754), .B1(new_n685), .B2(new_n688), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT114), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n755), .A2(new_n756), .A3(new_n650), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n753), .A2(G85gat), .A3(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT115), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n750), .B1(new_n686), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(KEYINPUT115), .B1(new_n499), .B2(new_n599), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT51), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n760), .A2(KEYINPUT51), .A3(new_n761), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n646), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n766), .A2(new_n570), .A3(new_n650), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n758), .A2(new_n767), .ZN(G1336gat));
  INV_X1    g567(.A(new_n569), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(new_n752), .B2(new_n654), .ZN(new_n770));
  INV_X1    g569(.A(G92gat), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n646), .A2(new_n654), .ZN(new_n772));
  AND3_X1   g571(.A1(new_n760), .A2(KEYINPUT51), .A3(new_n761), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT51), .B1(new_n760), .B2(new_n761), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n771), .B(new_n772), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  XNOR2_X1  g574(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n770), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n776), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n569), .B1(new_n755), .B2(new_n452), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n772), .A2(new_n771), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n780), .B1(new_n764), .B2(new_n765), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n778), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n777), .A2(new_n782), .ZN(G1337gat));
  INV_X1    g582(.A(G99gat), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n766), .A2(new_n784), .A3(new_n308), .ZN(new_n785));
  OAI21_X1  g584(.A(G99gat), .B1(new_n752), .B2(new_n665), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(G1338gat));
  INV_X1    g586(.A(new_n646), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n399), .A2(G106gat), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n788), .B(new_n789), .C1(new_n773), .C2(new_n774), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n598), .A2(new_n684), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n724), .A2(new_n725), .A3(new_n791), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n497), .B(new_n751), .C1(new_n792), .C2(new_n687), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(G106gat), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n790), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT53), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n790), .A2(new_n797), .A3(new_n794), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(G1339gat));
  NOR2_X1   g598(.A1(new_n647), .A2(new_n561), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n634), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n632), .A2(new_n629), .A3(new_n633), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n634), .A2(new_n801), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n805), .B1(new_n806), .B2(new_n640), .ZN(new_n807));
  AOI211_X1 g606(.A(KEYINPUT117), .B(new_n639), .C1(new_n634), .C2(new_n801), .ZN(new_n808));
  OAI211_X1 g607(.A(KEYINPUT55), .B(new_n804), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n809), .A2(new_n641), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n540), .A2(new_n541), .ZN(new_n811));
  OAI22_X1  g610(.A1(new_n811), .A2(KEYINPUT118), .B1(new_n551), .B2(new_n550), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n557), .A2(KEYINPUT118), .A3(new_n558), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n503), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n814), .A2(new_n560), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n804), .B1(new_n807), .B2(new_n808), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n810), .A2(new_n815), .A3(new_n598), .A4(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n788), .A2(new_n560), .A3(new_n814), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n818), .A2(new_n561), .A3(new_n641), .A4(new_n809), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n819), .B1(new_n822), .B2(new_n598), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n800), .B1(new_n823), .B2(new_n674), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n824), .A2(new_n649), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n497), .A2(new_n307), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n825), .A2(new_n654), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n827), .A2(new_n205), .A3(new_n561), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT119), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n824), .A2(new_n497), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n649), .A2(new_n452), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n308), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n561), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n829), .B1(new_n835), .B2(G113gat), .ZN(new_n836));
  AOI211_X1 g635(.A(KEYINPUT119), .B(new_n205), .C1(new_n834), .C2(new_n561), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n828), .B1(new_n836), .B2(new_n837), .ZN(G1340gat));
  NOR3_X1   g637(.A1(new_n833), .A2(new_n203), .A3(new_n646), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n827), .A2(new_n788), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n839), .B1(new_n840), .B2(new_n203), .ZN(G1341gat));
  INV_X1    g640(.A(G127gat), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n827), .A2(new_n842), .A3(new_n627), .ZN(new_n843));
  OAI21_X1  g642(.A(G127gat), .B1(new_n833), .B2(new_n674), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(G1342gat));
  NOR3_X1   g644(.A1(new_n599), .A2(new_n211), .A3(new_n212), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n827), .A2(new_n846), .ZN(new_n847));
  OR2_X1    g646(.A1(new_n847), .A2(KEYINPUT56), .ZN(new_n848));
  OAI21_X1  g647(.A(G134gat), .B1(new_n833), .B2(new_n599), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(KEYINPUT56), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(G1343gat));
  AOI21_X1  g650(.A(new_n399), .B1(new_n663), .B2(new_n664), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n825), .A2(new_n654), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n853), .A2(new_n328), .A3(new_n561), .ZN(new_n854));
  AND3_X1   g653(.A1(new_n561), .A2(new_n641), .A3(new_n809), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n816), .A2(KEYINPUT120), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT120), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n857), .B(new_n804), .C1(new_n807), .C2(new_n808), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n856), .A2(new_n817), .A3(new_n858), .ZN(new_n859));
  AOI22_X1  g658(.A1(new_n855), .A2(new_n859), .B1(new_n788), .B2(new_n815), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n819), .B1(new_n860), .B2(new_n598), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n800), .B1(new_n861), .B2(new_n674), .ZN(new_n862));
  OAI21_X1  g661(.A(KEYINPUT57), .B1(new_n862), .B2(new_n399), .ZN(new_n863));
  INV_X1    g662(.A(new_n819), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n598), .B1(new_n820), .B2(new_n821), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n674), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n800), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT57), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n868), .A2(new_n869), .A3(new_n497), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n467), .A2(new_n831), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n863), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(G141gat), .B1(new_n872), .B2(new_n562), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n854), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(KEYINPUT58), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT58), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n854), .A2(new_n873), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n877), .ZN(G1344gat));
  NAND3_X1  g677(.A1(new_n853), .A2(new_n326), .A3(new_n788), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT121), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n627), .B1(new_n861), .B2(new_n881), .ZN(new_n882));
  OAI211_X1 g681(.A(KEYINPUT121), .B(new_n819), .C1(new_n860), .C2(new_n598), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n800), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n399), .A2(KEYINPUT57), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT57), .B1(new_n824), .B2(new_n399), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n887), .A2(new_n788), .A3(new_n871), .A4(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n880), .B1(new_n889), .B2(G148gat), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n872), .A2(new_n646), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n891), .A2(KEYINPUT59), .A3(new_n326), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n879), .B1(new_n890), .B2(new_n892), .ZN(G1345gat));
  NAND3_X1  g692(.A1(new_n853), .A2(new_n319), .A3(new_n627), .ZN(new_n894));
  OAI21_X1  g693(.A(G155gat), .B1(new_n872), .B2(new_n674), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1346gat));
  AOI21_X1  g695(.A(G162gat), .B1(new_n853), .B2(new_n598), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n872), .A2(new_n320), .A3(new_n599), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n897), .A2(new_n898), .ZN(G1347gat));
  AOI21_X1  g698(.A(new_n650), .B1(new_n866), .B2(new_n867), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n826), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n901), .A2(new_n654), .ZN(new_n902));
  AOI21_X1  g701(.A(G169gat), .B1(new_n902), .B2(new_n561), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n650), .A2(new_n654), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n904), .A2(new_n308), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n830), .A2(new_n905), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n906), .A2(new_n226), .A3(new_n562), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n903), .A2(new_n907), .ZN(G1348gat));
  OAI21_X1  g707(.A(G176gat), .B1(new_n906), .B2(new_n646), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n772), .A2(new_n227), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n901), .B2(new_n910), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT122), .ZN(G1349gat));
  NAND4_X1  g711(.A1(new_n868), .A2(new_n399), .A3(new_n627), .A4(new_n905), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n243), .B1(new_n913), .B2(KEYINPUT123), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n914), .B1(KEYINPUT123), .B2(new_n913), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n902), .A2(new_n257), .A3(new_n627), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g717(.A1(new_n902), .A2(new_n247), .A3(new_n598), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n830), .A2(new_n598), .A3(new_n905), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n920), .A2(new_n921), .A3(G190gat), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n921), .B1(new_n920), .B2(G190gat), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n919), .B1(new_n922), .B2(new_n923), .ZN(G1351gat));
  AND2_X1   g723(.A1(new_n665), .A2(new_n904), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n888), .B(new_n925), .C1(new_n884), .C2(new_n886), .ZN(new_n926));
  INV_X1    g725(.A(G197gat), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n926), .A2(new_n927), .A3(new_n562), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n900), .A2(new_n852), .A3(new_n452), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT124), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n561), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n928), .B1(new_n931), .B2(new_n927), .ZN(G1352gat));
  XNOR2_X1  g731(.A(KEYINPUT125), .B(G204gat), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n934), .B1(new_n926), .B2(new_n646), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n900), .A2(new_n852), .A3(new_n772), .A4(new_n933), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT62), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n936), .B(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT126), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n935), .A2(KEYINPUT126), .A3(new_n938), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(G1353gat));
  INV_X1    g742(.A(G211gat), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n930), .A2(new_n944), .A3(new_n627), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n887), .A2(new_n627), .A3(new_n888), .A4(new_n925), .ZN(new_n946));
  AOI21_X1  g745(.A(KEYINPUT63), .B1(new_n946), .B2(G211gat), .ZN(new_n947));
  OAI211_X1 g746(.A(KEYINPUT63), .B(G211gat), .C1(new_n926), .C2(new_n674), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n945), .B1(new_n947), .B2(new_n949), .ZN(G1354gat));
  AOI21_X1  g749(.A(G218gat), .B1(new_n930), .B2(new_n598), .ZN(new_n951));
  INV_X1    g750(.A(new_n926), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n598), .A2(G218gat), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT127), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n951), .B1(new_n952), .B2(new_n954), .ZN(G1355gat));
endmodule


