//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 1 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 1 0 0 1 0 0 0 0 0 1 0 0 0 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n851, new_n852, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976;
  INV_X1    g000(.A(KEYINPUT99), .ZN(new_n202));
  AND2_X1   g001(.A1(G232gat), .A2(G233gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT41), .ZN(new_n204));
  AOI21_X1  g003(.A(KEYINPUT84), .B1(G29gat), .B2(G36gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  NAND3_X1  g005(.A1(KEYINPUT84), .A2(G29gat), .A3(G36gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(KEYINPUT85), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT85), .ZN(new_n209));
  INV_X1    g008(.A(new_n207), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n209), .B1(new_n210), .B2(new_n205), .ZN(new_n211));
  AND2_X1   g010(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G50gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G43gat), .ZN(new_n214));
  INV_X1    g013(.A(G43gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G50gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT15), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n214), .A2(new_n216), .A3(KEYINPUT15), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT14), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(G29gat), .B2(G36gat), .ZN(new_n222));
  INV_X1    g021(.A(G29gat), .ZN(new_n223));
  INV_X1    g022(.A(G36gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT14), .ZN(new_n225));
  AND3_X1   g024(.A1(new_n220), .A2(new_n222), .A3(new_n225), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n212), .A2(KEYINPUT86), .A3(new_n219), .A4(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT86), .ZN(new_n228));
  AND2_X1   g027(.A1(new_n225), .A2(new_n222), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n219), .A2(new_n229), .A3(new_n220), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n208), .A2(new_n211), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n228), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n229), .A2(new_n207), .A3(new_n206), .ZN(new_n233));
  INV_X1    g032(.A(new_n220), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n227), .A2(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT7), .ZN(new_n236));
  OAI211_X1 g035(.A(G85gat), .B(G92gat), .C1(new_n236), .C2(KEYINPUT96), .ZN(new_n237));
  NAND2_X1  g036(.A1(G85gat), .A2(G92gat), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT96), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n238), .A2(new_n239), .A3(KEYINPUT7), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G99gat), .B(G106gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(G99gat), .A2(G106gat), .ZN(new_n243));
  INV_X1    g042(.A(G85gat), .ZN(new_n244));
  INV_X1    g043(.A(G92gat), .ZN(new_n245));
  AOI22_X1  g044(.A1(KEYINPUT8), .A2(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  AND4_X1   g045(.A1(KEYINPUT97), .A2(new_n241), .A3(new_n242), .A4(new_n246), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n241), .A2(new_n242), .A3(new_n246), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n242), .B1(new_n241), .B2(new_n246), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT97), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n247), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n204), .B1(new_n235), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n227), .A2(new_n232), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n233), .A2(new_n234), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT87), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT17), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT17), .ZN(new_n259));
  NOR3_X1   g058(.A1(new_n235), .A2(KEYINPUT87), .A3(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n252), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT98), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n256), .A2(new_n257), .A3(KEYINPUT17), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n259), .B1(new_n235), .B2(KEYINPUT87), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n266), .A2(KEYINPUT98), .A3(new_n252), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n253), .B1(new_n263), .B2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G190gat), .B(G218gat), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n202), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n203), .A2(KEYINPUT41), .ZN(new_n272));
  XNOR2_X1  g071(.A(G134gat), .B(G162gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n268), .A2(new_n270), .ZN(new_n276));
  AOI211_X1 g075(.A(new_n269), .B(new_n253), .C1(new_n263), .C2(new_n267), .ZN(new_n277));
  OAI22_X1  g076(.A1(new_n271), .A2(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n263), .A2(new_n267), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n269), .B1(new_n279), .B2(new_n253), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n268), .A2(new_n270), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n280), .A2(new_n202), .A3(new_n281), .A4(new_n274), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G127gat), .ZN(new_n285));
  INV_X1    g084(.A(G57gat), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT93), .B1(new_n286), .B2(G64gat), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT93), .ZN(new_n288));
  INV_X1    g087(.A(G64gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n288), .A2(new_n289), .A3(G57gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n286), .A2(G64gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n287), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT94), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT94), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n287), .A2(new_n290), .A3(new_n294), .A4(new_n291), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT9), .ZN(new_n297));
  OR3_X1    g096(.A1(new_n297), .A2(G71gat), .A3(G78gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(G71gat), .A2(G78gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT95), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n289), .A2(G57gat), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n297), .B1(new_n303), .B2(new_n291), .ZN(new_n304));
  NOR3_X1   g103(.A1(KEYINPUT92), .A2(G71gat), .A3(G78gat), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT92), .B1(G71gat), .B2(G78gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(new_n299), .ZN(new_n307));
  NOR3_X1   g106(.A1(new_n304), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n301), .A2(new_n302), .A3(new_n309), .ZN(new_n310));
  AOI22_X1  g109(.A1(new_n293), .A2(new_n295), .B1(new_n299), .B2(new_n298), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT95), .B1(new_n311), .B2(new_n308), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G231gat), .ZN(new_n314));
  INV_X1    g113(.A(G233gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OR3_X1    g115(.A1(new_n313), .A2(KEYINPUT21), .A3(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n316), .B1(new_n313), .B2(KEYINPUT21), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n285), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n313), .A2(KEYINPUT21), .ZN(new_n321));
  XNOR2_X1  g120(.A(G15gat), .B(G22gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT16), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n322), .B1(new_n323), .B2(G1gat), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT88), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n324), .B(new_n325), .C1(G1gat), .C2(new_n322), .ZN(new_n326));
  XOR2_X1   g125(.A(new_n326), .B(G8gat), .Z(new_n327));
  AND2_X1   g126(.A1(new_n321), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n317), .A2(new_n285), .A3(new_n318), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n320), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n329), .B1(new_n320), .B2(new_n330), .ZN(new_n332));
  XNOR2_X1  g131(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n333));
  INV_X1    g132(.A(G155gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  XOR2_X1   g134(.A(G183gat), .B(G211gat), .Z(new_n336));
  XNOR2_X1  g135(.A(new_n335), .B(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  OR3_X1    g137(.A1(new_n331), .A2(new_n332), .A3(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n338), .B1(new_n331), .B2(new_n332), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n252), .A2(new_n310), .A3(new_n312), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT100), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n252), .A2(new_n310), .A3(new_n312), .A4(KEYINPUT100), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n301), .A2(new_n250), .A3(new_n309), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT101), .B(KEYINPUT10), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n344), .A2(new_n345), .A3(new_n346), .A4(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT10), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n252), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(new_n313), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(G230gat), .A2(G233gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n346), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n355), .B1(new_n342), .B2(new_n343), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n353), .B1(new_n356), .B2(new_n345), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G120gat), .B(G148gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(G176gat), .B(G204gat), .ZN(new_n360));
  XOR2_X1   g159(.A(new_n359), .B(new_n360), .Z(new_n361));
  NAND3_X1  g160(.A1(new_n354), .A2(new_n358), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n361), .ZN(new_n363));
  INV_X1    g162(.A(new_n353), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n364), .B1(new_n348), .B2(new_n351), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n363), .B1(new_n365), .B2(new_n357), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n284), .A2(new_n341), .A3(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G197gat), .B(G204gat), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT22), .ZN(new_n371));
  INV_X1    g170(.A(G211gat), .ZN(new_n372));
  INV_X1    g171(.A(G218gat), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT72), .ZN(new_n376));
  XNOR2_X1  g175(.A(G211gat), .B(G218gat), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n375), .A2(KEYINPUT72), .A3(new_n377), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(G226gat), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n383), .A2(new_n315), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n384), .A2(KEYINPUT29), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT73), .ZN(new_n387));
  INV_X1    g186(.A(G169gat), .ZN(new_n388));
  INV_X1    g187(.A(G176gat), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n389), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n390), .B1(KEYINPUT26), .B2(new_n391), .ZN(new_n392));
  NOR3_X1   g191(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n393));
  AND2_X1   g192(.A1(new_n393), .A2(KEYINPUT66), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n393), .A2(KEYINPUT66), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n392), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(G183gat), .A2(G190gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n399));
  XOR2_X1   g198(.A(KEYINPUT64), .B(G190gat), .Z(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT27), .B(G183gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g201(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n399), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OR2_X1    g203(.A1(new_n402), .A2(new_n399), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n398), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n390), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT23), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n391), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n388), .A2(new_n389), .A3(KEYINPUT23), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n407), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n411), .A2(KEYINPUT25), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n397), .A2(KEYINPUT24), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT24), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n414), .A2(G183gat), .A3(G190gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n416), .B1(G183gat), .B2(G190gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n412), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT25), .ZN(new_n419));
  INV_X1    g218(.A(G183gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n400), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n411), .B1(new_n421), .B2(new_n416), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n418), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n387), .B1(new_n406), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n405), .A2(new_n404), .ZN(new_n425));
  AND2_X1   g224(.A1(new_n396), .A2(new_n397), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n421), .A2(new_n416), .ZN(new_n428));
  INV_X1    g227(.A(new_n411), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI22_X1  g229(.A1(new_n430), .A2(KEYINPUT25), .B1(new_n417), .B2(new_n412), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n427), .A2(new_n431), .A3(KEYINPUT73), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n386), .B1(new_n424), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n427), .A2(new_n431), .A3(new_n384), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n382), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n424), .A2(new_n384), .A3(new_n432), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n427), .A2(new_n431), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n385), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n437), .A2(new_n381), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n436), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT74), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT74), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n436), .A2(new_n443), .A3(new_n440), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  XOR2_X1   g244(.A(G8gat), .B(G36gat), .Z(new_n446));
  XNOR2_X1  g245(.A(G64gat), .B(G92gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n446), .B(new_n447), .ZN(new_n448));
  XOR2_X1   g247(.A(new_n448), .B(KEYINPUT75), .Z(new_n449));
  NAND3_X1  g248(.A1(new_n436), .A2(new_n448), .A3(new_n440), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT76), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI22_X1  g251(.A1(new_n445), .A2(new_n449), .B1(new_n452), .B2(KEYINPUT30), .ZN(new_n453));
  XNOR2_X1  g252(.A(G78gat), .B(G106gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n454), .B(G22gat), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(G141gat), .B(G148gat), .ZN(new_n457));
  NAND2_X1  g256(.A1(G155gat), .A2(G162gat), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n458), .A2(KEYINPUT2), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(G162gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n334), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n458), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT77), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n462), .A2(KEYINPUT77), .A3(new_n458), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n460), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n464), .B(new_n463), .C1(new_n457), .C2(new_n459), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT79), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT78), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n377), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n375), .A2(new_n472), .A3(new_n377), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n377), .A2(new_n472), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n475), .A2(new_n374), .A3(new_n370), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n473), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n471), .B1(new_n477), .B2(KEYINPUT29), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT3), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR3_X1   g279(.A1(new_n477), .A2(new_n471), .A3(KEYINPUT29), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n470), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(G228gat), .A2(G233gat), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT3), .B1(new_n467), .B2(new_n468), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n381), .B1(new_n484), .B2(KEYINPUT29), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n482), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n483), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT29), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n379), .A2(new_n488), .A3(new_n380), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n469), .B1(new_n489), .B2(new_n479), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT80), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n485), .B1(new_n490), .B2(new_n491), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n487), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(KEYINPUT31), .B(G50gat), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n486), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n496), .B1(new_n486), .B2(new_n494), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n456), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n486), .A2(new_n494), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n495), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n486), .A2(new_n494), .A3(new_n496), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(new_n455), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT35), .ZN(new_n504));
  AND3_X1   g303(.A1(new_n499), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n484), .ZN(new_n506));
  INV_X1    g305(.A(G134gat), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT67), .B1(new_n507), .B2(G127gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(G113gat), .B(G120gat), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n508), .B1(new_n509), .B2(KEYINPUT1), .ZN(new_n510));
  XNOR2_X1  g309(.A(G127gat), .B(G134gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n467), .A2(KEYINPUT3), .A3(new_n468), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n506), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n511), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n510), .B(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n469), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT4), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(G225gat), .A2(G233gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n516), .A2(new_n469), .A3(KEYINPUT4), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n514), .A2(new_n519), .A3(new_n520), .A4(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT5), .ZN(new_n523));
  OR2_X1    g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n512), .B(new_n469), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT5), .B1(new_n525), .B2(new_n520), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(new_n522), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G1gat), .B(G29gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(KEYINPUT0), .ZN(new_n530));
  XNOR2_X1  g329(.A(G57gat), .B(G85gat), .ZN(new_n531));
  XOR2_X1   g330(.A(new_n530), .B(new_n531), .Z(new_n532));
  NAND2_X1  g331(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT6), .ZN(new_n534));
  INV_X1    g333(.A(new_n532), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n524), .A2(new_n527), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n533), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n524), .A2(new_n527), .A3(KEYINPUT6), .A4(new_n535), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT30), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n450), .A2(new_n451), .A3(new_n540), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n453), .A2(new_n505), .A3(new_n539), .A4(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT68), .B1(new_n406), .B2(new_n423), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT68), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n427), .A2(new_n431), .A3(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n543), .A2(new_n512), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(G227gat), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n547), .A2(new_n315), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n438), .A2(KEYINPUT68), .A3(new_n516), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n546), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT32), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT33), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(G15gat), .B(G43gat), .Z(new_n554));
  XNOR2_X1  g353(.A(G71gat), .B(G99gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n551), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n556), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n550), .B(KEYINPUT32), .C1(new_n552), .C2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n546), .A2(new_n549), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT34), .ZN(new_n562));
  INV_X1    g361(.A(new_n548), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n562), .B1(new_n561), .B2(new_n563), .ZN(new_n566));
  OAI21_X1  g365(.A(KEYINPUT71), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n566), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT71), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n568), .A2(new_n569), .A3(new_n564), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n560), .A2(new_n567), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n568), .A2(new_n564), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n572), .A2(KEYINPUT71), .A3(new_n557), .A4(new_n559), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(KEYINPUT82), .B1(new_n542), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n444), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n443), .B1(new_n436), .B2(new_n440), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n449), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n452), .A2(KEYINPUT30), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n579), .A2(new_n580), .A3(new_n541), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n537), .A2(new_n538), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT82), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n583), .A2(new_n584), .A3(new_n574), .A4(new_n505), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n499), .A2(new_n503), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(KEYINPUT69), .B1(new_n565), .B2(new_n566), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n560), .A2(new_n588), .ZN(new_n589));
  AOI22_X1  g388(.A1(new_n572), .A2(KEYINPUT69), .B1(new_n557), .B2(new_n559), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n587), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n539), .A2(new_n579), .A3(new_n580), .A4(new_n541), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT35), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n576), .A2(new_n585), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n525), .A2(new_n520), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT39), .ZN(new_n596));
  INV_X1    g395(.A(new_n520), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n514), .A2(new_n519), .A3(new_n521), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n597), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n532), .B1(new_n600), .B2(KEYINPUT39), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT40), .ZN(new_n602));
  OR3_X1    g401(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n602), .B1(new_n599), .B2(new_n601), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n604), .A2(new_n536), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n581), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT81), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n607), .B1(new_n441), .B2(KEYINPUT37), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT37), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n436), .A2(KEYINPUT81), .A3(new_n609), .A4(new_n440), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT38), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n449), .A2(new_n612), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n437), .A2(new_n439), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n609), .B1(new_n614), .B2(new_n382), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n381), .B1(new_n433), .B2(new_n435), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n613), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n611), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n582), .A2(new_n618), .A3(new_n450), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n445), .A2(KEYINPUT37), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n448), .B1(new_n608), .B2(new_n610), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n612), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n606), .B(new_n587), .C1(new_n619), .C2(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(KEYINPUT36), .B1(new_n589), .B2(new_n590), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT70), .B(KEYINPUT36), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n624), .B1(new_n574), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n592), .A2(new_n586), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n623), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n594), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G113gat), .B(G141gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(KEYINPUT83), .B(KEYINPUT11), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G169gat), .B(G197gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n634), .B(KEYINPUT12), .Z(new_n635));
  XNOR2_X1  g434(.A(new_n327), .B(new_n235), .ZN(new_n636));
  NAND2_X1  g435(.A1(G229gat), .A2(G233gat), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n637), .B(KEYINPUT89), .Z(new_n638));
  XOR2_X1   g437(.A(KEYINPUT90), .B(KEYINPUT13), .Z(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n327), .A2(new_n235), .ZN(new_n642));
  AOI211_X1 g441(.A(new_n638), .B(new_n642), .C1(new_n266), .C2(new_n327), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n641), .B1(new_n643), .B2(KEYINPUT18), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n642), .B1(new_n266), .B2(new_n327), .ZN(new_n645));
  INV_X1    g444(.A(new_n638), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT18), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n635), .B1(new_n644), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n647), .A2(new_n648), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n643), .A2(KEYINPUT18), .ZN(new_n652));
  INV_X1    g451(.A(new_n635), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n651), .A2(new_n652), .A3(new_n641), .A4(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n629), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT91), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n629), .A2(KEYINPUT91), .A3(new_n655), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n369), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(new_n582), .ZN(new_n661));
  XOR2_X1   g460(.A(KEYINPUT102), .B(G1gat), .Z(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(G1324gat));
  XOR2_X1   g462(.A(KEYINPUT16), .B(G8gat), .Z(new_n664));
  AND3_X1   g463(.A1(new_n660), .A2(new_n581), .A3(new_n664), .ZN(new_n665));
  AND3_X1   g464(.A1(new_n665), .A2(KEYINPUT103), .A3(KEYINPUT42), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT42), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n658), .A2(new_n659), .ZN(new_n668));
  INV_X1    g467(.A(new_n369), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n668), .A2(new_n581), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n667), .B1(new_n670), .B2(G8gat), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n671), .A2(new_n665), .ZN(new_n672));
  AOI21_X1  g471(.A(KEYINPUT103), .B1(new_n665), .B2(KEYINPUT42), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n666), .B1(new_n672), .B2(new_n673), .ZN(G1325gat));
  AOI21_X1  g473(.A(G15gat), .B1(new_n660), .B2(new_n574), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT104), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n675), .A2(new_n676), .ZN(new_n678));
  INV_X1    g477(.A(new_n626), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n679), .A2(G15gat), .ZN(new_n680));
  AOI22_X1  g479(.A1(new_n677), .A2(new_n678), .B1(new_n660), .B2(new_n680), .ZN(G1326gat));
  NAND2_X1  g480(.A1(new_n660), .A2(new_n586), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT43), .B(G22gat), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(G1327gat));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685));
  INV_X1    g484(.A(new_n628), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n594), .A2(KEYINPUT106), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT106), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n576), .A2(new_n585), .A3(new_n688), .A4(new_n593), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n686), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n685), .B1(new_n690), .B2(new_n284), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n629), .A2(KEYINPUT44), .A3(new_n283), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n341), .A2(new_n367), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n655), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n691), .A2(new_n582), .A3(new_n692), .A4(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n223), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n698), .B1(new_n697), .B2(new_n696), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n693), .A2(new_n283), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT105), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n668), .A2(new_n223), .A3(new_n582), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT45), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n699), .A2(new_n703), .ZN(G1328gat));
  AND2_X1   g503(.A1(new_n668), .A2(new_n701), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n705), .A2(new_n224), .A3(new_n581), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n706), .A2(KEYINPUT46), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n691), .A2(new_n692), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n708), .A2(new_n581), .A3(new_n695), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(G36gat), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n706), .A2(KEYINPUT46), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n707), .A2(new_n710), .A3(new_n711), .ZN(G1329gat));
  NAND4_X1  g511(.A1(new_n691), .A2(new_n679), .A3(new_n692), .A4(new_n695), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(G43gat), .ZN(new_n714));
  AOI21_X1  g513(.A(KEYINPUT47), .B1(new_n714), .B2(KEYINPUT109), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT108), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n575), .A2(G43gat), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n668), .A2(new_n716), .A3(new_n701), .A4(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(KEYINPUT91), .B1(new_n629), .B2(new_n655), .ZN(new_n719));
  INV_X1    g518(.A(new_n655), .ZN(new_n720));
  AOI211_X1 g519(.A(new_n657), .B(new_n720), .C1(new_n594), .C2(new_n628), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n701), .B(new_n717), .C1(new_n719), .C2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(KEYINPUT108), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n718), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n714), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n715), .A2(new_n725), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n724), .B(new_n714), .C1(KEYINPUT109), .C2(KEYINPUT47), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(G1330gat));
  NAND4_X1  g527(.A1(new_n691), .A2(new_n586), .A3(new_n692), .A4(new_n695), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(G50gat), .ZN(new_n730));
  AOI21_X1  g529(.A(KEYINPUT48), .B1(new_n730), .B2(KEYINPUT111), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n586), .A2(new_n213), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT110), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n705), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n730), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n734), .B(new_n730), .C1(KEYINPUT111), .C2(KEYINPUT48), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(G1331gat));
  NAND4_X1  g537(.A1(new_n284), .A2(new_n720), .A3(new_n341), .A4(new_n367), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n690), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n539), .B(KEYINPUT112), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(G57gat), .ZN(G1332gat));
  INV_X1    g542(.A(KEYINPUT49), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n581), .B1(new_n744), .B2(new_n289), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT113), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n740), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT114), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n744), .A2(new_n289), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1333gat));
  INV_X1    g549(.A(G71gat), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n740), .A2(new_n751), .A3(new_n574), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n690), .A2(new_n626), .A3(new_n739), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n753), .B2(new_n751), .ZN(new_n754));
  XOR2_X1   g553(.A(new_n754), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n586), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g556(.A1(new_n687), .A2(new_n689), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n284), .B1(new_n758), .B2(new_n628), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n341), .A2(new_n655), .ZN(new_n760));
  AOI21_X1  g559(.A(KEYINPUT51), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762));
  INV_X1    g561(.A(new_n760), .ZN(new_n763));
  NOR4_X1   g562(.A1(new_n690), .A2(new_n762), .A3(new_n284), .A4(new_n763), .ZN(new_n764));
  OR2_X1    g563(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n765), .A2(new_n244), .A3(new_n582), .A4(new_n367), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n763), .A2(new_n368), .ZN(new_n767));
  AND3_X1   g566(.A1(new_n691), .A2(new_n692), .A3(new_n767), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n768), .A2(new_n582), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n766), .B1(new_n244), .B2(new_n769), .ZN(G1336gat));
  INV_X1    g569(.A(new_n581), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n771), .A2(G92gat), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n367), .B(new_n772), .C1(new_n761), .C2(new_n764), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n691), .A2(new_n581), .A3(new_n692), .A4(new_n767), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(G92gat), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT52), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n773), .A2(new_n778), .A3(new_n775), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(G1337gat));
  NOR2_X1   g579(.A1(new_n575), .A2(G99gat), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n765), .A2(new_n367), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n768), .A2(new_n679), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(G99gat), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(G1338gat));
  NOR2_X1   g584(.A1(new_n587), .A2(G106gat), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n367), .B(new_n786), .C1(new_n761), .C2(new_n764), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n691), .A2(new_n586), .A3(new_n692), .A4(new_n767), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G106gat), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT53), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n768), .A2(KEYINPUT115), .A3(new_n586), .ZN(new_n792));
  INV_X1    g591(.A(G106gat), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n793), .B1(new_n788), .B2(new_n794), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n787), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n791), .B1(new_n796), .B2(new_n798), .ZN(G1339gat));
  INV_X1    g598(.A(new_n341), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n353), .B1(new_n350), .B2(new_n313), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n348), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(KEYINPUT54), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT55), .B1(new_n803), .B2(new_n365), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n352), .A2(new_n805), .A3(new_n353), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n363), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n362), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n805), .B1(new_n348), .B2(new_n801), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n354), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n361), .B1(new_n365), .B2(new_n805), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT55), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(KEYINPUT116), .B1(new_n808), .B2(new_n812), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n365), .A2(new_n357), .A3(new_n363), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n815), .B1(new_n354), .B2(new_n809), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n814), .B1(new_n816), .B2(new_n811), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n806), .B(new_n363), .C1(new_n803), .C2(new_n365), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n815), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT116), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n817), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n813), .A2(new_n821), .A3(new_n655), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n645), .A2(new_n646), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n636), .A2(new_n640), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n634), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n654), .A2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n367), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n283), .B1(new_n822), .B2(new_n828), .ZN(new_n829));
  AND4_X1   g628(.A1(new_n283), .A2(new_n827), .A3(new_n813), .A4(new_n821), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n800), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n284), .A2(new_n341), .A3(new_n720), .A4(new_n368), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n833), .A2(new_n741), .ZN(new_n834));
  INV_X1    g633(.A(new_n591), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n836), .A2(new_n771), .ZN(new_n837));
  AOI21_X1  g636(.A(G113gat), .B1(new_n837), .B2(new_n655), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT117), .B1(new_n833), .B2(new_n587), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n840));
  AOI211_X1 g639(.A(new_n840), .B(new_n586), .C1(new_n831), .C2(new_n832), .ZN(new_n841));
  OR2_X1    g640(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n575), .A2(new_n539), .A3(new_n581), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n655), .A2(G113gat), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n838), .B1(new_n845), .B2(new_n846), .ZN(G1340gat));
  AOI21_X1  g646(.A(G120gat), .B1(new_n837), .B2(new_n367), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n367), .A2(G120gat), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n848), .B1(new_n845), .B2(new_n849), .ZN(G1341gat));
  NAND3_X1  g649(.A1(new_n837), .A2(new_n285), .A3(new_n341), .ZN(new_n851));
  OAI21_X1  g650(.A(G127gat), .B1(new_n844), .B2(new_n800), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(G1342gat));
  NAND2_X1  g652(.A1(new_n283), .A2(new_n771), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT118), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n836), .A2(new_n507), .A3(new_n856), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n857), .A2(KEYINPUT56), .ZN(new_n858));
  OAI21_X1  g657(.A(G134gat), .B1(new_n844), .B2(new_n284), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(KEYINPUT56), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(G1343gat));
  NOR2_X1   g660(.A1(new_n679), .A2(new_n587), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n834), .A2(new_n862), .ZN(new_n863));
  NOR4_X1   g662(.A1(new_n863), .A2(G141gat), .A3(new_n581), .A4(new_n720), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT58), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n626), .A2(new_n582), .A3(new_n771), .ZN(new_n867));
  XOR2_X1   g666(.A(new_n867), .B(KEYINPUT119), .Z(new_n868));
  AOI21_X1  g667(.A(KEYINPUT57), .B1(new_n833), .B2(new_n586), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n586), .A2(KEYINPUT57), .ZN(new_n870));
  XNOR2_X1  g669(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n818), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n655), .A2(new_n817), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n283), .B1(new_n828), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n800), .B1(new_n830), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n870), .B1(new_n875), .B2(new_n832), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n868), .B1(new_n869), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(G141gat), .B1(new_n877), .B2(new_n720), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n865), .A2(new_n866), .A3(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n875), .A2(new_n832), .ZN(new_n882));
  INV_X1    g681(.A(new_n870), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n587), .B1(new_n831), .B2(new_n832), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n884), .B1(new_n885), .B2(KEYINPUT57), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(KEYINPUT121), .A3(new_n868), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n881), .A2(new_n655), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n864), .B1(new_n888), .B2(G141gat), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n879), .B1(new_n889), .B2(new_n866), .ZN(G1344gat));
  AND3_X1   g689(.A1(new_n886), .A2(KEYINPUT121), .A3(new_n868), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT121), .B1(new_n886), .B2(new_n868), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n891), .A2(new_n892), .A3(new_n368), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(G148gat), .ZN(new_n895));
  INV_X1    g694(.A(G148gat), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT57), .ZN(new_n897));
  AND4_X1   g696(.A1(new_n283), .A2(new_n827), .A3(new_n817), .A4(new_n819), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n800), .B1(new_n898), .B2(new_n874), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n899), .A2(new_n832), .ZN(new_n900));
  OAI211_X1 g699(.A(KEYINPUT122), .B(new_n897), .C1(new_n900), .C2(new_n587), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT122), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n587), .B1(new_n899), .B2(new_n832), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n902), .B1(new_n903), .B2(KEYINPUT57), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n833), .A2(new_n883), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n901), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n868), .A2(new_n367), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n896), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI22_X1  g707(.A1(new_n893), .A2(new_n895), .B1(new_n894), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n863), .A2(new_n581), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(new_n896), .A3(new_n367), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n911), .ZN(G1345gat));
  NAND2_X1  g711(.A1(new_n881), .A2(new_n887), .ZN(new_n913));
  OAI21_X1  g712(.A(G155gat), .B1(new_n913), .B2(new_n800), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n910), .A2(new_n334), .A3(new_n341), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1346gat));
  OAI21_X1  g715(.A(G162gat), .B1(new_n913), .B2(new_n284), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n856), .A2(new_n461), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n863), .B2(new_n918), .ZN(G1347gat));
  NOR2_X1   g718(.A1(new_n771), .A2(new_n582), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n833), .A2(new_n920), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n921), .A2(new_n835), .ZN(new_n922));
  AOI21_X1  g721(.A(G169gat), .B1(new_n922), .B2(new_n655), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n741), .A2(new_n771), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT123), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n925), .A2(new_n575), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n842), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n720), .A2(new_n388), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n923), .B1(new_n927), .B2(new_n928), .ZN(G1348gat));
  AOI21_X1  g728(.A(new_n389), .B1(new_n927), .B2(new_n367), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n922), .A2(new_n389), .A3(new_n367), .ZN(new_n931));
  OR2_X1    g730(.A1(new_n930), .A2(new_n931), .ZN(G1349gat));
  NAND3_X1  g731(.A1(new_n922), .A2(new_n401), .A3(new_n341), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n926), .B(new_n341), .C1(new_n839), .C2(new_n841), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(G183gat), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n936), .B(KEYINPUT60), .ZN(G1350gat));
  OAI211_X1 g736(.A(new_n926), .B(new_n283), .C1(new_n839), .C2(new_n841), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n938), .A2(KEYINPUT61), .A3(G190gat), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n283), .A2(new_n400), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n833), .A2(new_n835), .A3(new_n920), .A4(new_n940), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT124), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(KEYINPUT61), .B1(new_n938), .B2(G190gat), .ZN(new_n944));
  OAI21_X1  g743(.A(KEYINPUT125), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(new_n944), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT125), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n946), .A2(new_n947), .A3(new_n939), .A4(new_n942), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n945), .A2(new_n948), .ZN(G1351gat));
  NOR2_X1   g748(.A1(new_n925), .A2(new_n679), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n906), .A2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(G197gat), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n951), .A2(new_n952), .A3(new_n720), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n921), .A2(new_n862), .ZN(new_n954));
  AOI21_X1  g753(.A(G197gat), .B1(new_n954), .B2(new_n655), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n953), .A2(new_n955), .ZN(G1352gat));
  OAI21_X1  g755(.A(KEYINPUT126), .B1(new_n951), .B2(new_n368), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT126), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n906), .A2(new_n958), .A3(new_n367), .A4(new_n950), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n957), .A2(G204gat), .A3(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(G204gat), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n954), .A2(new_n961), .A3(new_n367), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT62), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n962), .B(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n960), .A2(new_n964), .ZN(G1353gat));
  NAND3_X1  g764(.A1(new_n954), .A2(new_n372), .A3(new_n341), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n906), .A2(new_n341), .A3(new_n950), .ZN(new_n967));
  AND3_X1   g766(.A1(new_n967), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n968));
  AOI21_X1  g767(.A(KEYINPUT63), .B1(new_n967), .B2(G211gat), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n966), .B1(new_n968), .B2(new_n969), .ZN(G1354gat));
  INV_X1    g769(.A(KEYINPUT127), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n906), .A2(new_n971), .A3(new_n950), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(new_n283), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n971), .B1(new_n906), .B2(new_n950), .ZN(new_n974));
  OAI21_X1  g773(.A(G218gat), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n954), .A2(new_n373), .A3(new_n283), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(G1355gat));
endmodule


