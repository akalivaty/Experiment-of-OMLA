

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749;

  NOR2_X1 U367 ( .A1(n633), .A2(n718), .ZN(n635) );
  OR2_X1 U368 ( .A1(n630), .A2(n402), .ZN(n401) );
  NOR2_X1 U369 ( .A1(n642), .A2(n718), .ZN(n643) );
  XNOR2_X2 U370 ( .A(n441), .B(G469), .ZN(n522) );
  XNOR2_X2 U371 ( .A(KEYINPUT4), .B(G101), .ZN(n448) );
  NOR2_X1 U372 ( .A1(n544), .A2(n429), .ZN(n688) );
  XNOR2_X2 U373 ( .A(n389), .B(KEYINPUT31), .ZN(n667) );
  NOR2_X2 U374 ( .A1(n692), .A2(n565), .ZN(n389) );
  NAND2_X1 U375 ( .A1(n549), .A2(n688), .ZN(n550) );
  NOR2_X1 U376 ( .A1(n627), .A2(n718), .ZN(n628) );
  XNOR2_X1 U377 ( .A(n600), .B(KEYINPUT19), .ZN(n605) );
  XNOR2_X1 U378 ( .A(n383), .B(G478), .ZN(n569) );
  NAND2_X1 U379 ( .A1(n400), .A2(n405), .ZN(n600) );
  AND2_X2 U380 ( .A1(n401), .A2(n352), .ZN(n400) );
  OR2_X1 U381 ( .A1(n648), .A2(G902), .ZN(n362) );
  XNOR2_X1 U382 ( .A(n430), .B(G131), .ZN(n493) );
  INV_X2 U383 ( .A(G953), .ZN(n742) );
  XNOR2_X2 U384 ( .A(n550), .B(KEYINPUT75), .ZN(n561) );
  AND2_X1 U385 ( .A1(n613), .A2(n372), .ZN(n371) );
  XNOR2_X1 U386 ( .A(G146), .B(G125), .ZN(n471) );
  XNOR2_X1 U387 ( .A(n431), .B(n502), .ZN(n737) );
  XNOR2_X1 U388 ( .A(n493), .B(G137), .ZN(n431) );
  AND2_X1 U389 ( .A1(n586), .A2(n587), .ZN(n681) );
  XNOR2_X1 U390 ( .A(G119), .B(G116), .ZN(n444) );
  INV_X1 U391 ( .A(G237), .ZN(n459) );
  INV_X1 U392 ( .A(KEYINPUT33), .ZN(n551) );
  OR2_X1 U393 ( .A1(n569), .A2(n567), .ZN(n382) );
  NOR2_X1 U394 ( .A1(n521), .A2(n679), .ZN(n364) );
  XNOR2_X1 U395 ( .A(n516), .B(KEYINPUT0), .ZN(n553) );
  NAND2_X1 U396 ( .A1(n605), .A2(n515), .ZN(n516) );
  XNOR2_X1 U397 ( .A(n455), .B(n454), .ZN(n648) );
  AND2_X1 U398 ( .A1(n390), .A2(n353), .ZN(n741) );
  XNOR2_X1 U399 ( .A(n393), .B(KEYINPUT45), .ZN(n719) );
  AND2_X1 U400 ( .A1(n585), .A2(n584), .ZN(n394) );
  XNOR2_X1 U401 ( .A(G119), .B(G137), .ZN(n407) );
  XOR2_X1 U402 ( .A(KEYINPUT88), .B(KEYINPUT23), .Z(n408) );
  XNOR2_X1 U403 ( .A(n737), .B(G146), .ZN(n455) );
  XOR2_X1 U404 ( .A(G107), .B(G140), .Z(n433) );
  NAND2_X1 U405 ( .A1(n397), .A2(n357), .ZN(n398) );
  NAND2_X1 U406 ( .A1(n719), .A2(n741), .ZN(n672) );
  INV_X1 U407 ( .A(KEYINPUT46), .ZN(n368) );
  INV_X1 U408 ( .A(n675), .ZN(n387) );
  INV_X1 U409 ( .A(KEYINPUT2), .ZN(n399) );
  INV_X1 U410 ( .A(KEYINPUT48), .ZN(n391) );
  INV_X1 U411 ( .A(KEYINPUT44), .ZN(n377) );
  XNOR2_X1 U412 ( .A(KEYINPUT83), .B(KEYINPUT3), .ZN(n445) );
  XNOR2_X1 U413 ( .A(G113), .B(KEYINPUT69), .ZN(n443) );
  XNOR2_X1 U414 ( .A(G143), .B(G128), .ZN(n470) );
  NOR2_X1 U415 ( .A1(G953), .A2(G237), .ZN(n486) );
  XOR2_X1 U416 ( .A(KEYINPUT11), .B(KEYINPUT100), .Z(n485) );
  NAND2_X1 U417 ( .A1(KEYINPUT79), .A2(n399), .ZN(n396) );
  NAND2_X1 U418 ( .A1(n672), .A2(n399), .ZN(n397) );
  NAND2_X1 U419 ( .A1(G234), .A2(G237), .ZN(n461) );
  NAND2_X1 U420 ( .A1(n618), .A2(n483), .ZN(n404) );
  NAND2_X1 U421 ( .A1(n481), .A2(n403), .ZN(n402) );
  INV_X1 U422 ( .A(n483), .ZN(n403) );
  BUF_X1 U423 ( .A(n522), .Z(n595) );
  XNOR2_X1 U424 ( .A(G128), .B(G110), .ZN(n412) );
  XNOR2_X1 U425 ( .A(G122), .B(G107), .ZN(n505) );
  XNOR2_X1 U426 ( .A(n381), .B(n379), .ZN(n503) );
  XNOR2_X1 U427 ( .A(KEYINPUT8), .B(KEYINPUT66), .ZN(n381) );
  NOR2_X1 U428 ( .A1(n380), .A2(G953), .ZN(n379) );
  INV_X1 U429 ( .A(G234), .ZN(n380) );
  XNOR2_X1 U430 ( .A(G116), .B(KEYINPUT9), .ZN(n499) );
  XOR2_X1 U431 ( .A(G104), .B(G122), .Z(n491) );
  XNOR2_X1 U432 ( .A(G113), .B(G143), .ZN(n490) );
  XNOR2_X1 U433 ( .A(n471), .B(n409), .ZN(n735) );
  XNOR2_X1 U434 ( .A(n591), .B(n590), .ZN(n703) );
  INV_X1 U435 ( .A(KEYINPUT112), .ZN(n589) );
  XNOR2_X1 U436 ( .A(n520), .B(n519), .ZN(n526) );
  BUF_X1 U437 ( .A(n549), .Z(n687) );
  XNOR2_X1 U438 ( .A(n364), .B(n355), .ZN(n363) );
  XNOR2_X1 U439 ( .A(n425), .B(n424), .ZN(n544) );
  NAND2_X1 U440 ( .A1(n384), .A2(n460), .ZN(n383) );
  XNOR2_X1 U441 ( .A(n498), .B(n497), .ZN(n567) );
  XNOR2_X1 U442 ( .A(n496), .B(G475), .ZN(n497) );
  BUF_X1 U443 ( .A(n553), .Z(n565) );
  XNOR2_X1 U444 ( .A(n455), .B(n440), .ZN(n639) );
  XNOR2_X1 U445 ( .A(n434), .B(KEYINPUT77), .ZN(n435) );
  AND2_X1 U446 ( .A1(n645), .A2(G469), .ZN(n386) );
  BUF_X1 U447 ( .A(n672), .Z(n673) );
  XNOR2_X1 U448 ( .A(n543), .B(n542), .ZN(n598) );
  NAND2_X1 U449 ( .A1(n361), .A2(n360), .ZN(n359) );
  INV_X1 U450 ( .A(n718), .ZN(n360) );
  XNOR2_X1 U451 ( .A(n649), .B(n356), .ZN(n361) );
  NAND2_X1 U452 ( .A1(n405), .A2(n354), .ZN(n347) );
  XNOR2_X1 U453 ( .A(n382), .B(KEYINPUT107), .ZN(n586) );
  XOR2_X1 U454 ( .A(n501), .B(KEYINPUT103), .Z(n348) );
  AND2_X1 U455 ( .A1(n586), .A2(n517), .ZN(n349) );
  OR2_X1 U456 ( .A1(n560), .A2(n375), .ZN(n350) );
  OR2_X1 U457 ( .A1(n748), .A2(KEYINPUT46), .ZN(n351) );
  AND2_X1 U458 ( .A1(n404), .A2(n588), .ZN(n352) );
  AND2_X1 U459 ( .A1(n617), .A2(n616), .ZN(n353) );
  AND2_X1 U460 ( .A1(n401), .A2(n404), .ZN(n354) );
  XNOR2_X1 U461 ( .A(KEYINPUT110), .B(KEYINPUT30), .ZN(n355) );
  XOR2_X1 U462 ( .A(n648), .B(KEYINPUT62), .Z(n356) );
  AND2_X1 U463 ( .A1(n618), .A2(n396), .ZN(n357) );
  XNOR2_X1 U464 ( .A(n358), .B(KEYINPUT106), .ZN(n576) );
  NAND2_X1 U465 ( .A1(n388), .A2(n387), .ZN(n358) );
  XNOR2_X1 U466 ( .A(n359), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X2 U467 ( .A(n362), .B(n458), .ZN(n521) );
  NAND2_X1 U468 ( .A1(n365), .A2(n363), .ZN(n540) );
  AND2_X1 U469 ( .A1(n564), .A2(n366), .ZN(n365) );
  INV_X1 U470 ( .A(n532), .ZN(n366) );
  NAND2_X1 U471 ( .A1(n369), .A2(n367), .ZN(n373) );
  NAND2_X1 U472 ( .A1(n598), .A2(n368), .ZN(n367) );
  NAND2_X1 U473 ( .A1(n370), .A2(n351), .ZN(n369) );
  INV_X1 U474 ( .A(n598), .ZN(n370) );
  NAND2_X1 U475 ( .A1(n373), .A2(n371), .ZN(n392) );
  NAND2_X1 U476 ( .A1(n748), .A2(KEYINPUT46), .ZN(n372) );
  NAND2_X1 U477 ( .A1(n526), .A2(n603), .ZN(n571) );
  NAND2_X1 U478 ( .A1(n350), .A2(n374), .ZN(n395) );
  NAND2_X1 U479 ( .A1(n376), .A2(n375), .ZN(n374) );
  INV_X1 U480 ( .A(KEYINPUT71), .ZN(n375) );
  NAND2_X1 U481 ( .A1(n378), .A2(n377), .ZN(n376) );
  INV_X1 U482 ( .A(n560), .ZN(n378) );
  INV_X1 U483 ( .A(n710), .ZN(n384) );
  AND2_X1 U484 ( .A1(n647), .A2(n645), .ZN(n713) );
  NAND2_X1 U485 ( .A1(n647), .A2(n385), .ZN(n632) );
  AND2_X1 U486 ( .A1(n645), .A2(G210), .ZN(n385) );
  NAND2_X1 U487 ( .A1(n647), .A2(n386), .ZN(n641) );
  NAND2_X1 U488 ( .A1(n713), .A2(G478), .ZN(n711) );
  NAND2_X1 U489 ( .A1(n667), .A2(n653), .ZN(n388) );
  XNOR2_X1 U490 ( .A(n392), .B(n391), .ZN(n390) );
  NAND2_X1 U491 ( .A1(n395), .A2(n394), .ZN(n393) );
  XNOR2_X1 U492 ( .A(n552), .B(n551), .ZN(n674) );
  NOR2_X2 U493 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U494 ( .A(n563), .B(n562), .ZN(n692) );
  NAND2_X2 U495 ( .A1(n621), .A2(n398), .ZN(n647) );
  NAND2_X1 U496 ( .A1(n630), .A2(n483), .ZN(n405) );
  XOR2_X1 U497 ( .A(n410), .B(n735), .Z(n406) );
  INV_X1 U498 ( .A(KEYINPUT86), .ZN(n434) );
  INV_X1 U499 ( .A(KEYINPUT89), .ZN(n411) );
  XNOR2_X1 U500 ( .A(n412), .B(n411), .ZN(n414) );
  XNOR2_X1 U501 ( .A(n436), .B(n435), .ZN(n439) );
  INV_X1 U502 ( .A(n676), .ZN(n587) );
  XNOR2_X1 U503 ( .A(n414), .B(n413), .ZN(n415) );
  BUF_X1 U504 ( .A(n674), .Z(n702) );
  XNOR2_X1 U505 ( .A(n406), .B(n415), .ZN(n416) );
  XNOR2_X1 U506 ( .A(n589), .B(KEYINPUT41), .ZN(n590) );
  XNOR2_X1 U507 ( .A(n479), .B(n478), .ZN(n729) );
  INV_X1 U508 ( .A(KEYINPUT108), .ZN(n546) );
  NAND2_X1 U509 ( .A1(n503), .A2(G221), .ZN(n417) );
  XNOR2_X1 U510 ( .A(n408), .B(n407), .ZN(n410) );
  XNOR2_X1 U511 ( .A(KEYINPUT10), .B(G140), .ZN(n409) );
  XOR2_X1 U512 ( .A(KEYINPUT87), .B(KEYINPUT24), .Z(n413) );
  XNOR2_X1 U513 ( .A(n417), .B(n416), .ZN(n714) );
  NOR2_X1 U514 ( .A1(G902), .A2(n714), .ZN(n425) );
  XOR2_X1 U515 ( .A(KEYINPUT20), .B(KEYINPUT91), .Z(n419) );
  XNOR2_X1 U516 ( .A(G902), .B(KEYINPUT15), .ZN(n481) );
  NAND2_X1 U517 ( .A1(G234), .A2(n481), .ZN(n418) );
  XNOR2_X1 U518 ( .A(n419), .B(n418), .ZN(n426) );
  NAND2_X1 U519 ( .A1(n426), .A2(G217), .ZN(n423) );
  XOR2_X1 U520 ( .A(KEYINPUT25), .B(KEYINPUT93), .Z(n421) );
  XOR2_X1 U521 ( .A(KEYINPUT90), .B(KEYINPUT92), .Z(n420) );
  XNOR2_X1 U522 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U523 ( .A(n423), .B(n422), .ZN(n424) );
  NAND2_X1 U524 ( .A1(G221), .A2(n426), .ZN(n428) );
  INV_X1 U525 ( .A(KEYINPUT21), .ZN(n427) );
  XNOR2_X1 U526 ( .A(n428), .B(n427), .ZN(n683) );
  XNOR2_X1 U527 ( .A(n683), .B(KEYINPUT94), .ZN(n517) );
  INV_X1 U528 ( .A(n517), .ZN(n429) );
  XNOR2_X2 U529 ( .A(KEYINPUT67), .B(KEYINPUT68), .ZN(n430) );
  XNOR2_X1 U530 ( .A(n470), .B(G134), .ZN(n502) );
  NAND2_X1 U531 ( .A1(G227), .A2(n742), .ZN(n432) );
  XNOR2_X1 U532 ( .A(n433), .B(n432), .ZN(n436) );
  XNOR2_X1 U533 ( .A(KEYINPUT82), .B(G110), .ZN(n437) );
  XNOR2_X1 U534 ( .A(n437), .B(G104), .ZN(n727) );
  XNOR2_X1 U535 ( .A(n448), .B(KEYINPUT70), .ZN(n438) );
  XNOR2_X1 U536 ( .A(n727), .B(n438), .ZN(n476) );
  XNOR2_X1 U537 ( .A(n439), .B(n476), .ZN(n440) );
  INV_X1 U538 ( .A(G902), .ZN(n460) );
  NAND2_X1 U539 ( .A1(n639), .A2(n460), .ZN(n441) );
  NAND2_X1 U540 ( .A1(n688), .A2(n595), .ZN(n442) );
  XNOR2_X1 U541 ( .A(n442), .B(KEYINPUT95), .ZN(n564) );
  XNOR2_X1 U542 ( .A(n444), .B(n443), .ZN(n446) );
  XNOR2_X1 U543 ( .A(n446), .B(n445), .ZN(n479) );
  XNOR2_X1 U544 ( .A(KEYINPUT76), .B(KEYINPUT96), .ZN(n447) );
  XNOR2_X1 U545 ( .A(n448), .B(n447), .ZN(n452) );
  XNOR2_X1 U546 ( .A(KEYINPUT97), .B(KEYINPUT5), .ZN(n450) );
  NAND2_X1 U547 ( .A1(G210), .A2(n486), .ZN(n449) );
  XNOR2_X1 U548 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U549 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U550 ( .A(n479), .B(n453), .ZN(n454) );
  XNOR2_X1 U551 ( .A(G472), .B(KEYINPUT98), .ZN(n457) );
  INV_X1 U552 ( .A(KEYINPUT72), .ZN(n456) );
  XNOR2_X1 U553 ( .A(n457), .B(n456), .ZN(n458) );
  INV_X1 U554 ( .A(n521), .ZN(n593) );
  NAND2_X1 U555 ( .A1(n460), .A2(n459), .ZN(n482) );
  NAND2_X1 U556 ( .A1(n482), .A2(G214), .ZN(n588) );
  INV_X1 U557 ( .A(n588), .ZN(n679) );
  XNOR2_X1 U558 ( .A(n461), .B(KEYINPUT14), .ZN(n465) );
  NAND2_X1 U559 ( .A1(G902), .A2(n465), .ZN(n462) );
  XNOR2_X1 U560 ( .A(KEYINPUT85), .B(n462), .ZN(n463) );
  NAND2_X1 U561 ( .A1(n463), .A2(G953), .ZN(n510) );
  XOR2_X1 U562 ( .A(KEYINPUT109), .B(n510), .Z(n464) );
  NOR2_X1 U563 ( .A1(n464), .A2(G900), .ZN(n469) );
  NAND2_X1 U564 ( .A1(n465), .A2(G952), .ZN(n466) );
  XNOR2_X1 U565 ( .A(n466), .B(KEYINPUT84), .ZN(n701) );
  INV_X1 U566 ( .A(n701), .ZN(n467) );
  NAND2_X1 U567 ( .A1(n467), .A2(n742), .ZN(n514) );
  INV_X1 U568 ( .A(n514), .ZN(n468) );
  NOR2_X1 U569 ( .A1(n469), .A2(n468), .ZN(n532) );
  INV_X1 U570 ( .A(n540), .ZN(n509) );
  XNOR2_X1 U571 ( .A(n471), .B(n470), .ZN(n475) );
  NAND2_X1 U572 ( .A1(n742), .A2(G224), .ZN(n473) );
  XNOR2_X1 U573 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n472) );
  XNOR2_X1 U574 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U575 ( .A(n475), .B(n474), .ZN(n477) );
  XNOR2_X1 U576 ( .A(n477), .B(n476), .ZN(n480) );
  XNOR2_X1 U577 ( .A(n505), .B(KEYINPUT16), .ZN(n478) );
  XNOR2_X1 U578 ( .A(n480), .B(n729), .ZN(n630) );
  INV_X1 U579 ( .A(n481), .ZN(n618) );
  NAND2_X1 U580 ( .A1(n482), .A2(G210), .ZN(n483) );
  XNOR2_X1 U581 ( .A(KEYINPUT12), .B(KEYINPUT101), .ZN(n484) );
  XNOR2_X1 U582 ( .A(n485), .B(n484), .ZN(n488) );
  NAND2_X1 U583 ( .A1(G214), .A2(n486), .ZN(n487) );
  XNOR2_X1 U584 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U585 ( .A(n489), .B(n735), .ZN(n495) );
  XNOR2_X1 U586 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U587 ( .A(n493), .B(n492), .Z(n494) );
  XNOR2_X1 U588 ( .A(n495), .B(n494), .ZN(n623) );
  NOR2_X1 U589 ( .A1(n623), .A2(G902), .ZN(n498) );
  XNOR2_X1 U590 ( .A(KEYINPUT102), .B(KEYINPUT13), .ZN(n496) );
  XOR2_X1 U591 ( .A(KEYINPUT104), .B(KEYINPUT7), .Z(n500) );
  XNOR2_X1 U592 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U593 ( .A(n348), .B(n502), .ZN(n507) );
  NAND2_X1 U594 ( .A1(G217), .A2(n503), .ZN(n504) );
  XOR2_X1 U595 ( .A(n505), .B(n504), .Z(n506) );
  XNOR2_X1 U596 ( .A(n507), .B(n506), .ZN(n710) );
  NAND2_X1 U597 ( .A1(n567), .A2(n569), .ZN(n556) );
  NOR2_X1 U598 ( .A1(n347), .A2(n556), .ZN(n508) );
  NAND2_X1 U599 ( .A1(n509), .A2(n508), .ZN(n611) );
  XNOR2_X1 U600 ( .A(n611), .B(G143), .ZN(G45) );
  INV_X1 U601 ( .A(n510), .ZN(n512) );
  INV_X1 U602 ( .A(G898), .ZN(n511) );
  NAND2_X1 U603 ( .A1(n512), .A2(n511), .ZN(n513) );
  NAND2_X1 U604 ( .A1(n514), .A2(n513), .ZN(n515) );
  INV_X1 U605 ( .A(n553), .ZN(n518) );
  NAND2_X1 U606 ( .A1(n518), .A2(n349), .ZN(n520) );
  XNOR2_X1 U607 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n519) );
  INV_X1 U608 ( .A(n544), .ZN(n684) );
  XNOR2_X1 U609 ( .A(n521), .B(KEYINPUT6), .ZN(n570) );
  NOR2_X1 U610 ( .A1(n684), .A2(n570), .ZN(n523) );
  XNOR2_X1 U611 ( .A(n522), .B(KEYINPUT1), .ZN(n549) );
  NAND2_X1 U612 ( .A1(n523), .A2(n687), .ZN(n524) );
  XOR2_X1 U613 ( .A(KEYINPUT78), .B(n524), .Z(n525) );
  NAND2_X1 U614 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U615 ( .A(n527), .B(KEYINPUT32), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n548), .B(G119), .ZN(G21) );
  INV_X1 U617 ( .A(n569), .ZN(n528) );
  NAND2_X1 U618 ( .A1(n528), .A2(n567), .ZN(n530) );
  INV_X1 U619 ( .A(KEYINPUT105), .ZN(n529) );
  XNOR2_X1 U620 ( .A(n530), .B(n529), .ZN(n663) );
  NAND2_X1 U621 ( .A1(n544), .A2(n683), .ZN(n531) );
  NOR2_X1 U622 ( .A1(n532), .A2(n531), .ZN(n592) );
  INV_X1 U623 ( .A(n592), .ZN(n533) );
  NOR2_X1 U624 ( .A1(n663), .A2(n533), .ZN(n534) );
  NAND2_X1 U625 ( .A1(n534), .A2(n570), .ZN(n599) );
  NOR2_X1 U626 ( .A1(n687), .A2(n599), .ZN(n535) );
  NAND2_X1 U627 ( .A1(n588), .A2(n535), .ZN(n536) );
  XNOR2_X1 U628 ( .A(n536), .B(KEYINPUT43), .ZN(n537) );
  NAND2_X1 U629 ( .A1(n347), .A2(n537), .ZN(n616) );
  XNOR2_X1 U630 ( .A(n616), .B(G140), .ZN(G42) );
  INV_X1 U631 ( .A(KEYINPUT74), .ZN(n538) );
  XNOR2_X1 U632 ( .A(n538), .B(KEYINPUT38), .ZN(n539) );
  XNOR2_X1 U633 ( .A(n347), .B(n539), .ZN(n676) );
  NOR2_X1 U634 ( .A1(n540), .A2(n676), .ZN(n541) );
  XNOR2_X1 U635 ( .A(n541), .B(KEYINPUT39), .ZN(n614) );
  NOR2_X1 U636 ( .A1(n614), .A2(n663), .ZN(n543) );
  XOR2_X1 U637 ( .A(KEYINPUT111), .B(KEYINPUT40), .Z(n542) );
  XOR2_X1 U638 ( .A(G131), .B(n598), .Z(G33) );
  INV_X1 U639 ( .A(n687), .ZN(n603) );
  NAND2_X1 U640 ( .A1(n544), .A2(n521), .ZN(n545) );
  NOR2_X2 U641 ( .A1(n571), .A2(n545), .ZN(n547) );
  XNOR2_X1 U642 ( .A(n547), .B(n546), .ZN(n644) );
  NAND2_X1 U643 ( .A1(n644), .A2(n548), .ZN(n580) );
  XNOR2_X1 U644 ( .A(n580), .B(KEYINPUT81), .ZN(n559) );
  INV_X1 U645 ( .A(KEYINPUT34), .ZN(n555) );
  NAND2_X1 U646 ( .A1(n561), .A2(n570), .ZN(n552) );
  NOR2_X1 U647 ( .A1(n674), .A2(n565), .ZN(n554) );
  XNOR2_X1 U648 ( .A(n555), .B(n554), .ZN(n557) );
  XNOR2_X2 U649 ( .A(n558), .B(KEYINPUT35), .ZN(n747) );
  NAND2_X1 U650 ( .A1(n559), .A2(n747), .ZN(n560) );
  NAND2_X1 U651 ( .A1(n561), .A2(n593), .ZN(n563) );
  INV_X1 U652 ( .A(KEYINPUT99), .ZN(n562) );
  NAND2_X1 U653 ( .A1(n564), .A2(n521), .ZN(n566) );
  OR2_X1 U654 ( .A1(n566), .A2(n565), .ZN(n653) );
  INV_X1 U655 ( .A(n567), .ZN(n568) );
  NAND2_X1 U656 ( .A1(n569), .A2(n568), .ZN(n668) );
  AND2_X1 U657 ( .A1(n663), .A2(n668), .ZN(n675) );
  OR2_X1 U658 ( .A1(n571), .A2(n570), .ZN(n573) );
  INV_X1 U659 ( .A(KEYINPUT80), .ZN(n572) );
  XNOR2_X1 U660 ( .A(n573), .B(n572), .ZN(n574) );
  AND2_X1 U661 ( .A1(n574), .A2(n684), .ZN(n650) );
  INV_X1 U662 ( .A(n650), .ZN(n575) );
  NAND2_X1 U663 ( .A1(n576), .A2(n575), .ZN(n579) );
  AND2_X1 U664 ( .A1(n580), .A2(KEYINPUT44), .ZN(n577) );
  NOR2_X1 U665 ( .A1(n577), .A2(KEYINPUT64), .ZN(n578) );
  NOR2_X1 U666 ( .A1(n579), .A2(n578), .ZN(n585) );
  AND2_X1 U667 ( .A1(n580), .A2(KEYINPUT64), .ZN(n581) );
  NOR2_X1 U668 ( .A1(n581), .A2(KEYINPUT71), .ZN(n582) );
  NAND2_X1 U669 ( .A1(n747), .A2(n582), .ZN(n583) );
  NAND2_X1 U670 ( .A1(n583), .A2(KEYINPUT44), .ZN(n584) );
  NAND2_X1 U671 ( .A1(n588), .A2(n681), .ZN(n591) );
  NAND2_X1 U672 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U673 ( .A(KEYINPUT28), .B(n594), .Z(n596) );
  NAND2_X1 U674 ( .A1(n596), .A2(n595), .ZN(n607) );
  NOR2_X1 U675 ( .A1(n703), .A2(n607), .ZN(n597) );
  XNOR2_X1 U676 ( .A(n597), .B(KEYINPUT42), .ZN(n748) );
  XOR2_X1 U677 ( .A(KEYINPUT113), .B(n599), .Z(n601) );
  NOR2_X1 U678 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U679 ( .A(KEYINPUT36), .B(n602), .Z(n604) );
  NOR2_X1 U680 ( .A1(n604), .A2(n603), .ZN(n670) );
  INV_X1 U681 ( .A(n605), .ZN(n606) );
  NOR2_X1 U682 ( .A1(n607), .A2(n606), .ZN(n661) );
  NOR2_X1 U683 ( .A1(KEYINPUT65), .A2(n675), .ZN(n608) );
  NAND2_X1 U684 ( .A1(n661), .A2(n608), .ZN(n609) );
  XOR2_X1 U685 ( .A(KEYINPUT47), .B(n609), .Z(n610) );
  NAND2_X1 U686 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U687 ( .A1(n670), .A2(n612), .ZN(n613) );
  NOR2_X1 U688 ( .A1(n614), .A2(n668), .ZN(n615) );
  XNOR2_X1 U689 ( .A(n615), .B(KEYINPUT114), .ZN(n749) );
  INV_X1 U690 ( .A(n749), .ZN(n617) );
  INV_X1 U691 ( .A(n672), .ZN(n619) );
  NAND2_X1 U692 ( .A1(n619), .A2(KEYINPUT2), .ZN(n645) );
  AND2_X1 U693 ( .A1(G475), .A2(n645), .ZN(n622) );
  NAND2_X1 U694 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U695 ( .A1(n620), .A2(KEYINPUT79), .ZN(n621) );
  NAND2_X1 U696 ( .A1(n622), .A2(n647), .ZN(n625) );
  XOR2_X1 U697 ( .A(KEYINPUT59), .B(n623), .Z(n624) );
  XNOR2_X1 U698 ( .A(n625), .B(n624), .ZN(n627) );
  INV_X1 U699 ( .A(G952), .ZN(n626) );
  AND2_X1 U700 ( .A1(n626), .A2(G953), .ZN(n718) );
  XNOR2_X1 U701 ( .A(n628), .B(KEYINPUT60), .ZN(G60) );
  XOR2_X1 U702 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n629) );
  XNOR2_X1 U703 ( .A(n630), .B(n629), .ZN(n631) );
  XNOR2_X1 U704 ( .A(n632), .B(n631), .ZN(n633) );
  XOR2_X1 U705 ( .A(KEYINPUT119), .B(KEYINPUT56), .Z(n634) );
  XNOR2_X1 U706 ( .A(n635), .B(n634), .ZN(G51) );
  XOR2_X1 U707 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n637) );
  XNOR2_X1 U708 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n636) );
  XNOR2_X1 U709 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U710 ( .A(n639), .B(n638), .ZN(n640) );
  XNOR2_X1 U711 ( .A(n641), .B(n640), .ZN(n642) );
  XNOR2_X1 U712 ( .A(n643), .B(KEYINPUT122), .ZN(G54) );
  XNOR2_X1 U713 ( .A(n644), .B(G110), .ZN(G12) );
  AND2_X1 U714 ( .A1(G472), .A2(n645), .ZN(n646) );
  NAND2_X1 U715 ( .A1(n647), .A2(n646), .ZN(n649) );
  XNOR2_X1 U716 ( .A(G101), .B(n650), .ZN(n651) );
  XNOR2_X1 U717 ( .A(n651), .B(KEYINPUT115), .ZN(G3) );
  NOR2_X1 U718 ( .A1(n653), .A2(n663), .ZN(n652) );
  XOR2_X1 U719 ( .A(G104), .B(n652), .Z(G6) );
  NOR2_X1 U720 ( .A1(n653), .A2(n668), .ZN(n655) );
  XNOR2_X1 U721 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n654) );
  XNOR2_X1 U722 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U723 ( .A(G107), .B(n656), .ZN(G9) );
  XOR2_X1 U724 ( .A(G128), .B(KEYINPUT29), .Z(n659) );
  INV_X1 U725 ( .A(n668), .ZN(n657) );
  NAND2_X1 U726 ( .A1(n661), .A2(n657), .ZN(n658) );
  XNOR2_X1 U727 ( .A(n659), .B(n658), .ZN(G30) );
  INV_X1 U728 ( .A(n663), .ZN(n660) );
  NAND2_X1 U729 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U730 ( .A(n662), .B(G146), .ZN(G48) );
  NOR2_X1 U731 ( .A1(n663), .A2(n667), .ZN(n665) );
  XNOR2_X1 U732 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n664) );
  XNOR2_X1 U733 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U734 ( .A(G113), .B(n666), .ZN(G15) );
  NOR2_X1 U735 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U736 ( .A(G116), .B(n669), .Z(G18) );
  XNOR2_X1 U737 ( .A(G125), .B(n670), .ZN(n671) );
  XNOR2_X1 U738 ( .A(n671), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U739 ( .A(KEYINPUT2), .B(n673), .Z(n707) );
  NOR2_X1 U740 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U741 ( .A1(n586), .A2(n677), .ZN(n678) );
  NOR2_X1 U742 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U743 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U744 ( .A1(n702), .A2(n682), .ZN(n698) );
  NOR2_X1 U745 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U746 ( .A(n685), .B(KEYINPUT49), .ZN(n686) );
  NAND2_X1 U747 ( .A1(n686), .A2(n521), .ZN(n691) );
  NOR2_X1 U748 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U749 ( .A(n689), .B(KEYINPUT50), .ZN(n690) );
  OR2_X1 U750 ( .A1(n691), .A2(n690), .ZN(n693) );
  NAND2_X1 U751 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U752 ( .A(n694), .B(KEYINPUT51), .ZN(n695) );
  XNOR2_X1 U753 ( .A(n695), .B(KEYINPUT118), .ZN(n696) );
  NOR2_X1 U754 ( .A1(n703), .A2(n696), .ZN(n697) );
  NOR2_X1 U755 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U756 ( .A(n699), .B(KEYINPUT52), .ZN(n700) );
  NOR2_X1 U757 ( .A1(n701), .A2(n700), .ZN(n705) );
  NOR2_X1 U758 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U759 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U760 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U761 ( .A1(n708), .A2(G953), .ZN(n709) );
  XNOR2_X1 U762 ( .A(n709), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U763 ( .A(n711), .B(n710), .ZN(n712) );
  NOR2_X1 U764 ( .A1(n718), .A2(n712), .ZN(G63) );
  NAND2_X1 U765 ( .A1(n713), .A2(G217), .ZN(n716) );
  XOR2_X1 U766 ( .A(n714), .B(KEYINPUT123), .Z(n715) );
  XNOR2_X1 U767 ( .A(n716), .B(n715), .ZN(n717) );
  NOR2_X1 U768 ( .A1(n718), .A2(n717), .ZN(G66) );
  BUF_X1 U769 ( .A(n719), .Z(n720) );
  NAND2_X1 U770 ( .A1(n720), .A2(n742), .ZN(n726) );
  NAND2_X1 U771 ( .A1(G224), .A2(G953), .ZN(n721) );
  XNOR2_X1 U772 ( .A(n721), .B(KEYINPUT61), .ZN(n722) );
  XNOR2_X1 U773 ( .A(KEYINPUT124), .B(n722), .ZN(n723) );
  NAND2_X1 U774 ( .A1(n723), .A2(G898), .ZN(n724) );
  XOR2_X1 U775 ( .A(KEYINPUT125), .B(n724), .Z(n725) );
  NAND2_X1 U776 ( .A1(n726), .A2(n725), .ZN(n733) );
  XNOR2_X1 U777 ( .A(n727), .B(G101), .ZN(n728) );
  XNOR2_X1 U778 ( .A(n729), .B(n728), .ZN(n731) );
  NOR2_X1 U779 ( .A1(G898), .A2(n742), .ZN(n730) );
  NOR2_X1 U780 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U781 ( .A(n733), .B(n732), .ZN(G69) );
  XNOR2_X1 U782 ( .A(KEYINPUT4), .B(KEYINPUT126), .ZN(n734) );
  XNOR2_X1 U783 ( .A(n735), .B(n734), .ZN(n736) );
  XNOR2_X1 U784 ( .A(n737), .B(n736), .ZN(n740) );
  XOR2_X1 U785 ( .A(G227), .B(n740), .Z(n738) );
  NOR2_X1 U786 ( .A1(n742), .A2(n738), .ZN(n739) );
  NAND2_X1 U787 ( .A1(n739), .A2(G900), .ZN(n745) );
  XNOR2_X1 U788 ( .A(n741), .B(n740), .ZN(n743) );
  NAND2_X1 U789 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U790 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U791 ( .A(KEYINPUT127), .B(n746), .ZN(G72) );
  XNOR2_X1 U792 ( .A(n747), .B(G122), .ZN(G24) );
  XOR2_X1 U793 ( .A(G137), .B(n748), .Z(G39) );
  XOR2_X1 U794 ( .A(G134), .B(n749), .Z(G36) );
endmodule

