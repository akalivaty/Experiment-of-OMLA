//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 1 1 1 1 1 1 0 1 0 0 0 1 1 0 1 1 1 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004;
  INV_X1    g000(.A(KEYINPUT76), .ZN(new_n187));
  INV_X1    g001(.A(G107), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(G104), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT3), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n188), .A2(G104), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n193));
  NAND4_X1  g007(.A1(new_n187), .A2(new_n193), .A3(new_n188), .A4(G104), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n190), .A2(new_n192), .A3(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G101), .ZN(new_n196));
  INV_X1    g010(.A(G101), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n190), .A2(new_n197), .A3(new_n192), .A4(new_n194), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(KEYINPUT4), .A3(new_n198), .ZN(new_n199));
  XOR2_X1   g013(.A(G116), .B(G119), .Z(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT2), .B(G113), .ZN(new_n201));
  XNOR2_X1  g015(.A(new_n200), .B(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT4), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n195), .A2(new_n203), .A3(G101), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n199), .A2(new_n202), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G104), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(G107), .ZN(new_n207));
  OAI21_X1  g021(.A(G101), .B1(new_n191), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n198), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  OR2_X1    g024(.A1(new_n200), .A2(new_n201), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT5), .ZN(new_n212));
  INV_X1    g026(.A(G119), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n213), .A3(G116), .ZN(new_n214));
  OAI211_X1 g028(.A(G113), .B(new_n214), .C1(new_n200), .C2(new_n212), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n210), .A2(new_n211), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n205), .A2(new_n216), .ZN(new_n217));
  XOR2_X1   g031(.A(G110), .B(G122), .Z(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n218), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n205), .A2(new_n216), .A3(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n219), .A2(KEYINPUT6), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT0), .ZN(new_n223));
  INV_X1    g037(.A(G128), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G143), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT64), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT64), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G143), .ZN(new_n229));
  INV_X1    g043(.A(G146), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n227), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(KEYINPUT65), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT65), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G146), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n232), .A2(new_n234), .A3(new_n226), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n225), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n223), .A2(new_n224), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n232), .A2(new_n234), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G143), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n228), .A2(G143), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n226), .A2(KEYINPUT64), .ZN(new_n242));
  OAI21_X1  g056(.A(G146), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n240), .A2(new_n243), .A3(new_n225), .ZN(new_n244));
  OR2_X1    g058(.A1(KEYINPUT74), .A2(G125), .ZN(new_n245));
  NAND2_X1  g059(.A1(KEYINPUT74), .A2(G125), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n238), .A2(new_n244), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n231), .A2(new_n235), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT1), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n251), .B1(new_n239), .B2(G143), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n250), .B1(new_n252), .B2(new_n224), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n240), .A2(new_n243), .A3(new_n251), .A4(G128), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n248), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n249), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G224), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(G953), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n258), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n260), .B1(new_n249), .B2(new_n255), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n217), .A2(new_n263), .A3(new_n218), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n222), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  OAI211_X1 g079(.A(KEYINPUT7), .B(new_n260), .C1(new_n249), .C2(new_n255), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n266), .A2(new_n221), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n215), .A2(new_n211), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n209), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n216), .A2(new_n269), .ZN(new_n270));
  XOR2_X1   g084(.A(new_n218), .B(KEYINPUT8), .Z(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT7), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n256), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n267), .A2(new_n259), .A3(new_n272), .A4(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G902), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n265), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(G210), .B1(G237), .B2(G902), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n265), .A2(new_n275), .A3(new_n276), .A4(new_n278), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT79), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT79), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(G214), .B1(G237), .B2(G902), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  OR2_X1    g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G469), .ZN(new_n290));
  XNOR2_X1  g104(.A(G110), .B(G140), .ZN(new_n291));
  INV_X1    g105(.A(G953), .ZN(new_n292));
  AND2_X1   g106(.A1(new_n292), .A2(G227), .ZN(new_n293));
  XOR2_X1   g107(.A(new_n291), .B(new_n293), .Z(new_n294));
  AOI21_X1  g108(.A(new_n230), .B1(new_n227), .B2(new_n229), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n295), .B1(G143), .B2(new_n239), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n296), .A2(new_n225), .B1(new_n236), .B2(new_n237), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n297), .A2(new_n199), .A3(new_n204), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT77), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n297), .A2(new_n199), .A3(KEYINPUT77), .A4(new_n204), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT64), .B(G143), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n251), .B1(new_n303), .B2(new_n230), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT65), .B(G146), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n305), .A2(new_n226), .ZN(new_n306));
  OAI22_X1  g120(.A1(new_n304), .A2(new_n224), .B1(new_n306), .B2(new_n295), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n209), .B1(new_n307), .B2(new_n254), .ZN(new_n308));
  OR2_X1    g122(.A1(new_n308), .A2(KEYINPUT10), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n253), .A2(new_n254), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(KEYINPUT10), .A3(new_n210), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n302), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G134), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT66), .B1(new_n313), .B2(G137), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT11), .ZN(new_n315));
  INV_X1    g129(.A(G137), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n316), .A2(G134), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT11), .ZN(new_n319));
  OAI211_X1 g133(.A(KEYINPUT66), .B(new_n319), .C1(new_n313), .C2(G137), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n315), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G131), .ZN(new_n322));
  INV_X1    g136(.A(G131), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n315), .A2(new_n323), .A3(new_n318), .A4(new_n320), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n312), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n325), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n302), .A2(new_n327), .A3(new_n309), .A4(new_n311), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n294), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  AND3_X1   g143(.A1(new_n253), .A2(new_n254), .A3(new_n209), .ZN(new_n330));
  OAI211_X1 g144(.A(KEYINPUT12), .B(new_n325), .C1(new_n330), .C2(new_n308), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT78), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n224), .B1(new_n231), .B2(KEYINPUT1), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n254), .B1(new_n296), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n210), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n253), .A2(new_n254), .A3(new_n209), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n338), .A2(KEYINPUT78), .A3(KEYINPUT12), .A4(new_n325), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n325), .B1(new_n330), .B2(new_n308), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT12), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n333), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  AND3_X1   g157(.A1(new_n343), .A2(new_n328), .A3(new_n294), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n290), .B(new_n276), .C1(new_n329), .C2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(G469), .A2(G902), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n343), .A2(new_n328), .ZN(new_n347));
  INV_X1    g161(.A(new_n294), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n326), .A2(new_n328), .A3(new_n294), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(new_n350), .A3(G469), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n345), .A2(new_n346), .A3(new_n351), .ZN(new_n352));
  XOR2_X1   g166(.A(KEYINPUT9), .B(G234), .Z(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(G221), .B1(new_n354), .B2(G902), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G116), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G122), .ZN(new_n358));
  INV_X1    g172(.A(G122), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G116), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G107), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n358), .A2(new_n360), .A3(new_n188), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT82), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n226), .A2(G128), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  OAI211_X1 g181(.A(KEYINPUT13), .B(new_n367), .C1(new_n303), .C2(new_n224), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n227), .A2(new_n229), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT13), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n370), .A3(G128), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n368), .A2(G134), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n369), .A2(G128), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(new_n313), .A3(new_n367), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT82), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n362), .A2(new_n375), .A3(new_n363), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n365), .A2(new_n372), .A3(new_n374), .A4(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT14), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n359), .A2(G116), .ZN(new_n379));
  AOI22_X1  g193(.A1(new_n378), .A2(new_n379), .B1(new_n360), .B2(KEYINPUT83), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n378), .A2(new_n357), .A3(KEYINPUT83), .A4(G122), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n381), .B1(new_n378), .B2(new_n379), .ZN(new_n382));
  OAI21_X1  g196(.A(G107), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n313), .B1(new_n373), .B2(new_n367), .ZN(new_n384));
  AOI211_X1 g198(.A(G134), .B(new_n366), .C1(new_n369), .C2(G128), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n383), .B(new_n363), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n377), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n353), .A2(G217), .A3(new_n292), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT84), .ZN(new_n390));
  INV_X1    g204(.A(new_n388), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n377), .A2(new_n386), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n389), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT85), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n387), .A2(KEYINPUT84), .A3(new_n388), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n393), .A2(new_n394), .A3(new_n276), .A4(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G478), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n397), .A2(KEYINPUT15), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n396), .A2(new_n398), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT86), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  OR2_X1    g217(.A1(new_n396), .A2(new_n398), .ZN(new_n404));
  AOI21_X1  g218(.A(KEYINPUT86), .B1(new_n404), .B2(new_n399), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G475), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT80), .ZN(new_n408));
  INV_X1    g222(.A(G214), .ZN(new_n409));
  NOR3_X1   g223(.A1(new_n409), .A2(G237), .A3(G953), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n303), .A2(new_n410), .ZN(new_n411));
  NOR4_X1   g225(.A1(new_n226), .A2(new_n409), .A3(G237), .A4(G953), .ZN(new_n412));
  OAI21_X1  g226(.A(G131), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NOR3_X1   g228(.A1(new_n411), .A2(G131), .A3(new_n412), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n408), .B(KEYINPUT18), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n411), .A2(new_n412), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n408), .A2(KEYINPUT18), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n245), .A2(G140), .A3(new_n246), .ZN(new_n420));
  OR2_X1    g234(.A1(G125), .A2(G140), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n420), .A2(KEYINPUT81), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(KEYINPUT81), .B1(new_n420), .B2(new_n421), .ZN(new_n423));
  OAI21_X1  g237(.A(G146), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(G125), .B(G140), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n239), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n416), .A2(new_n419), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n417), .A2(new_n323), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT17), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n429), .A2(new_n430), .A3(new_n413), .ZN(new_n431));
  NOR3_X1   g245(.A1(new_n247), .A2(KEYINPUT16), .A3(G140), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n420), .A2(new_n421), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n432), .B1(KEYINPUT16), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G146), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n414), .A2(KEYINPUT17), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n433), .A2(KEYINPUT16), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n230), .B1(new_n437), .B2(new_n432), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n431), .A2(new_n435), .A3(new_n436), .A4(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(G113), .B(G122), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n440), .B(new_n206), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n428), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  AOI22_X1  g257(.A1(G146), .A2(new_n434), .B1(new_n429), .B2(new_n413), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT19), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n422), .A2(new_n423), .A3(new_n445), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n425), .A2(KEYINPUT19), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n239), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n441), .B1(new_n449), .B2(new_n428), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n407), .B(new_n276), .C1(new_n443), .C2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT20), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n449), .A2(new_n428), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n442), .B1(new_n454), .B2(new_n441), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n455), .A2(KEYINPUT20), .A3(new_n407), .A4(new_n276), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n441), .B1(new_n428), .B2(new_n439), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n276), .B1(new_n443), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G475), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n453), .A2(new_n456), .A3(new_n459), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n292), .A2(G952), .ZN(new_n461));
  NAND2_X1  g275(.A1(G234), .A2(G237), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  XOR2_X1   g278(.A(KEYINPUT21), .B(G898), .Z(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n462), .A2(G902), .A3(G953), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n464), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  NOR3_X1   g283(.A1(new_n406), .A2(new_n460), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NOR3_X1   g285(.A1(new_n289), .A2(new_n356), .A3(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(KEYINPUT75), .A2(KEYINPUT25), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT23), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n474), .B1(G119), .B2(new_n224), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n213), .A2(KEYINPUT23), .A3(G128), .ZN(new_n476));
  OAI22_X1  g290(.A1(new_n475), .A2(new_n476), .B1(G119), .B2(new_n224), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(G110), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT72), .B1(new_n224), .B2(G119), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT72), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n480), .A2(new_n213), .A3(G128), .ZN(new_n481));
  AOI22_X1  g295(.A1(new_n479), .A2(new_n481), .B1(G119), .B2(new_n224), .ZN(new_n482));
  XOR2_X1   g296(.A(KEYINPUT24), .B(G110), .Z(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n484), .B(KEYINPUT73), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n434), .A2(G146), .ZN(new_n486));
  NOR3_X1   g300(.A1(new_n437), .A2(new_n230), .A3(new_n432), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n478), .B(new_n485), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  OAI22_X1  g302(.A1(new_n477), .A2(G110), .B1(new_n482), .B2(new_n483), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n435), .A2(new_n426), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n292), .A2(G221), .A3(G234), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(KEYINPUT22), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(G137), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n488), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n493), .B1(new_n488), .B2(new_n490), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n473), .B1(new_n496), .B2(new_n276), .ZN(new_n497));
  INV_X1    g311(.A(new_n473), .ZN(new_n498));
  NOR4_X1   g312(.A1(new_n494), .A2(new_n495), .A3(G902), .A4(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(G217), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n501), .B1(G234), .B2(new_n276), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n502), .A2(G902), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n496), .A2(new_n504), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n297), .A2(new_n325), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n313), .A2(G137), .ZN(new_n509));
  OAI21_X1  g323(.A(G131), .B1(new_n317), .B2(new_n509), .ZN(new_n510));
  AND2_X1   g324(.A1(new_n324), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(KEYINPUT1), .B1(new_n305), .B2(new_n226), .ZN(new_n512));
  AOI22_X1  g326(.A1(new_n512), .A2(G128), .B1(new_n231), .B2(new_n235), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n251), .A2(G128), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n306), .A2(new_n295), .A3(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n511), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n202), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n508), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT67), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n508), .A2(new_n516), .A3(KEYINPUT67), .A4(new_n517), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n520), .A2(KEYINPUT28), .A3(new_n521), .ZN(new_n522));
  AOI22_X1  g336(.A1(new_n310), .A2(new_n511), .B1(new_n297), .B2(new_n325), .ZN(new_n523));
  OR2_X1    g337(.A1(new_n523), .A2(new_n517), .ZN(new_n524));
  AOI21_X1  g338(.A(KEYINPUT28), .B1(new_n523), .B2(new_n517), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n522), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n528));
  INV_X1    g342(.A(G210), .ZN(new_n529));
  NOR3_X1   g343(.A1(new_n529), .A2(G237), .A3(G953), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n528), .B(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(KEYINPUT26), .B(G101), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n527), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT30), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n508), .A2(new_n535), .A3(new_n516), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n535), .B1(new_n508), .B2(new_n516), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n202), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n520), .A2(new_n521), .ZN(new_n539));
  INV_X1    g353(.A(new_n533), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT31), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT69), .B(KEYINPUT31), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n538), .A2(new_n539), .A3(new_n540), .A4(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n534), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT32), .ZN(new_n546));
  NOR2_X1   g360(.A1(G472), .A2(G902), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n546), .B1(new_n545), .B2(new_n547), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(G472), .ZN(new_n551));
  AOI21_X1  g365(.A(KEYINPUT67), .B1(new_n523), .B2(new_n517), .ZN(new_n552));
  INV_X1    g366(.A(new_n521), .ZN(new_n553));
  OAI21_X1  g367(.A(KEYINPUT70), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT70), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n520), .A2(new_n555), .A3(new_n521), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n554), .A2(new_n524), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n525), .B1(new_n557), .B2(KEYINPUT28), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT29), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n533), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(G902), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n538), .A2(new_n539), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n533), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n563), .B(new_n559), .C1(new_n533), .C2(new_n527), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n551), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(KEYINPUT71), .B1(new_n550), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n545), .A2(new_n547), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT32), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n557), .A2(KEYINPUT28), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n526), .ZN(new_n572));
  INV_X1    g386(.A(new_n560), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n564), .B(new_n276), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(G472), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT71), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n570), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n507), .B1(new_n566), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n472), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT87), .B(G101), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n579), .B(new_n580), .ZN(G3));
  INV_X1    g395(.A(new_n355), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n507), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n567), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n551), .B1(new_n545), .B2(new_n276), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n583), .A2(new_n586), .A3(new_n352), .ZN(new_n587));
  INV_X1    g401(.A(new_n460), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT33), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n393), .A2(new_n589), .A3(new_n395), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n389), .A2(KEYINPUT33), .A3(new_n392), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n397), .A2(G902), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n393), .A2(new_n276), .A3(new_n395), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n592), .A2(new_n593), .B1(new_n397), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n588), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n288), .B1(new_n280), .B2(new_n281), .ZN(new_n598));
  INV_X1    g412(.A(new_n469), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n587), .A2(new_n601), .ZN(new_n602));
  XOR2_X1   g416(.A(KEYINPUT34), .B(G104), .Z(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT88), .B(KEYINPUT89), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G6));
  INV_X1    g420(.A(new_n600), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n607), .A2(KEYINPUT90), .A3(new_n588), .A4(new_n406), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT90), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n406), .A2(new_n588), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n609), .B1(new_n610), .B2(new_n600), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n587), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT35), .B(G107), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G9));
  NAND2_X1  g429(.A1(new_n488), .A2(new_n490), .ZN(new_n616));
  INV_X1    g430(.A(new_n493), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n616), .B1(KEYINPUT36), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n617), .A2(KEYINPUT36), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n488), .A2(new_n490), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n618), .A2(new_n504), .A3(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT91), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n618), .A2(KEYINPUT91), .A3(new_n504), .A4(new_n620), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n500), .B2(new_n502), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(KEYINPUT92), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n586), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT93), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT93), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n627), .A2(new_n630), .A3(new_n586), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n472), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(new_n632), .B(KEYINPUT37), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G110), .ZN(G12));
  NAND2_X1  g448(.A1(new_n566), .A2(new_n577), .ZN(new_n635));
  INV_X1    g449(.A(G900), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n464), .B1(new_n468), .B2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n406), .A2(new_n588), .A3(new_n598), .A4(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT94), .ZN(new_n640));
  OR2_X1    g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n356), .B1(new_n639), .B2(new_n640), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n635), .A2(new_n627), .A3(new_n641), .A4(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G128), .ZN(G30));
  INV_X1    g458(.A(new_n406), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n645), .A2(new_n588), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT95), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n286), .B(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT38), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n286), .B(KEYINPUT95), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(KEYINPUT38), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n647), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n276), .B1(new_n557), .B2(new_n540), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n562), .A2(new_n540), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g471(.A(G472), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n570), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT96), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n637), .B(KEYINPUT97), .ZN(new_n661));
  XOR2_X1   g475(.A(new_n661), .B(KEYINPUT39), .Z(new_n662));
  AND3_X1   g476(.A1(new_n352), .A2(new_n355), .A3(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT40), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n288), .B1(new_n663), .B2(new_n664), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n654), .A2(new_n626), .A3(new_n666), .A4(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(new_n303), .ZN(G45));
  INV_X1    g483(.A(new_n598), .ZN(new_n670));
  INV_X1    g484(.A(new_n595), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n671), .A2(new_n460), .A3(new_n638), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n356), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n635), .A2(new_n627), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G146), .ZN(G48));
  OAI21_X1  g489(.A(new_n276), .B1(new_n329), .B2(new_n344), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(G469), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n677), .A2(new_n355), .A3(new_n345), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT98), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n677), .A2(KEYINPUT98), .A3(new_n355), .A4(new_n345), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n635), .A2(new_n682), .A3(new_n506), .A4(new_n601), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT41), .B(G113), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G15));
  NAND3_X1  g499(.A1(new_n578), .A2(new_n612), .A3(new_n682), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G116), .ZN(G18));
  NOR2_X1   g501(.A1(new_n678), .A2(new_n670), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n635), .A2(new_n470), .A3(new_n627), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G119), .ZN(G21));
  AOI21_X1  g504(.A(new_n600), .B1(new_n680), .B2(new_n681), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n572), .A2(KEYINPUT99), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT99), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n558), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n692), .A2(new_n533), .A3(new_n694), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n542), .A2(new_n544), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n585), .B1(new_n697), .B2(new_n547), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n691), .A2(new_n698), .A3(new_n506), .A4(new_n646), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G122), .ZN(G24));
  INV_X1    g514(.A(new_n626), .ZN(new_n701));
  INV_X1    g515(.A(new_n672), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n698), .A2(new_n701), .A3(new_n702), .A4(new_n688), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G125), .ZN(G27));
  NAND3_X1  g518(.A1(new_n283), .A2(new_n287), .A3(new_n285), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n705), .A2(new_n356), .A3(new_n672), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n550), .A2(new_n565), .A3(KEYINPUT71), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n576), .B1(new_n570), .B2(new_n575), .ZN(new_n708));
  OAI211_X1 g522(.A(new_n706), .B(new_n506), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT100), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT42), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n578), .A2(KEYINPUT100), .A3(new_n706), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n570), .B(KEYINPUT101), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n507), .B1(new_n715), .B2(new_n575), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(KEYINPUT42), .A3(new_n706), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(KEYINPUT102), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT102), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n714), .A2(new_n720), .A3(new_n717), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G131), .ZN(G33));
  NAND2_X1  g537(.A1(new_n588), .A2(new_n638), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n645), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n705), .A2(new_n356), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n578), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G134), .ZN(G36));
  INV_X1    g542(.A(KEYINPUT103), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT43), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n730), .B1(new_n460), .B2(new_n595), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n460), .A2(new_n595), .A3(new_n730), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n729), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n588), .A2(new_n671), .A3(KEYINPUT43), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(KEYINPUT103), .A3(new_n731), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g551(.A(KEYINPUT104), .B1(new_n586), .B2(new_n626), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT104), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n701), .B(new_n739), .C1(new_n584), .C2(new_n585), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n737), .A2(new_n738), .A3(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n349), .A2(new_n350), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT45), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n349), .A2(new_n350), .A3(KEYINPUT45), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(G469), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(KEYINPUT46), .B1(new_n748), .B2(new_n346), .ZN(new_n749));
  INV_X1    g563(.A(new_n345), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n748), .A2(KEYINPUT46), .A3(new_n346), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n582), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n743), .A2(new_n662), .A3(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n737), .A2(new_n738), .A3(KEYINPUT44), .A4(new_n740), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT105), .ZN(new_n756));
  INV_X1    g570(.A(new_n705), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n755), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n756), .B1(new_n755), .B2(new_n757), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n754), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(new_n316), .ZN(G39));
  INV_X1    g575(.A(KEYINPUT47), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n751), .A2(new_n752), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n762), .B1(new_n763), .B2(new_n582), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n753), .A2(KEYINPUT47), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n635), .A2(new_n506), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n766), .A2(new_n702), .A3(new_n757), .A4(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(KEYINPUT106), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G140), .ZN(G42));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT50), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n698), .A2(new_n506), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n463), .B1(new_n735), .B2(new_n731), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(new_n653), .A3(new_n651), .ZN(new_n776));
  INV_X1    g590(.A(new_n678), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n288), .ZN(new_n778));
  XOR2_X1   g592(.A(new_n778), .B(KEYINPUT112), .Z(new_n779));
  OAI21_X1  g593(.A(new_n772), .B1(new_n776), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n651), .A2(new_n653), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n773), .A2(new_n774), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n779), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(KEYINPUT50), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n780), .A2(new_n785), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n757), .A2(new_n774), .A3(new_n777), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n787), .A2(new_n701), .A3(new_n698), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n660), .A2(new_n464), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n507), .A2(new_n705), .A3(new_n678), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n789), .A2(new_n588), .A3(new_n595), .A4(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n786), .A2(new_n788), .A3(new_n791), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n677), .A2(new_n345), .ZN(new_n793));
  XOR2_X1   g607(.A(new_n793), .B(KEYINPUT111), .Z(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n582), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n764), .A2(new_n765), .A3(new_n795), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n796), .A2(new_n757), .A3(new_n775), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n771), .B1(new_n792), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n716), .A2(new_n787), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT48), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n796), .A2(KEYINPUT113), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n796), .A2(KEYINPUT113), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n801), .A2(new_n757), .A3(new_n775), .A4(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n791), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n804), .B1(new_n780), .B2(new_n785), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n803), .A2(new_n805), .A3(KEYINPUT51), .A4(new_n788), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n798), .A2(new_n461), .A3(new_n800), .A4(new_n806), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n782), .A2(new_n670), .A3(new_n678), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n789), .A2(new_n596), .A3(new_n790), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n406), .A2(new_n460), .A3(new_n598), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n811), .B1(new_n570), .B2(new_n658), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n352), .A2(new_n626), .A3(new_n355), .A4(new_n638), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT108), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n813), .A2(new_n814), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n812), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n643), .A2(new_n674), .A3(new_n703), .A4(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n818), .A2(new_n819), .ZN(new_n821));
  OAI21_X1  g635(.A(KEYINPUT109), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n643), .A2(new_n703), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n823), .A2(KEYINPUT52), .A3(new_n674), .A4(new_n817), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT109), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n818), .A2(new_n819), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n822), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n698), .A2(new_n701), .A3(new_n702), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n578), .A2(new_n725), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n400), .A2(new_n401), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n635), .A2(new_n831), .A3(new_n627), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n829), .B(new_n830), .C1(new_n724), .C2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n726), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n460), .A2(new_n831), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n596), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n289), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n587), .A2(new_n837), .A3(new_n599), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n632), .A2(new_n579), .A3(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n686), .A2(new_n689), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n683), .A2(new_n699), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT107), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n840), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n686), .A2(new_n689), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT107), .B1(new_n845), .B2(new_n841), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n839), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n828), .A2(new_n722), .A3(new_n834), .A4(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT53), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n722), .A2(new_n834), .A3(new_n847), .ZN(new_n850));
  AOI21_X1  g664(.A(KEYINPUT53), .B1(new_n824), .B2(new_n826), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n849), .A2(KEYINPUT54), .A3(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT53), .ZN(new_n854));
  INV_X1    g668(.A(new_n828), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n722), .A2(new_n847), .A3(new_n834), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT54), .ZN(new_n858));
  INV_X1    g672(.A(new_n839), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n859), .B(new_n718), .C1(new_n820), .C2(new_n821), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n834), .A2(KEYINPUT53), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n840), .A2(new_n842), .A3(KEYINPUT110), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT110), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n863), .B1(new_n845), .B2(new_n841), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n860), .A2(new_n861), .A3(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n857), .A2(new_n858), .A3(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n809), .A2(new_n810), .A3(new_n853), .A4(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n869), .B1(G952), .B2(G953), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT49), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n793), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n872), .A2(new_n588), .A3(new_n671), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n793), .A2(new_n871), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n781), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n875), .A2(new_n287), .A3(new_n583), .A4(new_n660), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n870), .A2(new_n876), .ZN(G75));
  AOI21_X1  g691(.A(new_n866), .B1(new_n848), .B2(new_n854), .ZN(new_n878));
  OAI21_X1  g692(.A(KEYINPUT114), .B1(new_n878), .B2(new_n276), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT114), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT53), .B1(new_n850), .B2(new_n828), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n880), .B(G902), .C1(new_n881), .C2(new_n866), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n879), .A2(new_n882), .A3(new_n279), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n222), .A2(new_n264), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(new_n262), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n885), .B(KEYINPUT55), .Z(new_n886));
  INV_X1    g700(.A(KEYINPUT115), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT116), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n889), .B1(new_n887), .B2(KEYINPUT56), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n888), .B(new_n890), .C1(new_n887), .C2(KEYINPUT56), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n891), .B1(KEYINPUT116), .B2(new_n888), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n883), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n292), .A2(G952), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n878), .A2(new_n529), .A3(new_n276), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n886), .B1(new_n896), .B2(KEYINPUT56), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n893), .A2(new_n895), .A3(new_n897), .ZN(G51));
  OR2_X1    g712(.A1(new_n329), .A2(new_n344), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n346), .B(KEYINPUT117), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT57), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI211_X1 g716(.A(KEYINPUT54), .B(new_n866), .C1(new_n848), .C2(new_n854), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n858), .B1(new_n857), .B2(new_n867), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n902), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n900), .A2(new_n901), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n899), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n748), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n879), .A2(new_n882), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n894), .B1(new_n907), .B2(new_n909), .ZN(G54));
  AND2_X1   g724(.A1(KEYINPUT58), .A2(G475), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n879), .A2(new_n882), .A3(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n455), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n879), .A2(new_n882), .A3(new_n455), .A4(new_n911), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n914), .A2(new_n895), .A3(new_n915), .ZN(G60));
  XNOR2_X1  g730(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n397), .A2(new_n276), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n917), .B(new_n918), .Z(new_n919));
  XOR2_X1   g733(.A(new_n592), .B(KEYINPUT118), .Z(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n919), .B(new_n921), .C1(new_n903), .C2(new_n904), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n895), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n853), .A2(new_n868), .ZN(new_n924));
  INV_X1    g738(.A(new_n919), .ZN(new_n925));
  OAI211_X1 g739(.A(KEYINPUT120), .B(new_n920), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT120), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n925), .B1(new_n853), .B2(new_n868), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n927), .B1(new_n928), .B2(new_n921), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n923), .B1(new_n926), .B2(new_n929), .ZN(G63));
  NAND2_X1  g744(.A1(new_n618), .A2(new_n620), .ZN(new_n931));
  NAND2_X1  g745(.A1(G217), .A2(G902), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT60), .ZN(new_n933));
  OR3_X1    g747(.A1(new_n878), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  OAI22_X1  g748(.A1(new_n878), .A2(new_n933), .B1(new_n494), .B2(new_n495), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n934), .A2(new_n935), .A3(new_n895), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n934), .A2(new_n935), .A3(KEYINPUT61), .A4(new_n895), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(G66));
  OAI21_X1  g754(.A(G953), .B1(new_n466), .B2(new_n257), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n941), .B1(new_n847), .B2(G953), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n884), .B1(G898), .B2(new_n292), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(G69));
  NOR2_X1   g758(.A1(new_n536), .A2(new_n537), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n446), .A2(new_n447), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n945), .B(new_n946), .Z(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(G900), .A2(G953), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n823), .A2(new_n674), .ZN(new_n950));
  OAI21_X1  g764(.A(KEYINPUT124), .B1(new_n760), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n758), .A2(new_n759), .ZN(new_n952));
  INV_X1    g766(.A(new_n754), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT124), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n823), .A2(new_n674), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n951), .A2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n768), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n959), .B1(new_n719), .B2(new_n721), .ZN(new_n960));
  INV_X1    g774(.A(new_n811), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n716), .A2(new_n662), .A3(new_n753), .A4(new_n961), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n958), .A2(new_n727), .A3(new_n960), .A4(new_n962), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n948), .B(new_n949), .C1(new_n963), .C2(G953), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n668), .A2(new_n956), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT62), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n668), .A2(new_n956), .A3(KEYINPUT62), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n836), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n578), .A2(new_n726), .A3(new_n662), .A4(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT122), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n971), .A2(new_n972), .ZN(new_n974));
  NOR4_X1   g788(.A1(new_n959), .A2(new_n760), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(G953), .B1(new_n969), .B2(new_n975), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n947), .A2(KEYINPUT121), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n947), .A2(KEYINPUT121), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(KEYINPUT123), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT123), .ZN(new_n982));
  NOR4_X1   g796(.A1(new_n976), .A2(new_n982), .A3(new_n979), .A4(new_n977), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n964), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n292), .B1(G227), .B2(G900), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n985), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n987), .B(new_n964), .C1(new_n981), .C2(new_n983), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n986), .A2(new_n988), .ZN(G72));
  NAND2_X1  g803(.A1(G472), .A2(G902), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT63), .Z(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT125), .Z(new_n992));
  INV_X1    g806(.A(new_n847), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n992), .B1(new_n963), .B2(new_n993), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n994), .A2(new_n533), .A3(new_n539), .A4(new_n538), .ZN(new_n995));
  AND3_X1   g809(.A1(new_n995), .A2(KEYINPUT126), .A3(new_n895), .ZN(new_n996));
  AOI21_X1  g810(.A(KEYINPUT126), .B1(new_n995), .B2(new_n895), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n969), .A2(new_n975), .A3(new_n847), .ZN(new_n998));
  AND2_X1   g812(.A1(new_n998), .A2(new_n992), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n849), .A2(new_n852), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n563), .A2(new_n541), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(new_n991), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(KEYINPUT127), .ZN(new_n1003));
  OAI22_X1  g817(.A1(new_n999), .A2(new_n656), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  NOR3_X1   g818(.A1(new_n996), .A2(new_n997), .A3(new_n1004), .ZN(G57));
endmodule


