

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590;

  XNOR2_X1 U324 ( .A(n331), .B(n330), .ZN(n335) );
  XNOR2_X1 U325 ( .A(n359), .B(n358), .ZN(n473) );
  XNOR2_X1 U326 ( .A(n428), .B(KEYINPUT64), .ZN(n574) );
  XNOR2_X1 U327 ( .A(n344), .B(n343), .ZN(n562) );
  XNOR2_X1 U328 ( .A(G120GAT), .B(n357), .ZN(n292) );
  XOR2_X1 U329 ( .A(n389), .B(n388), .Z(n293) );
  XNOR2_X1 U330 ( .A(KEYINPUT47), .B(KEYINPUT107), .ZN(n382) );
  XNOR2_X1 U331 ( .A(n383), .B(n382), .ZN(n384) );
  INV_X1 U332 ( .A(KEYINPUT92), .ZN(n392) );
  XNOR2_X1 U333 ( .A(n402), .B(KEYINPUT54), .ZN(n403) );
  XNOR2_X1 U334 ( .A(n329), .B(n357), .ZN(n330) );
  XNOR2_X1 U335 ( .A(n393), .B(n392), .ZN(n394) );
  INV_X1 U336 ( .A(KEYINPUT37), .ZN(n469) );
  XNOR2_X1 U337 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U338 ( .A(n397), .B(n292), .ZN(n358) );
  XNOR2_X1 U339 ( .A(n470), .B(n469), .ZN(n471) );
  XOR2_X1 U340 ( .A(n562), .B(KEYINPUT36), .Z(n587) );
  XNOR2_X1 U341 ( .A(n472), .B(n471), .ZN(n519) );
  NOR2_X1 U342 ( .A1(n503), .A2(n450), .ZN(n570) );
  XOR2_X1 U343 ( .A(KEYINPUT41), .B(n579), .Z(n557) );
  INV_X1 U344 ( .A(G50GAT), .ZN(n476) );
  XOR2_X1 U345 ( .A(n311), .B(n310), .Z(n532) );
  XNOR2_X1 U346 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U347 ( .A(n476), .B(KEYINPUT100), .ZN(n477) );
  XNOR2_X1 U348 ( .A(n482), .B(n481), .ZN(G1351GAT) );
  XNOR2_X1 U349 ( .A(n478), .B(n477), .ZN(G1331GAT) );
  XNOR2_X1 U350 ( .A(G43GAT), .B(G190GAT), .ZN(n294) );
  XNOR2_X1 U351 ( .A(n294), .B(G134GAT), .ZN(n296) );
  XNOR2_X1 U352 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n295) );
  XNOR2_X1 U353 ( .A(n295), .B(KEYINPUT18), .ZN(n388) );
  XOR2_X1 U354 ( .A(n296), .B(n388), .Z(n303) );
  XOR2_X1 U355 ( .A(G120GAT), .B(KEYINPUT81), .Z(n298) );
  XNOR2_X1 U356 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n297) );
  XNOR2_X1 U357 ( .A(n298), .B(n297), .ZN(n413) );
  XOR2_X1 U358 ( .A(n413), .B(KEYINPUT20), .Z(n300) );
  NAND2_X1 U359 ( .A1(G227GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U360 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U361 ( .A(n301), .B(G99GAT), .ZN(n302) );
  XNOR2_X1 U362 ( .A(n303), .B(n302), .ZN(n311) );
  XOR2_X1 U363 ( .A(G176GAT), .B(G71GAT), .Z(n305) );
  XNOR2_X1 U364 ( .A(G169GAT), .B(G127GAT), .ZN(n304) );
  XNOR2_X1 U365 ( .A(n305), .B(n304), .ZN(n309) );
  XOR2_X1 U366 ( .A(KEYINPUT82), .B(KEYINPUT83), .Z(n307) );
  XNOR2_X1 U367 ( .A(G15GAT), .B(G183GAT), .ZN(n306) );
  XNOR2_X1 U368 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U369 ( .A(n309), .B(n308), .Z(n310) );
  INV_X1 U370 ( .A(n532), .ZN(n503) );
  XNOR2_X1 U371 ( .A(G1GAT), .B(G22GAT), .ZN(n312) );
  XNOR2_X1 U372 ( .A(n312), .B(G15GAT), .ZN(n360) );
  XNOR2_X1 U373 ( .A(G8GAT), .B(G183GAT), .ZN(n313) );
  XNOR2_X1 U374 ( .A(n313), .B(G211GAT), .ZN(n391) );
  XNOR2_X1 U375 ( .A(n360), .B(n391), .ZN(n325) );
  XOR2_X1 U376 ( .A(G127GAT), .B(G155GAT), .Z(n416) );
  XOR2_X1 U377 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n315) );
  XNOR2_X1 U378 ( .A(G64GAT), .B(KEYINPUT15), .ZN(n314) );
  XNOR2_X1 U379 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U380 ( .A(n416), .B(n316), .Z(n318) );
  NAND2_X1 U381 ( .A1(G231GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U382 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U383 ( .A(n319), .B(KEYINPUT80), .Z(n323) );
  XOR2_X1 U384 ( .A(G78GAT), .B(KEYINPUT13), .Z(n321) );
  XNOR2_X1 U385 ( .A(G71GAT), .B(G57GAT), .ZN(n320) );
  XNOR2_X1 U386 ( .A(n321), .B(n320), .ZN(n347) );
  XNOR2_X1 U387 ( .A(n347), .B(KEYINPUT79), .ZN(n322) );
  XNOR2_X1 U388 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U389 ( .A(n325), .B(n324), .Z(n582) );
  INV_X1 U390 ( .A(n582), .ZN(n483) );
  XOR2_X1 U391 ( .A(KEYINPUT76), .B(G92GAT), .Z(n327) );
  XNOR2_X1 U392 ( .A(G50GAT), .B(G162GAT), .ZN(n326) );
  XNOR2_X1 U393 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U394 ( .A(n328), .B(G106GAT), .Z(n331) );
  XOR2_X1 U395 ( .A(G190GAT), .B(G218GAT), .Z(n389) );
  XNOR2_X1 U396 ( .A(G36GAT), .B(n389), .ZN(n329) );
  XOR2_X1 U397 ( .A(G99GAT), .B(G85GAT), .Z(n357) );
  XOR2_X1 U398 ( .A(G29GAT), .B(G43GAT), .Z(n333) );
  XNOR2_X1 U399 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n332) );
  XNOR2_X1 U400 ( .A(n333), .B(n332), .ZN(n362) );
  XOR2_X1 U401 ( .A(G134GAT), .B(KEYINPUT77), .Z(n417) );
  XOR2_X1 U402 ( .A(n362), .B(n417), .Z(n334) );
  XNOR2_X1 U403 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U404 ( .A(KEYINPUT78), .B(KEYINPUT73), .Z(n337) );
  NAND2_X1 U405 ( .A1(G232GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U406 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U407 ( .A(n339), .B(n338), .ZN(n344) );
  XOR2_X1 U408 ( .A(KEYINPUT74), .B(KEYINPUT75), .Z(n341) );
  XNOR2_X1 U409 ( .A(KEYINPUT9), .B(KEYINPUT10), .ZN(n340) );
  XNOR2_X1 U410 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U411 ( .A(n342), .B(KEYINPUT11), .ZN(n343) );
  NOR2_X1 U412 ( .A1(n483), .A2(n587), .ZN(n345) );
  XNOR2_X1 U413 ( .A(KEYINPUT45), .B(n345), .ZN(n376) );
  XNOR2_X1 U414 ( .A(G148GAT), .B(G106GAT), .ZN(n346) );
  XNOR2_X1 U415 ( .A(n346), .B(KEYINPUT71), .ZN(n442) );
  XNOR2_X1 U416 ( .A(n347), .B(n442), .ZN(n352) );
  XOR2_X1 U417 ( .A(KEYINPUT70), .B(KEYINPUT33), .Z(n349) );
  NAND2_X1 U418 ( .A1(G230GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U419 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U420 ( .A(n350), .B(KEYINPUT31), .Z(n351) );
  XNOR2_X1 U421 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U422 ( .A(n353), .B(KEYINPUT32), .ZN(n359) );
  XOR2_X1 U423 ( .A(G204GAT), .B(KEYINPUT72), .Z(n355) );
  XNOR2_X1 U424 ( .A(G176GAT), .B(G92GAT), .ZN(n354) );
  XNOR2_X1 U425 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U426 ( .A(G64GAT), .B(n356), .Z(n397) );
  INV_X1 U427 ( .A(n473), .ZN(n579) );
  XOR2_X1 U428 ( .A(G169GAT), .B(G36GAT), .Z(n398) );
  XOR2_X1 U429 ( .A(G50GAT), .B(G141GAT), .Z(n441) );
  XNOR2_X1 U430 ( .A(n398), .B(n441), .ZN(n361) );
  XNOR2_X1 U431 ( .A(n361), .B(n360), .ZN(n366) );
  XOR2_X1 U432 ( .A(n362), .B(KEYINPUT66), .Z(n364) );
  NAND2_X1 U433 ( .A1(G229GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U434 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U435 ( .A(n366), .B(n365), .Z(n374) );
  XOR2_X1 U436 ( .A(G197GAT), .B(G8GAT), .Z(n368) );
  XNOR2_X1 U437 ( .A(G113GAT), .B(KEYINPUT67), .ZN(n367) );
  XNOR2_X1 U438 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U439 ( .A(KEYINPUT29), .B(KEYINPUT68), .Z(n370) );
  XNOR2_X1 U440 ( .A(KEYINPUT30), .B(KEYINPUT65), .ZN(n369) );
  XNOR2_X1 U441 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U442 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U443 ( .A(n374), .B(n373), .Z(n508) );
  XNOR2_X1 U444 ( .A(n508), .B(KEYINPUT69), .ZN(n566) );
  NOR2_X1 U445 ( .A1(n579), .A2(n566), .ZN(n375) );
  AND2_X1 U446 ( .A1(n376), .A2(n375), .ZN(n377) );
  XOR2_X1 U447 ( .A(n377), .B(KEYINPUT108), .Z(n385) );
  XOR2_X1 U448 ( .A(KEYINPUT106), .B(n483), .Z(n569) );
  INV_X1 U449 ( .A(n508), .ZN(n575) );
  NAND2_X1 U450 ( .A1(n575), .A2(n557), .ZN(n378) );
  XOR2_X1 U451 ( .A(KEYINPUT46), .B(n378), .Z(n379) );
  NOR2_X1 U452 ( .A1(n569), .A2(n379), .ZN(n381) );
  INV_X1 U453 ( .A(n562), .ZN(n380) );
  NAND2_X1 U454 ( .A1(n381), .A2(n380), .ZN(n383) );
  AND2_X1 U455 ( .A1(n385), .A2(n384), .ZN(n387) );
  XOR2_X1 U456 ( .A(KEYINPUT109), .B(KEYINPUT48), .Z(n386) );
  XNOR2_X1 U457 ( .A(n387), .B(n386), .ZN(n531) );
  NAND2_X1 U458 ( .A1(G226GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U459 ( .A(n293), .B(n390), .ZN(n395) );
  XNOR2_X1 U460 ( .A(n391), .B(KEYINPUT91), .ZN(n393) );
  XOR2_X1 U461 ( .A(G197GAT), .B(KEYINPUT21), .Z(n431) );
  XOR2_X1 U462 ( .A(n396), .B(n431), .Z(n400) );
  XNOR2_X1 U463 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U464 ( .A(n400), .B(n399), .Z(n455) );
  XOR2_X1 U465 ( .A(n455), .B(KEYINPUT120), .Z(n401) );
  NOR2_X1 U466 ( .A1(n531), .A2(n401), .ZN(n404) );
  XOR2_X1 U467 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n402) );
  XNOR2_X1 U468 ( .A(n404), .B(n403), .ZN(n427) );
  XOR2_X1 U469 ( .A(KEYINPUT88), .B(G148GAT), .Z(n406) );
  XNOR2_X1 U470 ( .A(G1GAT), .B(G57GAT), .ZN(n405) );
  XNOR2_X1 U471 ( .A(n406), .B(n405), .ZN(n426) );
  XOR2_X1 U472 ( .A(KEYINPUT89), .B(KEYINPUT4), .Z(n408) );
  XNOR2_X1 U473 ( .A(G29GAT), .B(G85GAT), .ZN(n407) );
  XNOR2_X1 U474 ( .A(n408), .B(n407), .ZN(n412) );
  XOR2_X1 U475 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n410) );
  XNOR2_X1 U476 ( .A(G141GAT), .B(KEYINPUT90), .ZN(n409) );
  XNOR2_X1 U477 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U478 ( .A(n412), .B(n411), .Z(n424) );
  XOR2_X1 U479 ( .A(n413), .B(KEYINPUT5), .Z(n415) );
  NAND2_X1 U480 ( .A1(G225GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U481 ( .A(n415), .B(n414), .ZN(n422) );
  XNOR2_X1 U482 ( .A(n417), .B(n416), .ZN(n420) );
  XOR2_X1 U483 ( .A(KEYINPUT3), .B(KEYINPUT86), .Z(n419) );
  XNOR2_X1 U484 ( .A(G162GAT), .B(KEYINPUT2), .ZN(n418) );
  XNOR2_X1 U485 ( .A(n419), .B(n418), .ZN(n436) );
  XNOR2_X1 U486 ( .A(n420), .B(n436), .ZN(n421) );
  XNOR2_X1 U487 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U488 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U489 ( .A(n426), .B(n425), .ZN(n520) );
  INV_X1 U490 ( .A(n520), .ZN(n497) );
  NAND2_X1 U491 ( .A1(n427), .A2(n497), .ZN(n428) );
  XOR2_X1 U492 ( .A(G204GAT), .B(G78GAT), .Z(n430) );
  XNOR2_X1 U493 ( .A(G155GAT), .B(G218GAT), .ZN(n429) );
  XNOR2_X1 U494 ( .A(n430), .B(n429), .ZN(n432) );
  XOR2_X1 U495 ( .A(n432), .B(n431), .Z(n434) );
  XNOR2_X1 U496 ( .A(G22GAT), .B(G211GAT), .ZN(n433) );
  XNOR2_X1 U497 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U498 ( .A(n435), .B(KEYINPUT23), .Z(n438) );
  XNOR2_X1 U499 ( .A(n436), .B(KEYINPUT87), .ZN(n437) );
  XNOR2_X1 U500 ( .A(n438), .B(n437), .ZN(n448) );
  XOR2_X1 U501 ( .A(KEYINPUT85), .B(KEYINPUT22), .Z(n440) );
  XNOR2_X1 U502 ( .A(KEYINPUT24), .B(KEYINPUT84), .ZN(n439) );
  XNOR2_X1 U503 ( .A(n440), .B(n439), .ZN(n446) );
  XOR2_X1 U504 ( .A(n442), .B(n441), .Z(n444) );
  NAND2_X1 U505 ( .A1(G228GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U506 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U507 ( .A(n446), .B(n445), .Z(n447) );
  XNOR2_X1 U508 ( .A(n448), .B(n447), .ZN(n463) );
  NOR2_X1 U509 ( .A1(n574), .A2(n463), .ZN(n449) );
  XNOR2_X1 U510 ( .A(n449), .B(KEYINPUT55), .ZN(n450) );
  XOR2_X1 U511 ( .A(KEYINPUT101), .B(n557), .Z(n537) );
  NAND2_X1 U512 ( .A1(n570), .A2(n537), .ZN(n454) );
  XOR2_X1 U513 ( .A(G176GAT), .B(KEYINPUT124), .Z(n452) );
  XNOR2_X1 U514 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n451) );
  XNOR2_X1 U515 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U516 ( .A(n454), .B(n453), .ZN(G1349GAT) );
  INV_X1 U517 ( .A(n455), .ZN(n501) );
  NOR2_X1 U518 ( .A1(n501), .A2(n503), .ZN(n456) );
  NOR2_X1 U519 ( .A1(n463), .A2(n456), .ZN(n457) );
  XOR2_X1 U520 ( .A(KEYINPUT25), .B(n457), .Z(n460) );
  NAND2_X1 U521 ( .A1(n463), .A2(n503), .ZN(n458) );
  XNOR2_X1 U522 ( .A(n458), .B(KEYINPUT26), .ZN(n573) );
  XOR2_X1 U523 ( .A(n455), .B(KEYINPUT27), .Z(n462) );
  NOR2_X1 U524 ( .A1(n573), .A2(n462), .ZN(n459) );
  NOR2_X1 U525 ( .A1(n460), .A2(n459), .ZN(n461) );
  NOR2_X1 U526 ( .A1(n520), .A2(n461), .ZN(n465) );
  NOR2_X1 U527 ( .A1(n497), .A2(n462), .ZN(n549) );
  XNOR2_X1 U528 ( .A(KEYINPUT28), .B(n463), .ZN(n526) );
  INV_X1 U529 ( .A(n526), .ZN(n475) );
  NAND2_X1 U530 ( .A1(n549), .A2(n475), .ZN(n534) );
  NOR2_X1 U531 ( .A1(n532), .A2(n534), .ZN(n464) );
  NOR2_X1 U532 ( .A1(n465), .A2(n464), .ZN(n466) );
  XNOR2_X1 U533 ( .A(KEYINPUT93), .B(n466), .ZN(n485) );
  INV_X1 U534 ( .A(n485), .ZN(n467) );
  NOR2_X1 U535 ( .A1(n467), .A2(n587), .ZN(n468) );
  NAND2_X1 U536 ( .A1(n468), .A2(n483), .ZN(n472) );
  XOR2_X1 U537 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n470) );
  NAND2_X1 U538 ( .A1(n566), .A2(n473), .ZN(n487) );
  NOR2_X1 U539 ( .A1(n519), .A2(n487), .ZN(n474) );
  XOR2_X1 U540 ( .A(KEYINPUT38), .B(n474), .Z(n504) );
  NOR2_X1 U541 ( .A1(n504), .A2(n475), .ZN(n478) );
  NAND2_X1 U542 ( .A1(n570), .A2(n562), .ZN(n482) );
  XOR2_X1 U543 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n480) );
  INV_X1 U544 ( .A(G190GAT), .ZN(n479) );
  XNOR2_X1 U545 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n490) );
  NOR2_X1 U546 ( .A1(n483), .A2(n562), .ZN(n484) );
  XNOR2_X1 U547 ( .A(n484), .B(KEYINPUT16), .ZN(n486) );
  NAND2_X1 U548 ( .A1(n486), .A2(n485), .ZN(n509) );
  NOR2_X1 U549 ( .A1(n487), .A2(n509), .ZN(n488) );
  XNOR2_X1 U550 ( .A(KEYINPUT94), .B(n488), .ZN(n495) );
  NAND2_X1 U551 ( .A1(n520), .A2(n495), .ZN(n489) );
  XNOR2_X1 U552 ( .A(n490), .B(n489), .ZN(G1324GAT) );
  XOR2_X1 U553 ( .A(G8GAT), .B(KEYINPUT95), .Z(n492) );
  NAND2_X1 U554 ( .A1(n495), .A2(n455), .ZN(n491) );
  XNOR2_X1 U555 ( .A(n492), .B(n491), .ZN(G1325GAT) );
  XOR2_X1 U556 ( .A(G15GAT), .B(KEYINPUT35), .Z(n494) );
  NAND2_X1 U557 ( .A1(n532), .A2(n495), .ZN(n493) );
  XNOR2_X1 U558 ( .A(n494), .B(n493), .ZN(G1326GAT) );
  NAND2_X1 U559 ( .A1(n495), .A2(n526), .ZN(n496) );
  XNOR2_X1 U560 ( .A(n496), .B(G22GAT), .ZN(G1327GAT) );
  XNOR2_X1 U561 ( .A(KEYINPUT96), .B(KEYINPUT39), .ZN(n499) );
  NOR2_X1 U562 ( .A1(n497), .A2(n504), .ZN(n498) );
  XNOR2_X1 U563 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U564 ( .A(G29GAT), .B(n500), .ZN(G1328GAT) );
  NOR2_X1 U565 ( .A1(n501), .A2(n504), .ZN(n502) );
  XOR2_X1 U566 ( .A(G36GAT), .B(n502), .Z(G1329GAT) );
  NOR2_X1 U567 ( .A1(n504), .A2(n503), .ZN(n506) );
  XNOR2_X1 U568 ( .A(KEYINPUT40), .B(KEYINPUT99), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U570 ( .A(G43GAT), .B(n507), .ZN(G1330GAT) );
  XNOR2_X1 U571 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n511) );
  NAND2_X1 U572 ( .A1(n508), .A2(n537), .ZN(n518) );
  NOR2_X1 U573 ( .A1(n509), .A2(n518), .ZN(n515) );
  NAND2_X1 U574 ( .A1(n515), .A2(n520), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n511), .B(n510), .ZN(G1332GAT) );
  NAND2_X1 U576 ( .A1(n455), .A2(n515), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n512), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U578 ( .A1(n515), .A2(n532), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n513), .B(KEYINPUT102), .ZN(n514) );
  XNOR2_X1 U580 ( .A(G71GAT), .B(n514), .ZN(G1334GAT) );
  XOR2_X1 U581 ( .A(G78GAT), .B(KEYINPUT43), .Z(n517) );
  NAND2_X1 U582 ( .A1(n515), .A2(n526), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  XOR2_X1 U584 ( .A(G85GAT), .B(KEYINPUT103), .Z(n522) );
  NOR2_X1 U585 ( .A1(n519), .A2(n518), .ZN(n527) );
  NAND2_X1 U586 ( .A1(n527), .A2(n520), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n522), .B(n521), .ZN(G1336GAT) );
  NAND2_X1 U588 ( .A1(n455), .A2(n527), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n523), .B(KEYINPUT104), .ZN(n524) );
  XNOR2_X1 U590 ( .A(G92GAT), .B(n524), .ZN(G1337GAT) );
  NAND2_X1 U591 ( .A1(n527), .A2(n532), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n525), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT105), .B(KEYINPUT44), .Z(n529) );
  NAND2_X1 U594 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U595 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(n530), .ZN(G1339GAT) );
  XNOR2_X1 U597 ( .A(G113GAT), .B(KEYINPUT110), .ZN(n536) );
  INV_X1 U598 ( .A(n531), .ZN(n550) );
  NAND2_X1 U599 ( .A1(n532), .A2(n550), .ZN(n533) );
  NOR2_X1 U600 ( .A1(n534), .A2(n533), .ZN(n546) );
  NAND2_X1 U601 ( .A1(n566), .A2(n546), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n536), .B(n535), .ZN(G1340GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT49), .B(KEYINPUT112), .Z(n539) );
  NAND2_X1 U604 ( .A1(n546), .A2(n537), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(n541) );
  XOR2_X1 U606 ( .A(G120GAT), .B(KEYINPUT111), .Z(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  XNOR2_X1 U608 ( .A(G127GAT), .B(KEYINPUT113), .ZN(n545) );
  XOR2_X1 U609 ( .A(KEYINPUT114), .B(KEYINPUT50), .Z(n543) );
  NAND2_X1 U610 ( .A1(n546), .A2(n569), .ZN(n542) );
  XNOR2_X1 U611 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(G1342GAT) );
  XOR2_X1 U613 ( .A(G134GAT), .B(KEYINPUT51), .Z(n548) );
  NAND2_X1 U614 ( .A1(n546), .A2(n562), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(G1343GAT) );
  XOR2_X1 U616 ( .A(G141GAT), .B(KEYINPUT115), .Z(n553) );
  NAND2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X1 U618 ( .A1(n573), .A2(n551), .ZN(n563) );
  NAND2_X1 U619 ( .A1(n563), .A2(n575), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT117), .Z(n555) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U624 ( .A(KEYINPUT52), .B(n556), .Z(n559) );
  NAND2_X1 U625 ( .A1(n563), .A2(n557), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1345GAT) );
  NAND2_X1 U627 ( .A1(n582), .A2(n563), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n560), .B(KEYINPUT118), .ZN(n561) );
  XNOR2_X1 U629 ( .A(G155GAT), .B(n561), .ZN(G1346GAT) );
  XOR2_X1 U630 ( .A(G162GAT), .B(KEYINPUT119), .Z(n565) );
  NAND2_X1 U631 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(G1347GAT) );
  XOR2_X1 U633 ( .A(G169GAT), .B(KEYINPUT123), .Z(n568) );
  NAND2_X1 U634 ( .A1(n570), .A2(n566), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(G1348GAT) );
  XOR2_X1 U636 ( .A(G183GAT), .B(KEYINPUT125), .Z(n572) );
  NAND2_X1 U637 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(G1350GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n577) );
  NOR2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n585) );
  NAND2_X1 U641 ( .A1(n585), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT61), .Z(n581) );
  NAND2_X1 U645 ( .A1(n585), .A2(n579), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1353GAT) );
  XOR2_X1 U647 ( .A(G211GAT), .B(KEYINPUT127), .Z(n584) );
  NAND2_X1 U648 ( .A1(n585), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1354GAT) );
  INV_X1 U650 ( .A(KEYINPUT62), .ZN(n589) );
  INV_X1 U651 ( .A(n585), .ZN(n586) );
  NOR2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

