//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 1 0 0 0 0 0 0 0 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n808, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1024, new_n1025;
  INV_X1    g000(.A(G197gat), .ZN(new_n202));
  INV_X1    g001(.A(G204gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G197gat), .A2(G204gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT22), .ZN(new_n206));
  NAND2_X1  g005(.A1(G211gat), .A2(G218gat), .ZN(new_n207));
  AOI22_X1  g006(.A1(new_n204), .A2(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G211gat), .ZN(new_n209));
  INV_X1    g008(.A(G218gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT75), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n211), .A2(new_n212), .A3(new_n207), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n208), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n208), .A2(new_n213), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G183gat), .ZN(new_n217));
  INV_X1    g016(.A(G190gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n220));
  AND2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n223));
  AND2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n222), .A2(new_n223), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n221), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n229), .A2(G169gat), .A3(G176gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT23), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(G169gat), .B2(G176gat), .ZN(new_n233));
  AND2_X1   g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT65), .B(G176gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n232), .A2(G169gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n226), .A2(new_n234), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT25), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(G176gat), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n239), .B1(new_n236), .B2(new_n241), .ZN(new_n242));
  AND3_X1   g041(.A1(new_n242), .A2(new_n231), .A3(new_n233), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n217), .A2(new_n218), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n221), .B1(KEYINPUT24), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n240), .A2(new_n246), .ZN(new_n247));
  AND2_X1   g046(.A1(G226gat), .A2(G233gat), .ZN(new_n248));
  NOR3_X1   g047(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT68), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n231), .A2(KEYINPUT67), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT67), .B1(new_n231), .B2(new_n251), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n250), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT27), .B(G183gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(new_n218), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT28), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n255), .A2(KEYINPUT28), .A3(new_n218), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n244), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n254), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n247), .A2(new_n248), .A3(new_n261), .ZN(new_n262));
  AOI22_X1  g061(.A1(new_n238), .A2(new_n239), .B1(new_n245), .B2(new_n243), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n249), .B(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n229), .B1(G169gat), .B2(G176gat), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n251), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT67), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n231), .A2(KEYINPUT67), .A3(new_n251), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n266), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT28), .B1(new_n255), .B2(new_n218), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n217), .A2(KEYINPUT27), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT27), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G183gat), .ZN(new_n277));
  AND4_X1   g076(.A1(KEYINPUT28), .A2(new_n275), .A3(new_n277), .A4(new_n218), .ZN(new_n278));
  OAI22_X1  g077(.A1(new_n274), .A2(new_n278), .B1(new_n217), .B2(new_n218), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n264), .B1(new_n273), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n254), .A2(new_n260), .A3(KEYINPUT69), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n263), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n248), .A2(KEYINPUT29), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n216), .B(new_n262), .C1(new_n282), .C2(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n284), .B1(new_n247), .B2(new_n261), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n286), .B1(new_n248), .B2(new_n282), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n285), .B1(new_n287), .B2(new_n216), .ZN(new_n288));
  XNOR2_X1  g087(.A(G8gat), .B(G36gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(G64gat), .B(G92gat), .ZN(new_n290));
  XOR2_X1   g089(.A(new_n289), .B(new_n290), .Z(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT30), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n285), .B(new_n291), .C1(new_n287), .C2(new_n216), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n294), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  XOR2_X1   g098(.A(G141gat), .B(G148gat), .Z(new_n300));
  INV_X1    g099(.A(G155gat), .ZN(new_n301));
  INV_X1    g100(.A(G162gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(G155gat), .A2(G162gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(KEYINPUT2), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n300), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G141gat), .B(G148gat), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n304), .B(new_n303), .C1(new_n308), .C2(KEYINPUT2), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G127gat), .B(G134gat), .ZN(new_n311));
  INV_X1    g110(.A(G113gat), .ZN(new_n312));
  INV_X1    g111(.A(G120gat), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT1), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  OR2_X1    g114(.A1(KEYINPUT70), .A2(G113gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(KEYINPUT70), .A2(G113gat), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n313), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n312), .A2(new_n313), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT1), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n320), .B1(G113gat), .B2(G120gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  OAI22_X1  g121(.A1(new_n315), .A2(new_n318), .B1(new_n322), .B2(new_n311), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n310), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT4), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT78), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  XOR2_X1   g125(.A(KEYINPUT77), .B(KEYINPUT4), .Z(new_n327));
  NAND2_X1  g126(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n316), .A2(new_n317), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(G120gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n330), .A2(new_n314), .A3(new_n311), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n314), .B1(new_n312), .B2(new_n313), .ZN(new_n332));
  XOR2_X1   g131(.A(G127gat), .B(G134gat), .Z(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n331), .A2(new_n334), .A3(new_n309), .A4(new_n307), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT78), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n335), .A2(new_n336), .A3(KEYINPUT4), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n326), .A2(new_n328), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT5), .ZN(new_n339));
  NAND2_X1  g138(.A1(G225gat), .A2(G233gat), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT3), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n307), .A2(new_n309), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(new_n323), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n341), .B1(new_n307), .B2(new_n309), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n339), .B(new_n340), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n310), .A2(KEYINPUT3), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n347), .A2(new_n323), .A3(new_n342), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n335), .A2(new_n327), .ZN(new_n349));
  INV_X1    g148(.A(new_n323), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n307), .A2(new_n309), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n350), .A2(new_n351), .A3(KEYINPUT4), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n348), .A2(new_n349), .A3(new_n352), .A4(new_n340), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n310), .A2(new_n323), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(new_n335), .ZN(new_n355));
  INV_X1    g154(.A(new_n340), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n339), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI22_X1  g156(.A1(new_n338), .A2(new_n346), .B1(new_n353), .B2(new_n357), .ZN(new_n358));
  XOR2_X1   g157(.A(G1gat), .B(G29gat), .Z(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(KEYINPUT0), .ZN(new_n360));
  XNOR2_X1  g159(.A(G57gat), .B(G85gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT6), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n338), .A2(new_n346), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n353), .A2(new_n357), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n365), .A2(new_n366), .A3(new_n362), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT79), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT6), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n365), .A2(new_n366), .A3(KEYINPUT79), .A4(new_n362), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT85), .B1(new_n358), .B2(new_n362), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n365), .A2(new_n366), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT85), .ZN(new_n375));
  INV_X1    g174(.A(new_n362), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n364), .B1(new_n372), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n299), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT88), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT88), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n299), .A2(new_n382), .A3(new_n379), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NOR3_X1   g183(.A1(new_n273), .A2(new_n264), .A3(new_n279), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT69), .B1(new_n254), .B2(new_n260), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n247), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n350), .ZN(new_n388));
  INV_X1    g187(.A(G227gat), .ZN(new_n389));
  INV_X1    g188(.A(G233gat), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n323), .B(new_n247), .C1(new_n385), .C2(new_n386), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n388), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT32), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT33), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  XOR2_X1   g195(.A(G15gat), .B(G43gat), .Z(new_n397));
  XNOR2_X1  g196(.A(G71gat), .B(G99gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n397), .B(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n394), .A2(new_n396), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT34), .ZN(new_n401));
  INV_X1    g200(.A(new_n391), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n282), .A2(new_n323), .ZN(new_n403));
  AOI211_X1 g202(.A(new_n350), .B(new_n263), .C1(new_n280), .C2(new_n281), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n401), .B(new_n402), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n391), .B1(new_n388), .B2(new_n392), .ZN(new_n406));
  XOR2_X1   g205(.A(KEYINPUT71), .B(KEYINPUT34), .Z(new_n407));
  OAI21_X1  g206(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT72), .ZN(new_n409));
  INV_X1    g208(.A(new_n399), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n393), .B(KEYINPUT32), .C1(new_n395), .C2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n412));
  INV_X1    g211(.A(new_n407), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT72), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  AND4_X1   g214(.A1(new_n400), .A2(new_n409), .A3(new_n411), .A4(new_n415), .ZN(new_n416));
  AOI22_X1  g215(.A1(new_n409), .A2(new_n415), .B1(new_n400), .B2(new_n411), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(G78gat), .B(G106gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(KEYINPUT31), .B(G50gat), .ZN(new_n420));
  XOR2_X1   g219(.A(new_n419), .B(new_n420), .Z(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(G228gat), .A2(G233gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n423), .B(KEYINPUT81), .ZN(new_n424));
  INV_X1    g223(.A(new_n208), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n211), .A2(new_n207), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT29), .ZN(new_n428));
  INV_X1    g227(.A(new_n426), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n208), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n427), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n351), .B1(new_n431), .B2(new_n341), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n214), .A2(new_n215), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n433), .B1(new_n428), .B2(new_n342), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n424), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n342), .A2(new_n428), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n423), .B1(new_n436), .B2(new_n216), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT29), .B1(new_n214), .B2(new_n215), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n310), .B1(new_n438), .B2(KEYINPUT3), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n435), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(G22gat), .ZN(new_n442));
  INV_X1    g241(.A(G22gat), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n435), .A2(new_n440), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n422), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n443), .B1(new_n435), .B2(new_n440), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT82), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n444), .B(new_n422), .C1(new_n446), .C2(KEYINPUT82), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT83), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT82), .ZN(new_n451));
  INV_X1    g250(.A(new_n430), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n428), .B1(new_n429), .B2(new_n208), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n341), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n310), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n436), .A2(new_n216), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AOI22_X1  g256(.A1(new_n457), .A2(new_n424), .B1(new_n437), .B2(new_n439), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n451), .B1(new_n458), .B2(new_n443), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n421), .B1(new_n458), .B2(new_n443), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT83), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n447), .A2(new_n459), .A3(new_n460), .A4(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n445), .B1(new_n450), .B2(new_n462), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n463), .A2(KEYINPUT35), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n384), .A2(new_n418), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT73), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n400), .A2(new_n411), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n414), .B1(new_n408), .B2(KEYINPUT72), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n409), .A2(new_n415), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n400), .A2(new_n411), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(KEYINPUT73), .A3(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n445), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT82), .B1(new_n441), .B2(G22gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n444), .A2(new_n422), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n461), .B1(new_n476), .B2(new_n447), .ZN(new_n477));
  AND4_X1   g276(.A1(new_n461), .A2(new_n447), .A3(new_n459), .A4(new_n460), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n473), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n467), .A2(new_n468), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n469), .A2(new_n472), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT80), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n372), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n363), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n369), .A2(KEYINPUT80), .A3(new_n370), .A4(new_n371), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(new_n364), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n296), .A2(KEYINPUT76), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT76), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n293), .B(new_n489), .C1(new_n294), .C2(new_n295), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n490), .A2(new_n297), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n487), .A2(new_n488), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT35), .B1(new_n481), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n465), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n488), .A2(new_n490), .A3(new_n297), .ZN(new_n495));
  INV_X1    g294(.A(new_n364), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n363), .B1(new_n372), .B2(new_n482), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n496), .B1(new_n497), .B2(new_n485), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT84), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n479), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n463), .A2(KEYINPUT84), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n364), .B(new_n295), .C1(new_n372), .C2(new_n378), .ZN(new_n504));
  XNOR2_X1  g303(.A(KEYINPUT87), .B(KEYINPUT38), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT37), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n262), .B1(new_n282), .B2(new_n284), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(new_n433), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n508), .A2(KEYINPUT86), .B1(new_n216), .B2(new_n287), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT86), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n507), .A2(new_n510), .A3(new_n433), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n506), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n292), .B1(new_n288), .B2(KEYINPUT37), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n505), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n505), .B1(new_n288), .B2(KEYINPUT37), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n515), .B(new_n292), .C1(KEYINPUT37), .C2(new_n288), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n504), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n378), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n340), .B1(new_n338), .B2(new_n348), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT39), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(new_n362), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT39), .B1(new_n355), .B2(new_n356), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  NOR3_X1   g323(.A1(new_n522), .A2(KEYINPUT40), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT40), .ZN(new_n526));
  INV_X1    g325(.A(new_n524), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n376), .B1(new_n519), .B2(new_n520), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n518), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n479), .B1(new_n299), .B2(new_n530), .ZN(new_n531));
  OAI22_X1  g330(.A1(new_n499), .A2(new_n503), .B1(new_n517), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT36), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n533), .B1(new_n467), .B2(new_n468), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n469), .A2(new_n534), .A3(new_n472), .ZN(new_n535));
  XOR2_X1   g334(.A(KEYINPUT74), .B(KEYINPUT36), .Z(new_n536));
  OAI21_X1  g335(.A(new_n536), .B1(new_n416), .B2(new_n417), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n494), .B1(new_n532), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G113gat), .B(G141gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(G197gat), .ZN(new_n542));
  XOR2_X1   g341(.A(KEYINPUT11), .B(G169gat), .Z(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(KEYINPUT12), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  XOR2_X1   g345(.A(G43gat), .B(G50gat), .Z(new_n547));
  INV_X1    g346(.A(KEYINPUT89), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G43gat), .B(G50gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT89), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n549), .A2(KEYINPUT15), .A3(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(G29gat), .A2(G36gat), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT14), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  OR2_X1    g354(.A1(new_n550), .A2(KEYINPUT15), .ZN(new_n556));
  NAND2_X1  g355(.A1(G29gat), .A2(G36gat), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n557), .B(KEYINPUT90), .Z(new_n558));
  NAND4_X1  g357(.A1(new_n552), .A2(new_n555), .A3(new_n556), .A4(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n555), .A2(new_n557), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n560), .A2(KEYINPUT15), .A3(new_n549), .A4(new_n551), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT17), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G15gat), .B(G22gat), .ZN(new_n565));
  OR2_X1    g364(.A1(new_n565), .A2(G1gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT91), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT16), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n565), .B1(new_n568), .B2(G1gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n567), .A2(new_n570), .A3(G8gat), .ZN(new_n571));
  INV_X1    g370(.A(G8gat), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n566), .B(new_n569), .C1(KEYINPUT91), .C2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n559), .A2(KEYINPUT17), .A3(new_n561), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n564), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G229gat), .A2(G233gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n574), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT18), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n562), .B(new_n574), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n578), .B(KEYINPUT13), .Z(new_n583));
  AOI22_X1  g382(.A1(new_n580), .A2(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n577), .A2(KEYINPUT18), .A3(new_n578), .A4(new_n579), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT92), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n585), .A2(new_n586), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n546), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n589), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n591), .A2(new_n545), .A3(new_n584), .A4(new_n587), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n540), .A2(new_n593), .ZN(new_n594));
  AND2_X1   g393(.A1(G232gat), .A2(G233gat), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n595), .A2(KEYINPUT41), .ZN(new_n596));
  XNOR2_X1  g395(.A(G134gat), .B(G162gat), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n596), .B(new_n597), .Z(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT97), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT93), .ZN(new_n601));
  AND2_X1   g400(.A1(new_n564), .A2(new_n576), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT8), .ZN(new_n603));
  NAND2_X1  g402(.A1(G99gat), .A2(G106gat), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n603), .B1(new_n604), .B2(KEYINPUT95), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT95), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n606), .A2(G99gat), .A3(G106gat), .ZN(new_n607));
  INV_X1    g406(.A(G85gat), .ZN(new_n608));
  INV_X1    g407(.A(G92gat), .ZN(new_n609));
  AOI22_X1  g408(.A1(new_n605), .A2(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT7), .ZN(new_n611));
  OAI211_X1 g410(.A(KEYINPUT94), .B(new_n611), .C1(new_n608), .C2(new_n609), .ZN(new_n612));
  OAI21_X1  g411(.A(KEYINPUT94), .B1(new_n608), .B2(new_n609), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT94), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n614), .A2(G85gat), .A3(G92gat), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n613), .A2(new_n615), .A3(KEYINPUT7), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n610), .A2(new_n612), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G99gat), .B(G106gat), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n610), .A2(new_n618), .A3(new_n612), .A4(new_n616), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT96), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n620), .A2(KEYINPUT96), .A3(new_n621), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI22_X1  g425(.A1(new_n602), .A2(new_n626), .B1(KEYINPUT41), .B2(new_n595), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n624), .A2(new_n562), .A3(new_n625), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n627), .A2(new_n218), .A3(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n626), .A2(new_n564), .A3(new_n576), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n595), .A2(KEYINPUT41), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n630), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(G190gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n601), .B1(new_n634), .B2(new_n210), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n629), .A2(new_n633), .A3(G218gat), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n600), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n632), .A2(G190gat), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n632), .A2(G190gat), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n210), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AND4_X1   g439(.A1(KEYINPUT93), .A2(new_n640), .A3(new_n600), .A4(new_n636), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n599), .B1(new_n637), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n640), .A2(KEYINPUT93), .A3(new_n636), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(KEYINPUT97), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n635), .A2(new_n600), .A3(new_n636), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n644), .A2(new_n645), .A3(new_n598), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(G64gat), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n648), .A2(G57gat), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n648), .A2(G57gat), .ZN(new_n650));
  INV_X1    g449(.A(G71gat), .ZN(new_n651));
  INV_X1    g450(.A(G78gat), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  OAI22_X1  g452(.A1(new_n649), .A2(new_n650), .B1(new_n653), .B2(KEYINPUT9), .ZN(new_n654));
  XOR2_X1   g453(.A(G71gat), .B(G78gat), .Z(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT21), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(G231gat), .A2(G233gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(G127gat), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n575), .B1(new_n657), .B2(new_n656), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(new_n301), .ZN(new_n665));
  XOR2_X1   g464(.A(G183gat), .B(G211gat), .Z(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n663), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n663), .A2(new_n668), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n647), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(G230gat), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n674), .A2(new_n390), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT10), .ZN(new_n676));
  AND3_X1   g475(.A1(new_n656), .A2(new_n620), .A3(new_n621), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n656), .B1(new_n621), .B2(new_n620), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n656), .A2(new_n676), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n624), .A2(new_n625), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n675), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  NOR4_X1   g481(.A1(new_n677), .A2(new_n678), .A3(new_n674), .A4(new_n390), .ZN(new_n683));
  XNOR2_X1  g482(.A(G120gat), .B(G148gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(G176gat), .B(G204gat), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n684), .B(new_n685), .Z(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  OR3_X1    g486(.A1(new_n682), .A2(new_n683), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n687), .B1(new_n682), .B2(new_n683), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n594), .A2(new_n673), .A3(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n487), .ZN(new_n693));
  XOR2_X1   g492(.A(KEYINPUT98), .B(G1gat), .Z(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1324gat));
  XNOR2_X1  g494(.A(KEYINPUT16), .B(G8gat), .ZN(new_n696));
  NOR2_X1   g495(.A1(KEYINPUT100), .A2(KEYINPUT42), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n692), .A2(new_n299), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT99), .ZN(new_n702));
  OAI22_X1  g501(.A1(new_n699), .A2(new_n702), .B1(new_n700), .B2(G8gat), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n692), .A2(KEYINPUT99), .A3(new_n299), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n701), .B1(new_n703), .B2(new_n704), .ZN(G1325gat));
  AND3_X1   g504(.A1(new_n535), .A2(new_n537), .A3(KEYINPUT101), .ZN(new_n706));
  AOI21_X1  g505(.A(KEYINPUT101), .B1(new_n535), .B2(new_n537), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(G15gat), .B1(new_n692), .B2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n418), .ZN(new_n710));
  OR2_X1    g509(.A1(new_n710), .A2(G15gat), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n709), .B1(new_n692), .B2(new_n711), .ZN(G1326gat));
  NOR2_X1   g511(.A1(new_n692), .A2(new_n503), .ZN(new_n713));
  XOR2_X1   g512(.A(KEYINPUT43), .B(G22gat), .Z(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(G1327gat));
  NOR2_X1   g514(.A1(new_n671), .A2(new_n690), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n647), .A2(new_n716), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n717), .B(KEYINPUT102), .Z(new_n718));
  NAND2_X1  g517(.A1(new_n594), .A2(new_n718), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n719), .A2(G29gat), .A3(new_n487), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT45), .Z(new_n721));
  NOR3_X1   g520(.A1(new_n706), .A2(new_n707), .A3(new_n532), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n416), .A2(new_n463), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n499), .A2(new_n723), .A3(new_n469), .A4(new_n472), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n418), .A2(new_n464), .ZN(new_n725));
  AOI22_X1  g524(.A1(new_n724), .A2(KEYINPUT35), .B1(new_n725), .B2(new_n384), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n647), .B1(new_n722), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n637), .A2(new_n641), .A3(new_n599), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n598), .B1(new_n644), .B2(new_n645), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n731), .A2(new_n728), .ZN(new_n732));
  AOI22_X1  g531(.A1(new_n727), .A2(new_n728), .B1(new_n540), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g532(.A(KEYINPUT103), .B1(new_n590), .B2(new_n592), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n590), .A2(KEYINPUT103), .A3(new_n592), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n733), .A2(new_n716), .A3(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(G29gat), .B1(new_n739), .B2(new_n487), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n721), .A2(new_n740), .ZN(G1328gat));
  NOR3_X1   g540(.A1(new_n719), .A2(G36gat), .A3(new_n299), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT46), .ZN(new_n743));
  OAI21_X1  g542(.A(G36gat), .B1(new_n739), .B2(new_n299), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(G1329gat));
  OAI21_X1  g544(.A(G43gat), .B1(new_n739), .B2(new_n708), .ZN(new_n746));
  OR2_X1    g545(.A1(new_n710), .A2(G43gat), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n746), .B1(new_n719), .B2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT47), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1330gat));
  NOR2_X1   g549(.A1(new_n503), .A2(G50gat), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT105), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n752), .B1(new_n719), .B2(KEYINPUT104), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n753), .B1(KEYINPUT104), .B2(new_n719), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT48), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(G50gat), .B1(new_n739), .B2(new_n479), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OR2_X1    g557(.A1(new_n739), .A2(new_n503), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n754), .B1(G50gat), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n758), .B1(KEYINPUT48), .B2(new_n760), .ZN(G1331gat));
  INV_X1    g560(.A(KEYINPUT101), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n538), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n517), .ZN(new_n764));
  INV_X1    g563(.A(new_n531), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n450), .A2(new_n462), .ZN(new_n766));
  AOI21_X1  g565(.A(KEYINPUT84), .B1(new_n766), .B2(new_n473), .ZN(new_n767));
  AOI211_X1 g566(.A(new_n500), .B(new_n445), .C1(new_n450), .C2(new_n462), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI22_X1  g568(.A1(new_n764), .A2(new_n765), .B1(new_n492), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n535), .A2(new_n537), .A3(KEYINPUT101), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n763), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n494), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n642), .A2(new_n737), .A3(new_n671), .A4(new_n646), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n773), .A2(new_n690), .A3(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT106), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n498), .ZN(new_n779));
  XNOR2_X1  g578(.A(KEYINPUT107), .B(G57gat), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n779), .B(new_n780), .ZN(G1332gat));
  INV_X1    g580(.A(new_n299), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT49), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n782), .B1(new_n783), .B2(new_n648), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT108), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n778), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n786), .A2(KEYINPUT109), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(KEYINPUT109), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n788), .A2(new_n783), .A3(new_n648), .A4(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n789), .ZN(new_n791));
  OAI22_X1  g590(.A1(new_n791), .A2(new_n787), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n792), .ZN(G1333gat));
  OR2_X1    g592(.A1(new_n776), .A2(KEYINPUT106), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n776), .A2(KEYINPUT106), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XOR2_X1   g595(.A(new_n418), .B(KEYINPUT111), .Z(new_n797));
  OAI21_X1  g596(.A(new_n651), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT110), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n708), .A2(new_n651), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n799), .B1(new_n778), .B2(new_n800), .ZN(new_n801));
  AND4_X1   g600(.A1(new_n799), .A2(new_n794), .A3(new_n795), .A4(new_n800), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n798), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(KEYINPUT50), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n805), .B(new_n798), .C1(new_n801), .C2(new_n802), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(G1334gat));
  NAND2_X1  g606(.A1(new_n778), .A2(new_n769), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g608(.A1(new_n540), .A2(new_n732), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n738), .A2(new_n671), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n690), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n731), .B1(new_n772), .B2(new_n494), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n810), .B(new_n813), .C1(new_n814), .C2(KEYINPUT44), .ZN(new_n815));
  OAI21_X1  g614(.A(G85gat), .B1(new_n815), .B2(new_n487), .ZN(new_n816));
  NOR2_X1   g615(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n814), .A2(new_n811), .A3(new_n818), .ZN(new_n819));
  XOR2_X1   g618(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n820));
  AOI21_X1  g619(.A(new_n820), .B1(new_n814), .B2(new_n811), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n498), .A2(new_n608), .A3(new_n690), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n816), .B1(new_n822), .B2(new_n823), .ZN(G1336gat));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n299), .A2(G92gat), .A3(new_n691), .ZN(new_n827));
  NOR2_X1   g626(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  AND4_X1   g628(.A1(new_n647), .A2(new_n773), .A3(new_n811), .A4(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n829), .B1(new_n814), .B2(new_n811), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n827), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT114), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n727), .A2(new_n728), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n834), .A2(new_n782), .A3(new_n810), .A4(new_n813), .ZN(new_n835));
  AOI22_X1  g634(.A1(new_n832), .A2(new_n833), .B1(new_n835), .B2(G92gat), .ZN(new_n836));
  INV_X1    g635(.A(new_n827), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n773), .A2(new_n647), .A3(new_n811), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n828), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n814), .A2(new_n811), .A3(new_n829), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n837), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(KEYINPUT114), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n826), .B1(new_n836), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n827), .B1(new_n819), .B2(new_n821), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n826), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n733), .A2(new_n846), .A3(new_n782), .A4(new_n813), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n609), .B1(new_n835), .B2(KEYINPUT115), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n845), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n825), .B1(new_n843), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(G92gat), .B1(new_n815), .B2(new_n299), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n851), .B1(new_n841), .B2(KEYINPUT114), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n832), .A2(new_n833), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT52), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(KEYINPUT115), .B1(new_n815), .B2(new_n299), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n847), .A3(G92gat), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n856), .A2(new_n826), .A3(new_n844), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n854), .A2(KEYINPUT116), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n850), .A2(new_n858), .ZN(G1337gat));
  OAI21_X1  g658(.A(G99gat), .B1(new_n815), .B2(new_n708), .ZN(new_n860));
  OR3_X1    g659(.A1(new_n710), .A2(G99gat), .A3(new_n691), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n860), .B1(new_n822), .B2(new_n861), .ZN(G1338gat));
  OAI21_X1  g661(.A(G106gat), .B1(new_n815), .B2(new_n479), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n479), .A2(G106gat), .A3(new_n691), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n863), .B(new_n864), .C1(new_n822), .C2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n866), .B1(new_n839), .B2(new_n840), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n733), .A2(new_n769), .A3(new_n813), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n868), .B1(G106gat), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n867), .B1(new_n870), .B2(new_n864), .ZN(G1339gat));
  AND3_X1   g670(.A1(new_n590), .A2(KEYINPUT103), .A3(new_n592), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT55), .ZN(new_n873));
  INV_X1    g672(.A(new_n682), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n679), .A2(new_n675), .A3(new_n681), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n874), .A2(KEYINPUT54), .A3(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n686), .B1(new_n682), .B2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n873), .B1(new_n876), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n874), .A2(KEYINPUT54), .A3(new_n875), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(KEYINPUT55), .A3(new_n878), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n880), .A2(new_n688), .A3(new_n882), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n872), .A2(new_n734), .A3(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n582), .A2(new_n583), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n578), .B1(new_n577), .B2(new_n579), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n544), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n592), .A2(new_n690), .A3(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n646), .B(new_n642), .C1(new_n884), .C2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n592), .A2(new_n887), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n883), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n892), .B1(new_n729), .B2(new_n730), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n671), .B1(new_n890), .B2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n774), .A2(new_n690), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n769), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n487), .A2(new_n782), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n898), .A2(new_n418), .A3(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n593), .ZN(new_n901));
  OAI21_X1  g700(.A(G113gat), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(new_n899), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n903), .B1(new_n895), .B2(new_n897), .ZN(new_n904));
  INV_X1    g703(.A(new_n481), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n737), .A2(new_n329), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n902), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT117), .ZN(G1340gat));
  NOR3_X1   g708(.A1(new_n900), .A2(new_n313), .A3(new_n691), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n904), .A2(new_n905), .A3(new_n690), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n910), .B1(new_n313), .B2(new_n911), .ZN(G1341gat));
  OAI21_X1  g711(.A(KEYINPUT118), .B1(new_n906), .B2(new_n672), .ZN(new_n913));
  INV_X1    g712(.A(G127gat), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT118), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n904), .A2(new_n915), .A3(new_n905), .A4(new_n671), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n913), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n671), .A2(G127gat), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n900), .B2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT119), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n919), .B(new_n920), .ZN(G1342gat));
  OR3_X1    g720(.A1(new_n906), .A2(G134gat), .A3(new_n731), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n922), .A2(KEYINPUT56), .ZN(new_n923));
  OAI21_X1  g722(.A(G134gat), .B1(new_n900), .B2(new_n731), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(KEYINPUT56), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(G1343gat));
  OAI21_X1  g725(.A(new_n463), .B1(new_n894), .B2(new_n896), .ZN(new_n927));
  XOR2_X1   g726(.A(KEYINPUT120), .B(KEYINPUT57), .Z(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n769), .A2(KEYINPUT57), .ZN(new_n930));
  XNOR2_X1  g729(.A(KEYINPUT121), .B(KEYINPUT55), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n931), .B1(new_n876), .B2(new_n879), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n593), .A2(new_n688), .A3(new_n882), .A4(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(new_n888), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n934), .A2(new_n642), .A3(new_n646), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n671), .B1(new_n893), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n930), .B1(new_n936), .B2(new_n896), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT122), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g738(.A(KEYINPUT122), .B(new_n930), .C1(new_n936), .C2(new_n896), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n929), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(new_n708), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n942), .A2(new_n903), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g743(.A(G141gat), .B1(new_n944), .B2(new_n901), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT58), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n942), .A2(new_n479), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n901), .A2(G141gat), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n904), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n945), .A2(new_n946), .A3(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT123), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n941), .A2(new_n738), .A3(new_n943), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(G141gat), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(new_n950), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n952), .B1(new_n955), .B2(KEYINPUT58), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n949), .B1(new_n953), .B2(G141gat), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n957), .A2(KEYINPUT123), .A3(new_n946), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n951), .B1(new_n956), .B2(new_n958), .ZN(G1344gat));
  NAND2_X1  g758(.A1(new_n904), .A2(new_n947), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n960), .A2(G148gat), .A3(new_n691), .ZN(new_n961));
  XOR2_X1   g760(.A(new_n961), .B(KEYINPUT124), .Z(new_n962));
  INV_X1    g761(.A(KEYINPUT59), .ZN(new_n963));
  INV_X1    g762(.A(new_n936), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n673), .A2(new_n901), .A3(new_n691), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n503), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI22_X1  g765(.A1(new_n966), .A2(KEYINPUT57), .B1(new_n927), .B2(new_n928), .ZN(new_n967));
  NAND4_X1  g766(.A1(new_n967), .A2(new_n690), .A3(new_n708), .A4(new_n899), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n963), .B1(new_n968), .B2(G148gat), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n969), .A2(KEYINPUT125), .ZN(new_n970));
  OAI211_X1 g769(.A(new_n963), .B(G148gat), .C1(new_n944), .C2(new_n691), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n971), .B1(new_n969), .B2(KEYINPUT125), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n962), .B1(new_n970), .B2(new_n972), .ZN(G1345gat));
  NOR3_X1   g772(.A1(new_n944), .A2(new_n301), .A3(new_n672), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n960), .A2(new_n672), .ZN(new_n975));
  OR2_X1    g774(.A1(new_n975), .A2(KEYINPUT126), .ZN(new_n976));
  AOI21_X1  g775(.A(G155gat), .B1(new_n975), .B2(KEYINPUT126), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n974), .B1(new_n976), .B2(new_n977), .ZN(G1346gat));
  NAND4_X1  g777(.A1(new_n941), .A2(G162gat), .A3(new_n647), .A4(new_n943), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n302), .B1(new_n960), .B2(new_n731), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n979), .A2(new_n980), .ZN(G1347gat));
  NOR2_X1   g780(.A1(new_n498), .A2(new_n299), .ZN(new_n982));
  INV_X1    g781(.A(new_n982), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n797), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n898), .A2(new_n984), .ZN(new_n985));
  INV_X1    g784(.A(G169gat), .ZN(new_n986));
  NOR3_X1   g785(.A1(new_n985), .A2(new_n986), .A3(new_n901), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n983), .B1(new_n895), .B2(new_n897), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n988), .A2(new_n905), .ZN(new_n989));
  INV_X1    g788(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(new_n738), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n987), .B1(new_n986), .B2(new_n991), .ZN(G1348gat));
  NOR3_X1   g791(.A1(new_n985), .A2(new_n235), .A3(new_n691), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n990), .A2(new_n690), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n993), .B1(new_n241), .B2(new_n994), .ZN(G1349gat));
  OAI21_X1  g794(.A(G183gat), .B1(new_n985), .B2(new_n672), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n671), .A2(new_n255), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n996), .B1(new_n989), .B2(new_n997), .ZN(new_n998));
  XNOR2_X1  g797(.A(new_n998), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g798(.A1(new_n990), .A2(new_n218), .A3(new_n647), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n898), .A2(new_n647), .A3(new_n984), .ZN(new_n1001));
  NOR2_X1   g800(.A1(KEYINPUT127), .A2(KEYINPUT61), .ZN(new_n1002));
  AOI21_X1  g801(.A(new_n218), .B1(KEYINPUT127), .B2(KEYINPUT61), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g803(.A(new_n1004), .ZN(new_n1005));
  AOI21_X1  g804(.A(new_n1002), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n1000), .B1(new_n1005), .B2(new_n1006), .ZN(G1351gat));
  AND2_X1   g806(.A1(new_n988), .A2(new_n947), .ZN(new_n1008));
  AOI21_X1  g807(.A(G197gat), .B1(new_n1008), .B2(new_n738), .ZN(new_n1009));
  AND3_X1   g808(.A1(new_n967), .A2(new_n708), .A3(new_n982), .ZN(new_n1010));
  NOR2_X1   g809(.A1(new_n901), .A2(new_n202), .ZN(new_n1011));
  AOI21_X1  g810(.A(new_n1009), .B1(new_n1010), .B2(new_n1011), .ZN(G1352gat));
  AND3_X1   g811(.A1(new_n1008), .A2(new_n203), .A3(new_n690), .ZN(new_n1013));
  INV_X1    g812(.A(KEYINPUT62), .ZN(new_n1014));
  OR2_X1    g813(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1016));
  AND2_X1   g815(.A1(new_n1010), .A2(new_n690), .ZN(new_n1017));
  OAI211_X1 g816(.A(new_n1015), .B(new_n1016), .C1(new_n1017), .C2(new_n203), .ZN(G1353gat));
  NAND3_X1  g817(.A1(new_n1008), .A2(new_n209), .A3(new_n671), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n1010), .A2(new_n671), .ZN(new_n1020));
  AND3_X1   g819(.A1(new_n1020), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1021));
  AOI21_X1  g820(.A(KEYINPUT63), .B1(new_n1020), .B2(G211gat), .ZN(new_n1022));
  OAI21_X1  g821(.A(new_n1019), .B1(new_n1021), .B2(new_n1022), .ZN(G1354gat));
  NAND3_X1  g822(.A1(new_n1008), .A2(new_n210), .A3(new_n647), .ZN(new_n1024));
  AND2_X1   g823(.A1(new_n1010), .A2(new_n647), .ZN(new_n1025));
  OAI21_X1  g824(.A(new_n1024), .B1(new_n1025), .B2(new_n210), .ZN(G1355gat));
endmodule


