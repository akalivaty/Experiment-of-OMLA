

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588;

  XNOR2_X1 U324 ( .A(n367), .B(n366), .ZN(n408) );
  NOR2_X1 U325 ( .A1(n455), .A2(n533), .ZN(n574) );
  XNOR2_X1 U326 ( .A(n411), .B(KEYINPUT65), .ZN(n412) );
  XNOR2_X1 U327 ( .A(n365), .B(KEYINPUT112), .ZN(n366) );
  XNOR2_X1 U328 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U329 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U330 ( .A(n372), .B(n371), .ZN(n377) );
  XNOR2_X1 U331 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U332 ( .A(n319), .B(n318), .ZN(n452) );
  NOR2_X1 U333 ( .A1(n470), .A2(n421), .ZN(n484) );
  XNOR2_X1 U334 ( .A(n349), .B(n323), .ZN(n324) );
  XNOR2_X1 U335 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U336 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U337 ( .A(n364), .B(n363), .ZN(n577) );
  XNOR2_X1 U338 ( .A(n486), .B(KEYINPUT59), .ZN(n487) );
  XOR2_X1 U339 ( .A(n390), .B(n389), .Z(n573) );
  INV_X1 U340 ( .A(G36GAT), .ZN(n481) );
  XNOR2_X1 U341 ( .A(n488), .B(n487), .ZN(n490) );
  XNOR2_X1 U342 ( .A(n481), .B(KEYINPUT104), .ZN(n482) );
  XNOR2_X1 U343 ( .A(n458), .B(n457), .ZN(G1349GAT) );
  XNOR2_X1 U344 ( .A(n483), .B(n482), .ZN(G1329GAT) );
  XOR2_X1 U345 ( .A(KEYINPUT120), .B(KEYINPUT55), .Z(n440) );
  XOR2_X1 U346 ( .A(KEYINPUT1), .B(G148GAT), .Z(n293) );
  XNOR2_X1 U347 ( .A(G127GAT), .B(G155GAT), .ZN(n292) );
  XNOR2_X1 U348 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U349 ( .A(KEYINPUT92), .B(KEYINPUT94), .Z(n295) );
  XNOR2_X1 U350 ( .A(KEYINPUT6), .B(G57GAT), .ZN(n294) );
  XNOR2_X1 U351 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U352 ( .A(n297), .B(n296), .Z(n304) );
  XOR2_X1 U353 ( .A(G134GAT), .B(G85GAT), .Z(n301) );
  XOR2_X1 U354 ( .A(G141GAT), .B(KEYINPUT89), .Z(n299) );
  XNOR2_X1 U355 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n298) );
  XNOR2_X1 U356 ( .A(n299), .B(n298), .ZN(n428) );
  XNOR2_X1 U357 ( .A(G162GAT), .B(n428), .ZN(n300) );
  XNOR2_X1 U358 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U359 ( .A(G29GAT), .B(n302), .ZN(n303) );
  XNOR2_X1 U360 ( .A(n304), .B(n303), .ZN(n313) );
  XOR2_X1 U361 ( .A(KEYINPUT4), .B(KEYINPUT93), .Z(n306) );
  XNOR2_X1 U362 ( .A(KEYINPUT5), .B(G1GAT), .ZN(n305) );
  XNOR2_X1 U363 ( .A(n306), .B(n305), .ZN(n311) );
  XNOR2_X1 U364 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n307) );
  XNOR2_X1 U365 ( .A(n307), .B(G120GAT), .ZN(n441) );
  XOR2_X1 U366 ( .A(n441), .B(KEYINPUT91), .Z(n309) );
  NAND2_X1 U367 ( .A1(G225GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U368 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U369 ( .A(n311), .B(n310), .Z(n312) );
  XOR2_X1 U370 ( .A(n313), .B(n312), .Z(n470) );
  XOR2_X1 U371 ( .A(G211GAT), .B(G8GAT), .Z(n391) );
  XOR2_X1 U372 ( .A(KEYINPUT21), .B(G197GAT), .Z(n433) );
  XNOR2_X1 U373 ( .A(n391), .B(n433), .ZN(n327) );
  XOR2_X1 U374 ( .A(G169GAT), .B(KEYINPUT18), .Z(n315) );
  XNOR2_X1 U375 ( .A(KEYINPUT17), .B(KEYINPUT86), .ZN(n314) );
  XNOR2_X1 U376 ( .A(n315), .B(n314), .ZN(n319) );
  XNOR2_X1 U377 ( .A(G190GAT), .B(G176GAT), .ZN(n317) );
  INV_X1 U378 ( .A(KEYINPUT19), .ZN(n316) );
  XOR2_X1 U379 ( .A(KEYINPUT82), .B(G36GAT), .Z(n368) );
  XOR2_X1 U380 ( .A(n452), .B(n368), .Z(n321) );
  NAND2_X1 U381 ( .A1(G226GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U382 ( .A(n321), .B(n320), .ZN(n325) );
  XNOR2_X1 U383 ( .A(G92GAT), .B(G64GAT), .ZN(n322) );
  XNOR2_X1 U384 ( .A(n322), .B(G204GAT), .ZN(n349) );
  XOR2_X1 U385 ( .A(G218GAT), .B(G183GAT), .Z(n323) );
  XNOR2_X1 U386 ( .A(n327), .B(n326), .ZN(n530) );
  XOR2_X1 U387 ( .A(KEYINPUT115), .B(KEYINPUT48), .Z(n419) );
  XOR2_X1 U388 ( .A(G1GAT), .B(KEYINPUT71), .Z(n392) );
  XOR2_X1 U389 ( .A(G169GAT), .B(G36GAT), .Z(n329) );
  XNOR2_X1 U390 ( .A(G50GAT), .B(G43GAT), .ZN(n328) );
  XNOR2_X1 U391 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U392 ( .A(n392), .B(n330), .Z(n332) );
  NAND2_X1 U393 ( .A1(G229GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U394 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U395 ( .A(n333), .B(KEYINPUT68), .Z(n336) );
  XNOR2_X1 U396 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n334) );
  XNOR2_X1 U397 ( .A(n334), .B(KEYINPUT7), .ZN(n388) );
  XNOR2_X1 U398 ( .A(n388), .B(KEYINPUT66), .ZN(n335) );
  XNOR2_X1 U399 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U400 ( .A(G197GAT), .B(G22GAT), .Z(n338) );
  XNOR2_X1 U401 ( .A(G113GAT), .B(G15GAT), .ZN(n337) );
  XOR2_X1 U402 ( .A(n338), .B(n337), .Z(n339) );
  XNOR2_X1 U403 ( .A(n340), .B(n339), .ZN(n348) );
  XOR2_X1 U404 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n342) );
  XNOR2_X1 U405 ( .A(KEYINPUT30), .B(KEYINPUT72), .ZN(n341) );
  XNOR2_X1 U406 ( .A(n342), .B(n341), .ZN(n346) );
  XOR2_X1 U407 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n344) );
  XNOR2_X1 U408 ( .A(G141GAT), .B(G8GAT), .ZN(n343) );
  XNOR2_X1 U409 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U410 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U411 ( .A(n348), .B(n347), .ZN(n567) );
  XOR2_X1 U412 ( .A(G85GAT), .B(G99GAT), .Z(n370) );
  XNOR2_X1 U413 ( .A(n349), .B(n370), .ZN(n351) );
  AND2_X1 U414 ( .A1(G230GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U415 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U416 ( .A(KEYINPUT33), .B(n352), .Z(n364) );
  XOR2_X1 U417 ( .A(G71GAT), .B(KEYINPUT13), .Z(n354) );
  XNOR2_X1 U418 ( .A(G57GAT), .B(KEYINPUT74), .ZN(n353) );
  XNOR2_X1 U419 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U420 ( .A(KEYINPUT73), .B(n355), .Z(n405) );
  XOR2_X1 U421 ( .A(KEYINPUT76), .B(KEYINPUT32), .Z(n357) );
  XNOR2_X1 U422 ( .A(G120GAT), .B(G176GAT), .ZN(n356) );
  XNOR2_X1 U423 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U424 ( .A(n405), .B(n358), .ZN(n362) );
  XOR2_X1 U425 ( .A(KEYINPUT75), .B(G78GAT), .Z(n360) );
  XNOR2_X1 U426 ( .A(G148GAT), .B(G106GAT), .ZN(n359) );
  XNOR2_X1 U427 ( .A(n360), .B(n359), .ZN(n431) );
  XNOR2_X1 U428 ( .A(n431), .B(KEYINPUT31), .ZN(n361) );
  XOR2_X1 U429 ( .A(n577), .B(KEYINPUT41), .Z(n514) );
  INV_X1 U430 ( .A(n514), .ZN(n559) );
  NAND2_X1 U431 ( .A1(n567), .A2(n559), .ZN(n367) );
  XOR2_X1 U432 ( .A(KEYINPUT46), .B(KEYINPUT113), .Z(n365) );
  XOR2_X1 U433 ( .A(G134GAT), .B(G43GAT), .Z(n442) );
  XNOR2_X1 U434 ( .A(n442), .B(n368), .ZN(n372) );
  XNOR2_X1 U435 ( .A(KEYINPUT81), .B(KEYINPUT9), .ZN(n369) );
  XOR2_X1 U436 ( .A(KEYINPUT10), .B(G190GAT), .Z(n374) );
  NAND2_X1 U437 ( .A1(G232GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U438 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U439 ( .A(KEYINPUT79), .B(n375), .ZN(n376) );
  XNOR2_X1 U440 ( .A(n377), .B(n376), .ZN(n380) );
  XOR2_X1 U441 ( .A(KEYINPUT11), .B(G92GAT), .Z(n379) );
  XNOR2_X1 U442 ( .A(KEYINPUT80), .B(G106GAT), .ZN(n378) );
  XOR2_X1 U443 ( .A(n379), .B(n378), .Z(n381) );
  NAND2_X1 U444 ( .A1(n380), .A2(n381), .ZN(n385) );
  INV_X1 U445 ( .A(n380), .ZN(n383) );
  INV_X1 U446 ( .A(n381), .ZN(n382) );
  NAND2_X1 U447 ( .A1(n383), .A2(n382), .ZN(n384) );
  NAND2_X1 U448 ( .A1(n385), .A2(n384), .ZN(n390) );
  XOR2_X1 U449 ( .A(G50GAT), .B(KEYINPUT78), .Z(n387) );
  XNOR2_X1 U450 ( .A(G162GAT), .B(G218GAT), .ZN(n386) );
  XNOR2_X1 U451 ( .A(n387), .B(n386), .ZN(n427) );
  XNOR2_X1 U452 ( .A(n427), .B(n388), .ZN(n389) );
  INV_X1 U453 ( .A(n573), .ZN(n491) );
  XOR2_X1 U454 ( .A(n392), .B(n391), .Z(n394) );
  NAND2_X1 U455 ( .A1(G231GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U456 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U457 ( .A(G155GAT), .B(G22GAT), .Z(n434) );
  XOR2_X1 U458 ( .A(n395), .B(n434), .Z(n403) );
  XOR2_X1 U459 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n397) );
  XNOR2_X1 U460 ( .A(G78GAT), .B(G64GAT), .ZN(n396) );
  XNOR2_X1 U461 ( .A(n397), .B(n396), .ZN(n401) );
  XNOR2_X1 U462 ( .A(G127GAT), .B(G15GAT), .ZN(n398) );
  XNOR2_X1 U463 ( .A(n398), .B(G183GAT), .ZN(n446) );
  XNOR2_X1 U464 ( .A(n446), .B(KEYINPUT83), .ZN(n399) );
  XNOR2_X1 U465 ( .A(n399), .B(KEYINPUT12), .ZN(n400) );
  XNOR2_X1 U466 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U467 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U468 ( .A(n405), .B(n404), .ZN(n583) );
  XOR2_X1 U469 ( .A(KEYINPUT111), .B(n583), .Z(n569) );
  INV_X1 U470 ( .A(n569), .ZN(n406) );
  AND2_X1 U471 ( .A1(n491), .A2(n406), .ZN(n407) );
  AND2_X1 U472 ( .A1(n408), .A2(n407), .ZN(n409) );
  XNOR2_X1 U473 ( .A(n409), .B(KEYINPUT47), .ZN(n417) );
  XOR2_X1 U474 ( .A(n573), .B(KEYINPUT101), .Z(n410) );
  XNOR2_X1 U475 ( .A(n410), .B(KEYINPUT36), .ZN(n585) );
  NAND2_X1 U476 ( .A1(n585), .A2(n583), .ZN(n413) );
  XOR2_X1 U477 ( .A(KEYINPUT114), .B(KEYINPUT45), .Z(n411) );
  NOR2_X1 U478 ( .A1(n414), .A2(n567), .ZN(n415) );
  NAND2_X1 U479 ( .A1(n415), .A2(n577), .ZN(n416) );
  NAND2_X1 U480 ( .A1(n417), .A2(n416), .ZN(n418) );
  XNOR2_X1 U481 ( .A(n419), .B(n418), .ZN(n553) );
  INV_X1 U482 ( .A(n553), .ZN(n539) );
  NOR2_X1 U483 ( .A1(n530), .A2(n539), .ZN(n420) );
  XOR2_X1 U484 ( .A(KEYINPUT54), .B(n420), .Z(n421) );
  XOR2_X1 U485 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n423) );
  XNOR2_X1 U486 ( .A(G211GAT), .B(G204GAT), .ZN(n422) );
  XNOR2_X1 U487 ( .A(n423), .B(n422), .ZN(n438) );
  XOR2_X1 U488 ( .A(KEYINPUT88), .B(KEYINPUT90), .Z(n425) );
  NAND2_X1 U489 ( .A1(G228GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U490 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U491 ( .A(n426), .B(KEYINPUT23), .Z(n430) );
  XNOR2_X1 U492 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U493 ( .A(n430), .B(n429), .ZN(n432) );
  XOR2_X1 U494 ( .A(n432), .B(n431), .Z(n436) );
  XNOR2_X1 U495 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U496 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U497 ( .A(n438), .B(n437), .ZN(n472) );
  NAND2_X1 U498 ( .A1(n484), .A2(n472), .ZN(n439) );
  XNOR2_X1 U499 ( .A(n440), .B(n439), .ZN(n455) );
  XOR2_X1 U500 ( .A(n442), .B(n441), .Z(n444) );
  NAND2_X1 U501 ( .A1(G227GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U502 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U503 ( .A(n445), .B(KEYINPUT84), .Z(n448) );
  XNOR2_X1 U504 ( .A(G71GAT), .B(n446), .ZN(n447) );
  XNOR2_X1 U505 ( .A(n448), .B(n447), .ZN(n454) );
  XOR2_X1 U506 ( .A(KEYINPUT20), .B(KEYINPUT85), .Z(n450) );
  XNOR2_X1 U507 ( .A(G99GAT), .B(KEYINPUT64), .ZN(n449) );
  XNOR2_X1 U508 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U509 ( .A(n452), .B(n451), .Z(n453) );
  XOR2_X1 U510 ( .A(n454), .B(n453), .Z(n541) );
  INV_X1 U511 ( .A(n541), .ZN(n533) );
  NAND2_X1 U512 ( .A1(n574), .A2(n559), .ZN(n458) );
  XOR2_X1 U513 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n456) );
  XNOR2_X1 U514 ( .A(n456), .B(G176GAT), .ZN(n457) );
  XOR2_X1 U515 ( .A(KEYINPUT103), .B(KEYINPUT38), .Z(n480) );
  NAND2_X1 U516 ( .A1(n567), .A2(n577), .ZN(n459) );
  XNOR2_X1 U517 ( .A(n459), .B(KEYINPUT77), .ZN(n495) );
  NOR2_X1 U518 ( .A1(n530), .A2(n533), .ZN(n461) );
  INV_X1 U519 ( .A(KEYINPUT96), .ZN(n460) );
  XNOR2_X1 U520 ( .A(n461), .B(n460), .ZN(n462) );
  NAND2_X1 U521 ( .A1(n462), .A2(n472), .ZN(n463) );
  XNOR2_X1 U522 ( .A(n463), .B(KEYINPUT25), .ZN(n467) );
  XNOR2_X1 U523 ( .A(n530), .B(KEYINPUT27), .ZN(n471) );
  NOR2_X1 U524 ( .A1(n541), .A2(n472), .ZN(n465) );
  XNOR2_X1 U525 ( .A(KEYINPUT26), .B(KEYINPUT95), .ZN(n464) );
  XNOR2_X1 U526 ( .A(n465), .B(n464), .ZN(n556) );
  NOR2_X1 U527 ( .A1(n471), .A2(n556), .ZN(n466) );
  NOR2_X1 U528 ( .A1(n467), .A2(n466), .ZN(n468) );
  NOR2_X1 U529 ( .A1(n468), .A2(n470), .ZN(n469) );
  XNOR2_X1 U530 ( .A(n469), .B(KEYINPUT97), .ZN(n475) );
  INV_X1 U531 ( .A(n470), .ZN(n527) );
  NOR2_X1 U532 ( .A1(n527), .A2(n471), .ZN(n554) );
  XNOR2_X1 U533 ( .A(KEYINPUT28), .B(n472), .ZN(n536) );
  NAND2_X1 U534 ( .A1(n554), .A2(n536), .ZN(n540) );
  XOR2_X1 U535 ( .A(KEYINPUT87), .B(n541), .Z(n473) );
  OR2_X1 U536 ( .A1(n540), .A2(n473), .ZN(n474) );
  AND2_X1 U537 ( .A1(n475), .A2(n474), .ZN(n494) );
  NOR2_X1 U538 ( .A1(n494), .A2(n583), .ZN(n476) );
  XNOR2_X1 U539 ( .A(n476), .B(KEYINPUT102), .ZN(n477) );
  NAND2_X1 U540 ( .A1(n477), .A2(n585), .ZN(n478) );
  XNOR2_X1 U541 ( .A(n478), .B(KEYINPUT37), .ZN(n526) );
  NAND2_X1 U542 ( .A1(n495), .A2(n526), .ZN(n479) );
  XNOR2_X1 U543 ( .A(n480), .B(n479), .ZN(n512) );
  NOR2_X1 U544 ( .A1(n530), .A2(n512), .ZN(n483) );
  INV_X1 U545 ( .A(n484), .ZN(n485) );
  NOR2_X1 U546 ( .A1(n556), .A2(n485), .ZN(n586) );
  NAND2_X1 U547 ( .A1(n586), .A2(n567), .ZN(n488) );
  XOR2_X1 U548 ( .A(KEYINPUT60), .B(KEYINPUT124), .Z(n486) );
  XNOR2_X1 U549 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n489) );
  XOR2_X1 U550 ( .A(n490), .B(n489), .Z(G1352GAT) );
  NAND2_X1 U551 ( .A1(n491), .A2(n583), .ZN(n492) );
  XNOR2_X1 U552 ( .A(KEYINPUT16), .B(n492), .ZN(n493) );
  NOR2_X1 U553 ( .A1(n494), .A2(n493), .ZN(n515) );
  NAND2_X1 U554 ( .A1(n495), .A2(n515), .ZN(n504) );
  NOR2_X1 U555 ( .A1(n527), .A2(n504), .ZN(n497) );
  XNOR2_X1 U556 ( .A(KEYINPUT98), .B(KEYINPUT34), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U558 ( .A(G1GAT), .B(n498), .Z(G1324GAT) );
  NOR2_X1 U559 ( .A1(n530), .A2(n504), .ZN(n500) );
  XNOR2_X1 U560 ( .A(G8GAT), .B(KEYINPUT99), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(G1325GAT) );
  NOR2_X1 U562 ( .A1(n533), .A2(n504), .ZN(n502) );
  XNOR2_X1 U563 ( .A(KEYINPUT100), .B(KEYINPUT35), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U565 ( .A(G15GAT), .B(n503), .ZN(G1326GAT) );
  NOR2_X1 U566 ( .A1(n536), .A2(n504), .ZN(n505) );
  XOR2_X1 U567 ( .A(G22GAT), .B(n505), .Z(G1327GAT) );
  NOR2_X1 U568 ( .A1(n512), .A2(n527), .ZN(n506) );
  XNOR2_X1 U569 ( .A(G29GAT), .B(n506), .ZN(n507) );
  XNOR2_X1 U570 ( .A(n507), .B(KEYINPUT39), .ZN(G1328GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n509) );
  XNOR2_X1 U572 ( .A(G43GAT), .B(KEYINPUT106), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(n511) );
  NOR2_X1 U574 ( .A1(n512), .A2(n533), .ZN(n510) );
  XOR2_X1 U575 ( .A(n511), .B(n510), .Z(G1330GAT) );
  NOR2_X1 U576 ( .A1(n536), .A2(n512), .ZN(n513) );
  XOR2_X1 U577 ( .A(G50GAT), .B(n513), .Z(G1331GAT) );
  NOR2_X1 U578 ( .A1(n567), .A2(n514), .ZN(n525) );
  NAND2_X1 U579 ( .A1(n525), .A2(n515), .ZN(n521) );
  NOR2_X1 U580 ( .A1(n527), .A2(n521), .ZN(n516) );
  XOR2_X1 U581 ( .A(G57GAT), .B(n516), .Z(n517) );
  XNOR2_X1 U582 ( .A(KEYINPUT42), .B(n517), .ZN(G1332GAT) );
  NOR2_X1 U583 ( .A1(n530), .A2(n521), .ZN(n519) );
  XNOR2_X1 U584 ( .A(G64GAT), .B(KEYINPUT107), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(G1333GAT) );
  NOR2_X1 U586 ( .A1(n533), .A2(n521), .ZN(n520) );
  XOR2_X1 U587 ( .A(G71GAT), .B(n520), .Z(G1334GAT) );
  NOR2_X1 U588 ( .A1(n536), .A2(n521), .ZN(n523) );
  XNOR2_X1 U589 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n522) );
  XNOR2_X1 U590 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U591 ( .A(G78GAT), .B(n524), .ZN(G1335GAT) );
  NAND2_X1 U592 ( .A1(n526), .A2(n525), .ZN(n535) );
  NOR2_X1 U593 ( .A1(n527), .A2(n535), .ZN(n529) );
  XNOR2_X1 U594 ( .A(G85GAT), .B(KEYINPUT109), .ZN(n528) );
  XNOR2_X1 U595 ( .A(n529), .B(n528), .ZN(G1336GAT) );
  NOR2_X1 U596 ( .A1(n530), .A2(n535), .ZN(n531) );
  XOR2_X1 U597 ( .A(KEYINPUT110), .B(n531), .Z(n532) );
  XNOR2_X1 U598 ( .A(G92GAT), .B(n532), .ZN(G1337GAT) );
  NOR2_X1 U599 ( .A1(n533), .A2(n535), .ZN(n534) );
  XOR2_X1 U600 ( .A(G99GAT), .B(n534), .Z(G1338GAT) );
  NOR2_X1 U601 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U602 ( .A(KEYINPUT44), .B(n537), .Z(n538) );
  XNOR2_X1 U603 ( .A(G106GAT), .B(n538), .ZN(G1339GAT) );
  NOR2_X1 U604 ( .A1(n540), .A2(n539), .ZN(n542) );
  NAND2_X1 U605 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U606 ( .A(KEYINPUT116), .B(n543), .Z(n550) );
  NAND2_X1 U607 ( .A1(n550), .A2(n567), .ZN(n544) );
  XNOR2_X1 U608 ( .A(n544), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n546) );
  NAND2_X1 U610 ( .A1(n550), .A2(n559), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U612 ( .A(G120GAT), .B(n547), .Z(G1341GAT) );
  NAND2_X1 U613 ( .A1(n550), .A2(n569), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n548), .B(KEYINPUT50), .ZN(n549) );
  XNOR2_X1 U615 ( .A(G127GAT), .B(n549), .ZN(G1342GAT) );
  XOR2_X1 U616 ( .A(G134GAT), .B(KEYINPUT51), .Z(n552) );
  NAND2_X1 U617 ( .A1(n550), .A2(n573), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(G1343GAT) );
  XNOR2_X1 U619 ( .A(G141GAT), .B(KEYINPUT118), .ZN(n558) );
  NAND2_X1 U620 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U621 ( .A1(n556), .A2(n555), .ZN(n565) );
  NAND2_X1 U622 ( .A1(n567), .A2(n565), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n558), .B(n557), .ZN(G1344GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT53), .B(KEYINPUT119), .Z(n561) );
  NAND2_X1 U625 ( .A1(n565), .A2(n559), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n561), .B(n560), .ZN(n563) );
  XOR2_X1 U627 ( .A(G148GAT), .B(KEYINPUT52), .Z(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(G1345GAT) );
  NAND2_X1 U629 ( .A1(n583), .A2(n565), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U631 ( .A1(n573), .A2(n565), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U633 ( .A1(n574), .A2(n567), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U635 ( .A1(n569), .A2(n574), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U637 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n571), .B(KEYINPUT121), .ZN(n572) );
  XOR2_X1 U639 ( .A(KEYINPUT122), .B(n572), .Z(n576) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1351GAT) );
  INV_X1 U642 ( .A(n586), .ZN(n578) );
  NOR2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n582) );
  XOR2_X1 U644 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n580) );
  XNOR2_X1 U645 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  NAND2_X1 U648 ( .A1(n583), .A2(n586), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n584), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U651 ( .A(n587), .B(KEYINPUT62), .ZN(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

