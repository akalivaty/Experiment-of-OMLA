

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748;

  NOR2_X1 U370 ( .A1(n531), .A2(n361), .ZN(n360) );
  INV_X2 U371 ( .A(G953), .ZN(n737) );
  XNOR2_X1 U372 ( .A(n735), .B(n397), .ZN(n700) );
  BUF_X1 U373 ( .A(n705), .Z(n716) );
  BUF_X1 U374 ( .A(n615), .Z(n722) );
  XNOR2_X1 U375 ( .A(G116), .B(KEYINPUT3), .ZN(n452) );
  OR2_X1 U376 ( .A1(n689), .A2(n688), .ZN(n690) );
  AND2_X1 U377 ( .A1(n371), .A2(n370), .ZN(n407) );
  XNOR2_X1 U378 ( .A(n375), .B(n414), .ZN(n652) );
  NAND2_X1 U379 ( .A1(n391), .A2(n350), .ZN(n736) );
  XNOR2_X1 U380 ( .A(n696), .B(n695), .ZN(n697) );
  XNOR2_X1 U381 ( .A(n364), .B(n362), .ZN(n717) );
  XNOR2_X1 U382 ( .A(n366), .B(n365), .ZN(n364) );
  XNOR2_X1 U383 ( .A(n452), .B(KEYINPUT71), .ZN(n492) );
  XNOR2_X1 U384 ( .A(n421), .B(G146), .ZN(n455) );
  XNOR2_X1 U385 ( .A(KEYINPUT67), .B(G101), .ZN(n421) );
  XNOR2_X1 U386 ( .A(n383), .B(n530), .ZN(n562) );
  XNOR2_X2 U387 ( .A(n551), .B(KEYINPUT33), .ZN(n675) );
  XNOR2_X1 U388 ( .A(G134), .B(G131), .ZN(n426) );
  XNOR2_X1 U389 ( .A(n611), .B(n392), .ZN(n391) );
  INV_X1 U390 ( .A(KEYINPUT48), .ZN(n392) );
  XNOR2_X1 U391 ( .A(n445), .B(n444), .ZN(n531) );
  XNOR2_X1 U392 ( .A(n367), .B(n457), .ZN(n383) );
  AND2_X2 U393 ( .A1(n410), .A2(n413), .ZN(n705) );
  INV_X1 U394 ( .A(n652), .ZN(n413) );
  NAND2_X1 U395 ( .A1(n407), .A2(n405), .ZN(n410) );
  INV_X1 U396 ( .A(KEYINPUT80), .ZN(n417) );
  NOR2_X1 U397 ( .A1(G953), .A2(G237), .ZN(n477) );
  NAND2_X1 U398 ( .A1(n736), .A2(n411), .ZN(n409) );
  INV_X1 U399 ( .A(KEYINPUT78), .ZN(n393) );
  INV_X1 U400 ( .A(G902), .ZN(n459) );
  XNOR2_X1 U401 ( .A(G146), .B(G125), .ZN(n499) );
  XNOR2_X1 U402 ( .A(n440), .B(KEYINPUT8), .ZN(n464) );
  XNOR2_X1 U403 ( .A(KEYINPUT85), .B(KEYINPUT17), .ZN(n504) );
  XNOR2_X1 U404 ( .A(KEYINPUT18), .B(KEYINPUT82), .ZN(n503) );
  NAND2_X1 U405 ( .A1(G234), .A2(G237), .ZN(n429) );
  NOR2_X1 U406 ( .A1(n592), .A2(n666), .ZN(n387) );
  INV_X1 U407 ( .A(KEYINPUT68), .ZN(n359) );
  XNOR2_X1 U408 ( .A(n369), .B(n368), .ZN(n618) );
  INV_X1 U409 ( .A(n456), .ZN(n368) );
  XNOR2_X1 U410 ( .A(n453), .B(n492), .ZN(n404) );
  XNOR2_X1 U411 ( .A(n497), .B(n496), .ZN(n727) );
  XNOR2_X1 U412 ( .A(n493), .B(n492), .ZN(n497) );
  XNOR2_X1 U413 ( .A(n491), .B(n490), .ZN(n493) );
  XNOR2_X1 U414 ( .A(n499), .B(n439), .ZN(n733) );
  INV_X1 U415 ( .A(KEYINPUT10), .ZN(n439) );
  XNOR2_X1 U416 ( .A(G137), .B(G140), .ZN(n441) );
  XNOR2_X1 U417 ( .A(G119), .B(G110), .ZN(n494) );
  NAND2_X1 U418 ( .A1(n464), .A2(G221), .ZN(n366) );
  XNOR2_X1 U419 ( .A(n438), .B(n436), .ZN(n365) );
  XNOR2_X1 U420 ( .A(G128), .B(KEYINPUT24), .ZN(n437) );
  XNOR2_X1 U421 ( .A(n398), .B(n425), .ZN(n397) );
  XNOR2_X1 U422 ( .A(n455), .B(n399), .ZN(n398) );
  INV_X1 U423 ( .A(KEYINPUT72), .ZN(n414) );
  NOR2_X1 U424 ( .A1(n736), .A2(n616), .ZN(n408) );
  NAND2_X1 U425 ( .A1(n641), .A2(n377), .ZN(n600) );
  AND2_X1 U426 ( .A1(n539), .A2(n378), .ZN(n377) );
  INV_X1 U427 ( .A(n562), .ZN(n378) );
  XNOR2_X1 U428 ( .A(n389), .B(KEYINPUT39), .ZN(n546) );
  NAND2_X1 U429 ( .A1(n353), .A2(n390), .ZN(n389) );
  INV_X1 U430 ( .A(n667), .ZN(n390) );
  NOR2_X1 U431 ( .A1(n600), .A2(n516), .ZN(n602) );
  BUF_X1 U432 ( .A(n531), .Z(n653) );
  INV_X1 U433 ( .A(KEYINPUT1), .ZN(n395) );
  NOR2_X1 U434 ( .A1(n737), .A2(G952), .ZN(n721) );
  XNOR2_X1 U435 ( .A(n385), .B(n384), .ZN(n453) );
  XNOR2_X1 U436 ( .A(G137), .B(G113), .ZN(n384) );
  XNOR2_X1 U437 ( .A(n386), .B(G119), .ZN(n385) );
  INV_X1 U438 ( .A(KEYINPUT5), .ZN(n386) );
  XNOR2_X1 U439 ( .A(n382), .B(KEYINPUT45), .ZN(n615) );
  INV_X1 U440 ( .A(KEYINPUT16), .ZN(n490) );
  XOR2_X1 U441 ( .A(KEYINPUT93), .B(KEYINPUT12), .Z(n476) );
  XNOR2_X1 U442 ( .A(G143), .B(G122), .ZN(n482) );
  XOR2_X1 U443 ( .A(G140), .B(G131), .Z(n479) );
  XNOR2_X1 U444 ( .A(n422), .B(KEYINPUT88), .ZN(n399) );
  INV_X1 U445 ( .A(G110), .ZN(n422) );
  XOR2_X1 U446 ( .A(G107), .B(G104), .Z(n424) );
  INV_X1 U447 ( .A(n441), .ZN(n400) );
  INV_X1 U448 ( .A(n415), .ZN(n406) );
  AND2_X1 U449 ( .A1(n409), .A2(n357), .ZN(n370) );
  AND2_X1 U450 ( .A1(G953), .A2(G902), .ZN(n431) );
  INV_X1 U451 ( .A(G237), .ZN(n458) );
  XNOR2_X1 U452 ( .A(KEYINPUT15), .B(G902), .ZN(n614) );
  BUF_X1 U453 ( .A(n383), .Z(n374) );
  XOR2_X1 U454 ( .A(G122), .B(G107), .Z(n495) );
  INV_X1 U455 ( .A(KEYINPUT9), .ZN(n468) );
  XNOR2_X1 U456 ( .A(n727), .B(n510), .ZN(n693) );
  XNOR2_X1 U457 ( .A(n387), .B(KEYINPUT30), .ZN(n462) );
  NAND2_X1 U458 ( .A1(n394), .A2(n587), .ZN(n451) );
  XNOR2_X1 U459 ( .A(n618), .B(n617), .ZN(n619) );
  XNOR2_X1 U460 ( .A(n733), .B(n363), .ZN(n362) );
  XNOR2_X1 U461 ( .A(n441), .B(n494), .ZN(n363) );
  XNOR2_X1 U462 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U463 ( .A(n388), .B(n548), .ZN(n597) );
  OR2_X1 U464 ( .A1(n379), .A2(n603), .ZN(n604) );
  XNOR2_X1 U465 ( .A(n567), .B(KEYINPUT32), .ZN(n745) );
  NOR2_X1 U466 ( .A1(n595), .A2(n594), .ZN(n636) );
  AND2_X1 U467 ( .A1(n536), .A2(n535), .ZN(n641) );
  XNOR2_X1 U468 ( .A(n703), .B(n420), .ZN(n704) );
  NOR2_X1 U469 ( .A1(n691), .A2(G953), .ZN(n692) );
  XNOR2_X1 U470 ( .A(n635), .B(n402), .ZN(G30) );
  INV_X1 U471 ( .A(G128), .ZN(n402) );
  AND2_X1 U472 ( .A1(n391), .A2(n355), .ZN(n348) );
  XOR2_X1 U473 ( .A(n427), .B(G469), .Z(n349) );
  AND2_X1 U474 ( .A1(n613), .A2(n612), .ZN(n350) );
  AND2_X1 U475 ( .A1(n511), .A2(G210), .ZN(n351) );
  AND2_X1 U476 ( .A1(n580), .A2(n579), .ZN(n352) );
  AND2_X1 U477 ( .A1(n463), .A2(n462), .ZN(n353) );
  NOR2_X1 U478 ( .A1(n609), .A2(n608), .ZN(n354) );
  AND2_X1 U479 ( .A1(n350), .A2(KEYINPUT64), .ZN(n355) );
  OR2_X1 U480 ( .A1(n614), .A2(n616), .ZN(n356) );
  AND2_X1 U481 ( .A1(n356), .A2(n412), .ZN(n411) );
  OR2_X1 U482 ( .A1(n356), .A2(n412), .ZN(n357) );
  NAND2_X1 U483 ( .A1(n518), .A2(n517), .ZN(n520) );
  XNOR2_X2 U484 ( .A(n358), .B(n351), .ZN(n518) );
  NAND2_X1 U485 ( .A1(n693), .A2(n614), .ZN(n358) );
  XNOR2_X2 U486 ( .A(n360), .B(n359), .ZN(n655) );
  INV_X1 U487 ( .A(n588), .ZN(n361) );
  NAND2_X1 U488 ( .A1(n618), .A2(n459), .ZN(n367) );
  XNOR2_X1 U489 ( .A(n404), .B(n403), .ZN(n369) );
  NAND2_X1 U490 ( .A1(n415), .A2(n348), .ZN(n371) );
  XNOR2_X2 U491 ( .A(n381), .B(n393), .ZN(n415) );
  INV_X1 U492 ( .A(n502), .ZN(n498) );
  XNOR2_X1 U493 ( .A(n467), .B(KEYINPUT4), .ZN(n502) );
  XNOR2_X2 U494 ( .A(G143), .B(G128), .ZN(n467) );
  INV_X2 U495 ( .A(G113), .ZN(n372) );
  XNOR2_X2 U496 ( .A(n372), .B(G104), .ZN(n491) );
  XNOR2_X1 U497 ( .A(n373), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U498 ( .A1(n699), .A2(n721), .ZN(n373) );
  NAND2_X1 U499 ( .A1(n408), .A2(n722), .ZN(n375) );
  NAND2_X1 U500 ( .A1(n376), .A2(n610), .ZN(n611) );
  AND2_X1 U501 ( .A1(n354), .A2(n746), .ZN(n376) );
  XNOR2_X1 U502 ( .A(n486), .B(n487), .ZN(n489) );
  NOR2_X2 U503 ( .A1(n621), .A2(n721), .ZN(n623) );
  XNOR2_X1 U504 ( .A(n602), .B(n601), .ZN(n379) );
  NAND2_X1 U505 ( .A1(n584), .A2(n583), .ZN(n382) );
  NAND2_X1 U506 ( .A1(n615), .A2(n585), .ZN(n381) );
  NAND2_X1 U507 ( .A1(n705), .A2(G475), .ZN(n709) );
  NAND2_X1 U508 ( .A1(n416), .A2(n352), .ZN(n418) );
  XNOR2_X1 U509 ( .A(n418), .B(n417), .ZN(n584) );
  XNOR2_X1 U510 ( .A(n380), .B(n711), .ZN(G60) );
  NOR2_X2 U511 ( .A1(n710), .A2(n721), .ZN(n380) );
  NAND2_X1 U512 ( .A1(n394), .A2(n374), .ZN(n572) );
  XNOR2_X1 U513 ( .A(n383), .B(KEYINPUT100), .ZN(n592) );
  NOR2_X1 U514 ( .A1(n655), .A2(n374), .ZN(n569) );
  NAND2_X1 U515 ( .A1(n658), .A2(n374), .ZN(n659) );
  NAND2_X1 U516 ( .A1(n546), .A2(n641), .ZN(n388) );
  INV_X1 U517 ( .A(n396), .ZN(n394) );
  XNOR2_X2 U518 ( .A(n396), .B(n395), .ZN(n561) );
  XNOR2_X1 U519 ( .A(n396), .B(KEYINPUT104), .ZN(n594) );
  XNOR2_X2 U520 ( .A(n428), .B(n349), .ZN(n396) );
  XNOR2_X2 U521 ( .A(n456), .B(n400), .ZN(n735) );
  XNOR2_X2 U522 ( .A(n498), .B(n426), .ZN(n456) );
  NAND2_X1 U523 ( .A1(n401), .A2(KEYINPUT44), .ZN(n416) );
  NAND2_X1 U524 ( .A1(n568), .A2(n745), .ZN(n401) );
  INV_X1 U525 ( .A(n401), .ZN(n581) );
  NAND2_X1 U526 ( .A1(n717), .A2(n459), .ZN(n445) );
  XNOR2_X1 U527 ( .A(n455), .B(n454), .ZN(n403) );
  INV_X1 U528 ( .A(n518), .ZN(n516) );
  NAND2_X1 U529 ( .A1(n406), .A2(n411), .ZN(n405) );
  INV_X1 U530 ( .A(KEYINPUT64), .ZN(n412) );
  NAND2_X1 U531 ( .A1(n574), .A2(n675), .ZN(n553) );
  NOR2_X1 U532 ( .A1(n667), .A2(n666), .ZN(n419) );
  XOR2_X1 U533 ( .A(n702), .B(n701), .Z(n420) );
  XNOR2_X1 U534 ( .A(n469), .B(n468), .ZN(n470) );
  BUF_X1 U535 ( .A(n693), .Z(n696) );
  INV_X1 U536 ( .A(KEYINPUT34), .ZN(n552) );
  NAND2_X1 U537 ( .A1(G227), .A2(n737), .ZN(n423) );
  XNOR2_X1 U538 ( .A(n424), .B(n423), .ZN(n425) );
  NOR2_X2 U539 ( .A1(G902), .A2(n700), .ZN(n428) );
  XNOR2_X1 U540 ( .A(KEYINPUT70), .B(KEYINPUT69), .ZN(n427) );
  XNOR2_X1 U541 ( .A(n429), .B(KEYINPUT87), .ZN(n430) );
  XOR2_X1 U542 ( .A(KEYINPUT14), .B(n430), .Z(n433) );
  NAND2_X1 U543 ( .A1(n433), .A2(n431), .ZN(n521) );
  XNOR2_X1 U544 ( .A(KEYINPUT102), .B(n521), .ZN(n432) );
  NOR2_X1 U545 ( .A1(G900), .A2(n432), .ZN(n434) );
  NAND2_X1 U546 ( .A1(G952), .A2(n433), .ZN(n684) );
  NOR2_X1 U547 ( .A1(n684), .A2(G953), .ZN(n523) );
  OR2_X1 U548 ( .A1(n434), .A2(n523), .ZN(n435) );
  XNOR2_X1 U549 ( .A(n435), .B(KEYINPUT76), .ZN(n587) );
  XNOR2_X1 U550 ( .A(KEYINPUT89), .B(KEYINPUT23), .ZN(n436) );
  XNOR2_X1 U551 ( .A(n437), .B(KEYINPUT73), .ZN(n438) );
  AND2_X1 U552 ( .A1(G234), .A2(n737), .ZN(n440) );
  NAND2_X1 U553 ( .A1(n614), .A2(G234), .ZN(n442) );
  XNOR2_X1 U554 ( .A(n442), .B(KEYINPUT20), .ZN(n446) );
  NAND2_X1 U555 ( .A1(n446), .A2(G217), .ZN(n443) );
  XNOR2_X1 U556 ( .A(n443), .B(KEYINPUT25), .ZN(n444) );
  INV_X1 U557 ( .A(n446), .ZN(n448) );
  INV_X1 U558 ( .A(G221), .ZN(n447) );
  OR2_X1 U559 ( .A1(n448), .A2(n447), .ZN(n450) );
  INV_X1 U560 ( .A(KEYINPUT21), .ZN(n449) );
  XNOR2_X1 U561 ( .A(n450), .B(n449), .ZN(n588) );
  NOR2_X1 U562 ( .A1(n451), .A2(n655), .ZN(n463) );
  NAND2_X1 U563 ( .A1(n477), .A2(G210), .ZN(n454) );
  XOR2_X1 U564 ( .A(G472), .B(KEYINPUT90), .Z(n457) );
  NAND2_X1 U565 ( .A1(n459), .A2(n458), .ZN(n511) );
  NAND2_X1 U566 ( .A1(n511), .A2(G214), .ZN(n461) );
  INV_X1 U567 ( .A(KEYINPUT86), .ZN(n460) );
  XNOR2_X1 U568 ( .A(n461), .B(n460), .ZN(n666) );
  XNOR2_X1 U569 ( .A(G134), .B(n495), .ZN(n473) );
  XOR2_X1 U570 ( .A(KEYINPUT96), .B(KEYINPUT7), .Z(n466) );
  NAND2_X1 U571 ( .A1(G217), .A2(n464), .ZN(n465) );
  XNOR2_X1 U572 ( .A(n466), .B(n465), .ZN(n471) );
  XOR2_X1 U573 ( .A(n467), .B(G116), .Z(n469) );
  XNOR2_X1 U574 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U575 ( .A(n473), .B(n472), .ZN(n712) );
  NOR2_X1 U576 ( .A1(n712), .A2(G902), .ZN(n474) );
  XNOR2_X1 U577 ( .A(n474), .B(G478), .ZN(n536) );
  XNOR2_X1 U578 ( .A(KEYINPUT94), .B(KEYINPUT13), .ZN(n487) );
  XNOR2_X1 U579 ( .A(KEYINPUT11), .B(KEYINPUT92), .ZN(n475) );
  XNOR2_X1 U580 ( .A(n476), .B(n475), .ZN(n481) );
  NAND2_X1 U581 ( .A1(G214), .A2(n477), .ZN(n478) );
  XNOR2_X1 U582 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U583 ( .A(n481), .B(n480), .ZN(n485) );
  XNOR2_X1 U584 ( .A(n491), .B(n482), .ZN(n483) );
  XNOR2_X1 U585 ( .A(n483), .B(n733), .ZN(n484) );
  XNOR2_X1 U586 ( .A(n485), .B(n484), .ZN(n707) );
  NOR2_X1 U587 ( .A1(G902), .A2(n707), .ZN(n486) );
  INV_X1 U588 ( .A(G475), .ZN(n488) );
  XNOR2_X1 U589 ( .A(n489), .B(n488), .ZN(n526) );
  OR2_X1 U590 ( .A1(n536), .A2(n526), .ZN(n554) );
  XNOR2_X1 U591 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U592 ( .A(KEYINPUT67), .B(G101), .Z(n500) );
  XNOR2_X1 U593 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U594 ( .A(n502), .B(n501), .ZN(n509) );
  XNOR2_X1 U595 ( .A(n504), .B(n503), .ZN(n507) );
  NAND2_X1 U596 ( .A1(n737), .A2(G224), .ZN(n505) );
  XNOR2_X1 U597 ( .A(n505), .B(KEYINPUT74), .ZN(n506) );
  XNOR2_X1 U598 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U599 ( .A(n509), .B(n508), .ZN(n510) );
  NOR2_X1 U600 ( .A1(n554), .A2(n516), .ZN(n512) );
  AND2_X1 U601 ( .A1(n353), .A2(n512), .ZN(n608) );
  XOR2_X1 U602 ( .A(G143), .B(n608), .Z(G45) );
  XNOR2_X1 U603 ( .A(n526), .B(KEYINPUT95), .ZN(n535) );
  NOR2_X1 U604 ( .A1(n535), .A2(n536), .ZN(n513) );
  XNOR2_X1 U605 ( .A(n513), .B(KEYINPUT97), .ZN(n627) );
  XNOR2_X1 U606 ( .A(n627), .B(KEYINPUT98), .ZN(n577) );
  INV_X1 U607 ( .A(n577), .ZN(n515) );
  INV_X1 U608 ( .A(KEYINPUT38), .ZN(n514) );
  XNOR2_X1 U609 ( .A(n516), .B(n514), .ZN(n667) );
  NAND2_X1 U610 ( .A1(n515), .A2(n546), .ZN(n613) );
  XNOR2_X1 U611 ( .A(n613), .B(G134), .ZN(G36) );
  INV_X1 U612 ( .A(n666), .ZN(n517) );
  INV_X1 U613 ( .A(KEYINPUT19), .ZN(n519) );
  XNOR2_X2 U614 ( .A(n520), .B(n519), .ZN(n637) );
  NOR2_X1 U615 ( .A1(n521), .A2(G898), .ZN(n522) );
  NOR2_X1 U616 ( .A1(n523), .A2(n522), .ZN(n524) );
  NOR2_X2 U617 ( .A1(n637), .A2(n524), .ZN(n525) );
  XNOR2_X2 U618 ( .A(n525), .B(KEYINPUT0), .ZN(n574) );
  AND2_X1 U619 ( .A1(n536), .A2(n526), .ZN(n669) );
  AND2_X1 U620 ( .A1(n669), .A2(n588), .ZN(n527) );
  NAND2_X1 U621 ( .A1(n574), .A2(n527), .ZN(n529) );
  XNOR2_X1 U622 ( .A(KEYINPUT65), .B(KEYINPUT22), .ZN(n528) );
  XNOR2_X2 U623 ( .A(n529), .B(n528), .ZN(n565) );
  INV_X1 U624 ( .A(n561), .ZN(n656) );
  XNOR2_X1 U625 ( .A(KEYINPUT99), .B(KEYINPUT6), .ZN(n530) );
  INV_X1 U626 ( .A(n653), .ZN(n532) );
  NAND2_X1 U627 ( .A1(n562), .A2(n532), .ZN(n533) );
  NOR2_X1 U628 ( .A1(n561), .A2(n533), .ZN(n534) );
  NAND2_X1 U629 ( .A1(n565), .A2(n534), .ZN(n579) );
  XNOR2_X1 U630 ( .A(n579), .B(G101), .ZN(G3) );
  AND2_X1 U631 ( .A1(n588), .A2(n517), .ZN(n537) );
  AND2_X1 U632 ( .A1(n587), .A2(n537), .ZN(n538) );
  AND2_X1 U633 ( .A1(n538), .A2(n653), .ZN(n539) );
  XNOR2_X1 U634 ( .A(KEYINPUT103), .B(n600), .ZN(n540) );
  NAND2_X1 U635 ( .A1(n656), .A2(n540), .ZN(n541) );
  XNOR2_X1 U636 ( .A(n541), .B(KEYINPUT43), .ZN(n542) );
  NAND2_X1 U637 ( .A1(n542), .A2(n516), .ZN(n612) );
  XNOR2_X1 U638 ( .A(n612), .B(G140), .ZN(G42) );
  NAND2_X1 U639 ( .A1(n592), .A2(n653), .ZN(n543) );
  NOR2_X1 U640 ( .A1(n561), .A2(n543), .ZN(n544) );
  NAND2_X1 U641 ( .A1(n565), .A2(n544), .ZN(n545) );
  XNOR2_X1 U642 ( .A(n545), .B(KEYINPUT101), .ZN(n559) );
  XOR2_X1 U643 ( .A(n559), .B(G110), .Z(G12) );
  INV_X1 U644 ( .A(KEYINPUT105), .ZN(n547) );
  XNOR2_X1 U645 ( .A(n547), .B(KEYINPUT40), .ZN(n548) );
  XNOR2_X1 U646 ( .A(G131), .B(KEYINPUT126), .ZN(n549) );
  XNOR2_X1 U647 ( .A(n597), .B(n549), .ZN(G33) );
  NOR2_X1 U648 ( .A1(n562), .A2(n655), .ZN(n550) );
  NAND2_X1 U649 ( .A1(n561), .A2(n550), .ZN(n551) );
  XNOR2_X1 U650 ( .A(n553), .B(n552), .ZN(n556) );
  INV_X1 U651 ( .A(n554), .ZN(n555) );
  NAND2_X1 U652 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U653 ( .A(n557), .B(KEYINPUT35), .ZN(n560) );
  XNOR2_X1 U654 ( .A(G122), .B(KEYINPUT125), .ZN(n558) );
  XNOR2_X1 U655 ( .A(n560), .B(n558), .ZN(G24) );
  NOR2_X1 U656 ( .A1(n560), .A2(n559), .ZN(n568) );
  XNOR2_X1 U657 ( .A(n561), .B(KEYINPUT83), .ZN(n603) );
  NAND2_X1 U658 ( .A1(n562), .A2(n653), .ZN(n563) );
  OR2_X1 U659 ( .A1(n603), .A2(n563), .ZN(n564) );
  XNOR2_X1 U660 ( .A(n564), .B(KEYINPUT75), .ZN(n566) );
  NAND2_X1 U661 ( .A1(n566), .A2(n565), .ZN(n567) );
  INV_X1 U662 ( .A(KEYINPUT44), .ZN(n582) );
  AND2_X1 U663 ( .A1(n561), .A2(n569), .ZN(n662) );
  NAND2_X1 U664 ( .A1(n662), .A2(n574), .ZN(n571) );
  XOR2_X1 U665 ( .A(KEYINPUT91), .B(KEYINPUT31), .Z(n570) );
  XNOR2_X1 U666 ( .A(n571), .B(n570), .ZN(n644) );
  INV_X1 U667 ( .A(n644), .ZN(n575) );
  NOR2_X1 U668 ( .A1(n572), .A2(n655), .ZN(n573) );
  NAND2_X1 U669 ( .A1(n574), .A2(n573), .ZN(n624) );
  NAND2_X1 U670 ( .A1(n575), .A2(n624), .ZN(n578) );
  INV_X1 U671 ( .A(n641), .ZN(n576) );
  NAND2_X1 U672 ( .A1(n577), .A2(n576), .ZN(n671) );
  NAND2_X1 U673 ( .A1(n578), .A2(n671), .ZN(n580) );
  NAND2_X1 U674 ( .A1(n581), .A2(n582), .ZN(n583) );
  INV_X1 U675 ( .A(n614), .ZN(n585) );
  NAND2_X1 U676 ( .A1(n419), .A2(n669), .ZN(n586) );
  XNOR2_X1 U677 ( .A(KEYINPUT41), .B(n586), .ZN(n685) );
  INV_X1 U678 ( .A(n587), .ZN(n589) );
  NOR2_X1 U679 ( .A1(n589), .A2(n361), .ZN(n590) );
  NAND2_X1 U680 ( .A1(n590), .A2(n653), .ZN(n591) );
  NOR2_X1 U681 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U682 ( .A(KEYINPUT28), .B(n593), .Z(n595) );
  NAND2_X1 U683 ( .A1(n685), .A2(n636), .ZN(n596) );
  XNOR2_X1 U684 ( .A(n596), .B(KEYINPUT42), .ZN(n748) );
  NAND2_X1 U685 ( .A1(n748), .A2(n597), .ZN(n599) );
  XNOR2_X1 U686 ( .A(KEYINPUT79), .B(KEYINPUT46), .ZN(n598) );
  XNOR2_X1 U687 ( .A(n599), .B(n598), .ZN(n610) );
  INV_X1 U688 ( .A(KEYINPUT36), .ZN(n601) );
  XNOR2_X1 U689 ( .A(n604), .B(KEYINPUT106), .ZN(n746) );
  INV_X1 U690 ( .A(n637), .ZN(n605) );
  AND2_X1 U691 ( .A1(n636), .A2(n605), .ZN(n606) );
  NAND2_X1 U692 ( .A1(n671), .A2(n606), .ZN(n607) );
  XNOR2_X1 U693 ( .A(n607), .B(KEYINPUT47), .ZN(n609) );
  INV_X1 U694 ( .A(KEYINPUT2), .ZN(n616) );
  NAND2_X1 U695 ( .A1(n705), .A2(G472), .ZN(n620) );
  XNOR2_X1 U696 ( .A(KEYINPUT107), .B(KEYINPUT62), .ZN(n617) );
  XNOR2_X1 U697 ( .A(n620), .B(n619), .ZN(n621) );
  XNOR2_X1 U698 ( .A(KEYINPUT81), .B(KEYINPUT63), .ZN(n622) );
  XNOR2_X1 U699 ( .A(n623), .B(n622), .ZN(G57) );
  INV_X1 U700 ( .A(n624), .ZN(n628) );
  NAND2_X1 U701 ( .A1(n628), .A2(n641), .ZN(n625) );
  XNOR2_X1 U702 ( .A(n625), .B(KEYINPUT108), .ZN(n626) );
  XNOR2_X1 U703 ( .A(G104), .B(n626), .ZN(G6) );
  XOR2_X1 U704 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n630) );
  INV_X1 U705 ( .A(n627), .ZN(n643) );
  NAND2_X1 U706 ( .A1(n628), .A2(n643), .ZN(n629) );
  XNOR2_X1 U707 ( .A(n630), .B(n629), .ZN(n631) );
  XNOR2_X1 U708 ( .A(G107), .B(n631), .ZN(G9) );
  NAND2_X1 U709 ( .A1(n643), .A2(n636), .ZN(n632) );
  NOR2_X1 U710 ( .A1(n632), .A2(n637), .ZN(n634) );
  XNOR2_X1 U711 ( .A(KEYINPUT29), .B(KEYINPUT109), .ZN(n633) );
  XNOR2_X1 U712 ( .A(n634), .B(n633), .ZN(n635) );
  NAND2_X1 U713 ( .A1(n636), .A2(n641), .ZN(n638) );
  NOR2_X1 U714 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U715 ( .A(KEYINPUT110), .B(n639), .Z(n640) );
  XNOR2_X1 U716 ( .A(G146), .B(n640), .ZN(G48) );
  NAND2_X1 U717 ( .A1(n644), .A2(n641), .ZN(n642) );
  XNOR2_X1 U718 ( .A(n642), .B(G113), .ZN(G15) );
  XOR2_X1 U719 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n646) );
  NAND2_X1 U720 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U721 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U722 ( .A(G116), .B(n647), .ZN(G18) );
  INV_X1 U723 ( .A(n722), .ZN(n648) );
  NOR2_X1 U724 ( .A1(n648), .A2(n736), .ZN(n650) );
  XOR2_X1 U725 ( .A(KEYINPUT2), .B(KEYINPUT77), .Z(n649) );
  NOR2_X1 U726 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U727 ( .A1(n652), .A2(n651), .ZN(n689) );
  NAND2_X1 U728 ( .A1(n653), .A2(n361), .ZN(n654) );
  XNOR2_X1 U729 ( .A(n654), .B(KEYINPUT49), .ZN(n660) );
  NAND2_X1 U730 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U731 ( .A(KEYINPUT50), .B(n657), .ZN(n658) );
  NOR2_X1 U732 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U733 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U734 ( .A(KEYINPUT51), .B(n663), .ZN(n664) );
  NAND2_X1 U735 ( .A1(n664), .A2(n685), .ZN(n665) );
  XNOR2_X1 U736 ( .A(KEYINPUT113), .B(n665), .ZN(n680) );
  NAND2_X1 U737 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U738 ( .A(KEYINPUT114), .B(n668), .ZN(n670) );
  NAND2_X1 U739 ( .A1(n670), .A2(n669), .ZN(n673) );
  NAND2_X1 U740 ( .A1(n419), .A2(n671), .ZN(n672) );
  NAND2_X1 U741 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U742 ( .A(KEYINPUT115), .B(n674), .ZN(n677) );
  INV_X1 U743 ( .A(n675), .ZN(n676) );
  NOR2_X1 U744 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U745 ( .A(n678), .B(KEYINPUT116), .ZN(n679) );
  NOR2_X1 U746 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U747 ( .A(n681), .B(KEYINPUT52), .Z(n682) );
  XNOR2_X1 U748 ( .A(KEYINPUT117), .B(n682), .ZN(n683) );
  NOR2_X1 U749 ( .A1(n684), .A2(n683), .ZN(n687) );
  AND2_X1 U750 ( .A1(n675), .A2(n685), .ZN(n686) );
  OR2_X1 U751 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U752 ( .A(KEYINPUT118), .B(n690), .ZN(n691) );
  XNOR2_X1 U753 ( .A(n692), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U754 ( .A1(n705), .A2(G210), .ZN(n698) );
  XNOR2_X1 U755 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n694) );
  XOR2_X1 U756 ( .A(n694), .B(KEYINPUT55), .Z(n695) );
  XNOR2_X1 U757 ( .A(n698), .B(n697), .ZN(n699) );
  NAND2_X1 U758 ( .A1(n716), .A2(G469), .ZN(n703) );
  XNOR2_X1 U759 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n702) );
  XNOR2_X1 U760 ( .A(n700), .B(KEYINPUT57), .ZN(n701) );
  NOR2_X1 U761 ( .A1(n721), .A2(n704), .ZN(G54) );
  XOR2_X1 U762 ( .A(KEYINPUT59), .B(KEYINPUT84), .Z(n706) );
  XNOR2_X1 U763 ( .A(n709), .B(n708), .ZN(n710) );
  XNOR2_X1 U764 ( .A(KEYINPUT60), .B(KEYINPUT66), .ZN(n711) );
  NAND2_X1 U765 ( .A1(n716), .A2(G478), .ZN(n714) );
  XOR2_X1 U766 ( .A(n712), .B(KEYINPUT121), .Z(n713) );
  XNOR2_X1 U767 ( .A(n714), .B(n713), .ZN(n715) );
  NOR2_X1 U768 ( .A1(n721), .A2(n715), .ZN(G63) );
  NAND2_X1 U769 ( .A1(n716), .A2(G217), .ZN(n719) );
  XOR2_X1 U770 ( .A(KEYINPUT122), .B(n717), .Z(n718) );
  XNOR2_X1 U771 ( .A(n719), .B(n718), .ZN(n720) );
  NOR2_X1 U772 ( .A1(n721), .A2(n720), .ZN(G66) );
  NAND2_X1 U773 ( .A1(n722), .A2(n737), .ZN(n726) );
  NAND2_X1 U774 ( .A1(G953), .A2(G224), .ZN(n723) );
  XNOR2_X1 U775 ( .A(KEYINPUT61), .B(n723), .ZN(n724) );
  NAND2_X1 U776 ( .A1(n724), .A2(G898), .ZN(n725) );
  NAND2_X1 U777 ( .A1(n726), .A2(n725), .ZN(n732) );
  BUF_X1 U778 ( .A(n727), .Z(n728) );
  XNOR2_X1 U779 ( .A(n728), .B(G101), .ZN(n730) );
  NOR2_X1 U780 ( .A1(n737), .A2(G898), .ZN(n729) );
  NOR2_X1 U781 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U782 ( .A(n732), .B(n731), .ZN(G69) );
  XOR2_X1 U783 ( .A(KEYINPUT123), .B(n733), .Z(n734) );
  XNOR2_X1 U784 ( .A(n735), .B(n734), .ZN(n740) );
  XNOR2_X1 U785 ( .A(n736), .B(n740), .ZN(n738) );
  NAND2_X1 U786 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U787 ( .A(n739), .B(KEYINPUT124), .ZN(n744) );
  XNOR2_X1 U788 ( .A(G227), .B(n740), .ZN(n741) );
  NAND2_X1 U789 ( .A1(n741), .A2(G900), .ZN(n742) );
  NAND2_X1 U790 ( .A1(n742), .A2(G953), .ZN(n743) );
  NAND2_X1 U791 ( .A1(n744), .A2(n743), .ZN(G72) );
  XNOR2_X1 U792 ( .A(G119), .B(n745), .ZN(G21) );
  XOR2_X1 U793 ( .A(G125), .B(n746), .Z(n747) );
  XNOR2_X1 U794 ( .A(KEYINPUT37), .B(n747), .ZN(G27) );
  XNOR2_X1 U795 ( .A(G137), .B(n748), .ZN(G39) );
endmodule

