//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 0 0 0 1 1 0 1 1 0 0 0 0 1 0 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 1 1 0 1 1 0 0 1 0 0 1 0 1 0 0 1 0 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:05 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n558, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n847, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1264, new_n1265;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n459), .A2(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G101), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(new_n459), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n461), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n465), .A2(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n466), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n469), .A2(new_n472), .ZN(G160));
  AND2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(KEYINPUT66), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n467), .A2(new_n479), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n466), .B1(new_n463), .B2(new_n464), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  XOR2_X1   g059(.A(new_n484), .B(KEYINPUT67), .Z(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n482), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  OAI211_X1 g064(.A(G126), .B(G2105), .C1(new_n474), .C2(new_n475), .ZN(new_n490));
  OR2_X1    g065(.A1(KEYINPUT68), .A2(G114), .ZN(new_n491));
  NAND2_X1  g066(.A1(KEYINPUT68), .A2(G114), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n466), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n490), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g070(.A(G138), .B(new_n466), .C1(new_n474), .C2(new_n475), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n465), .A2(new_n498), .A3(G138), .A4(new_n466), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n495), .B1(new_n497), .B2(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT69), .ZN(new_n501));
  AND2_X1   g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G62), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT5), .B(G543), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(KEYINPUT69), .A3(G62), .ZN(new_n508));
  NAND2_X1  g083(.A1(G75), .A2(G543), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n506), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G651), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n507), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n512));
  AND2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OR2_X1    g090(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n511), .A2(new_n516), .ZN(G166));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  XOR2_X1   g093(.A(new_n518), .B(KEYINPUT7), .Z(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  XOR2_X1   g095(.A(KEYINPUT71), .B(G89), .Z(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT6), .B(G651), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n521), .A2(new_n522), .B1(G63), .B2(G651), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n520), .B1(new_n523), .B2(new_n504), .ZN(new_n524));
  OR2_X1    g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT70), .ZN(new_n526));
  NAND2_X1  g101(.A1(KEYINPUT6), .A2(G651), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  OAI21_X1  g103(.A(KEYINPUT70), .B1(new_n513), .B2(new_n514), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n528), .A2(new_n529), .A3(G543), .ZN(new_n530));
  INV_X1    g105(.A(G51), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n524), .A2(new_n532), .ZN(G168));
  INV_X1    g108(.A(G543), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n534), .B1(new_n522), .B2(KEYINPUT70), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n535), .A2(G52), .A3(new_n528), .ZN(new_n536));
  NAND2_X1  g111(.A1(G77), .A2(G543), .ZN(new_n537));
  INV_X1    g112(.A(G64), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n504), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G651), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n515), .A2(new_n504), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G90), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n536), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT72), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n543), .A2(KEYINPUT72), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n545), .A2(new_n546), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  AOI22_X1  g123(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G651), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AND3_X1   g126(.A1(new_n528), .A2(new_n529), .A3(G543), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G43), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n541), .A2(G81), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n551), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n558));
  XOR2_X1   g133(.A(new_n558), .B(KEYINPUT73), .Z(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  NAND4_X1  g137(.A1(new_n528), .A2(new_n529), .A3(G53), .A4(G543), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(KEYINPUT9), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n535), .A2(new_n565), .A3(G53), .A4(new_n528), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n504), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(G651), .A2(new_n570), .B1(new_n541), .B2(G91), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT74), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n567), .A2(KEYINPUT74), .A3(new_n571), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G299));
  INV_X1    g152(.A(G168), .ZN(G286));
  NAND2_X1  g153(.A1(new_n511), .A2(new_n516), .ZN(G303));
  NAND2_X1  g154(.A1(new_n552), .A2(G49), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n541), .A2(G87), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(G288));
  AOI22_X1  g158(.A1(new_n507), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n550), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n507), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(new_n515), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n585), .A2(new_n587), .ZN(G305));
  INV_X1    g163(.A(G60), .ZN(new_n589));
  INV_X1    g164(.A(G72), .ZN(new_n590));
  OAI22_X1  g165(.A1(new_n504), .A2(new_n589), .B1(new_n590), .B2(new_n534), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT75), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI221_X1 g168(.A(KEYINPUT75), .B1(new_n590), .B2(new_n534), .C1(new_n504), .C2(new_n589), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n593), .A2(G651), .A3(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n552), .A2(G47), .B1(new_n541), .B2(G85), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(new_n507), .A2(new_n522), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  OAI21_X1  g174(.A(KEYINPUT76), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT76), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n507), .A2(new_n522), .A3(new_n601), .A4(G92), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n600), .A2(KEYINPUT10), .A3(new_n602), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n504), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n552), .A2(G54), .B1(G651), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n605), .A2(new_n606), .A3(new_n610), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n612), .B1(G171), .B2(G868), .ZN(G321));
  XNOR2_X1  g188(.A(G321), .B(KEYINPUT77), .ZN(G284));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(new_n576), .B2(G868), .ZN(G297));
  OAI21_X1  g191(.A(new_n615), .B1(new_n576), .B2(G868), .ZN(G280));
  AND3_X1   g192(.A1(new_n605), .A2(new_n606), .A3(new_n610), .ZN(new_n618));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(G860), .ZN(G148));
  NOR2_X1   g195(.A1(new_n555), .A2(G868), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n611), .A2(G559), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT78), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n621), .B1(new_n623), .B2(G868), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n481), .A2(G135), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT79), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n483), .A2(G123), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT80), .ZN(new_n630));
  OAI21_X1  g205(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n631));
  INV_X1    g206(.A(G111), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n631), .B1(new_n632), .B2(G2105), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n628), .A2(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(G2096), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n635), .A2(G2096), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n465), .A2(new_n460), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT12), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT13), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2100), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n638), .A2(new_n639), .A3(new_n643), .ZN(G156));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT81), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2427), .B(G2430), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n647), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(KEYINPUT14), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2451), .B(G2454), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1341), .B(G1348), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n654), .B(new_n655), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n652), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2443), .B(G2446), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  AND2_X1   g234(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g235(.A(G14), .B1(new_n657), .B2(new_n659), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(G401));
  NOR2_X1   g237(.A1(G2072), .A2(G2078), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n442), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT17), .Z(new_n665));
  XNOR2_X1  g240(.A(G2084), .B(G2090), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT82), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT83), .Z(new_n669));
  NAND3_X1  g244(.A1(new_n665), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT84), .Z(new_n671));
  NAND3_X1  g246(.A1(new_n667), .A2(new_n664), .A3(new_n668), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT18), .Z(new_n673));
  INV_X1    g248(.A(new_n664), .ZN(new_n674));
  AND2_X1   g249(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n665), .A2(new_n669), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n676), .A2(new_n667), .ZN(new_n677));
  OAI211_X1 g252(.A(new_n671), .B(new_n673), .C1(new_n675), .C2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(new_n637), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT85), .B(G2100), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n678), .B(G2096), .ZN(new_n682));
  INV_X1    g257(.A(new_n680), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n681), .A2(new_n684), .ZN(G227));
  XNOR2_X1  g260(.A(G1991), .B(G1996), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G1971), .B(G1976), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT19), .ZN(new_n689));
  XOR2_X1   g264(.A(G1956), .B(G2474), .Z(new_n690));
  XOR2_X1   g265(.A(G1961), .B(G1966), .Z(new_n691));
  AND2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT20), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n690), .A2(new_n691), .ZN(new_n695));
  NOR3_X1   g270(.A1(new_n689), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n689), .B2(new_n695), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G1981), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G1986), .ZN(new_n700));
  INV_X1    g275(.A(G1981), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n698), .B(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G1986), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT86), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  AND3_X1   g282(.A1(new_n700), .A2(new_n704), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n707), .B1(new_n700), .B2(new_n704), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n687), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n700), .A2(new_n704), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(new_n706), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n700), .A2(new_n704), .A3(new_n707), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n712), .A2(new_n686), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n710), .A2(new_n714), .ZN(G229));
  NAND2_X1  g290(.A1(new_n481), .A2(G141), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n460), .A2(G105), .ZN(new_n717));
  NAND3_X1  g292(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT26), .ZN(new_n719));
  AOI211_X1 g294(.A(new_n717), .B(new_n719), .C1(G129), .C2(new_n483), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT93), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G29), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G29), .B2(G32), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT27), .B(G1996), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT94), .ZN(new_n727));
  NOR2_X1   g302(.A1(G5), .A2(G16), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G171), .B2(G16), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT96), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n730), .A2(G1961), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n730), .A2(G1961), .ZN(new_n732));
  NOR3_X1   g307(.A1(new_n727), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G29), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G35), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT97), .Z(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n488), .B2(G29), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT99), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G2090), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT89), .B(G16), .Z(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(G20), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT23), .Z(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G299), .B2(G16), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G1956), .ZN(new_n746));
  INV_X1    g321(.A(G16), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G4), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n618), .B2(new_n747), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G1348), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n749), .A2(G1348), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n750), .B(new_n751), .C1(new_n724), .C2(new_n725), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n734), .A2(G33), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n481), .A2(G139), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT25), .Z(new_n756));
  AOI22_X1  g331(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n757), .B2(new_n466), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n753), .B1(new_n759), .B2(new_n734), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n760), .A2(G2072), .ZN(new_n761));
  INV_X1    g336(.A(G1966), .ZN(new_n762));
  NOR2_X1   g337(.A1(G168), .A2(new_n747), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n747), .B2(G21), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n761), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n762), .B2(new_n764), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n636), .A2(G29), .B1(new_n760), .B2(G2072), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT31), .B(G11), .ZN(new_n768));
  INV_X1    g343(.A(G28), .ZN(new_n769));
  AOI21_X1  g344(.A(G29), .B1(new_n769), .B2(KEYINPUT30), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n770), .A2(KEYINPUT95), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(KEYINPUT30), .B2(new_n769), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n770), .A2(KEYINPUT95), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n768), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT24), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n734), .B1(new_n775), .B2(G34), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n775), .B2(G34), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G160), .B2(G29), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n774), .B1(new_n778), .B2(G2084), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n767), .B(new_n779), .C1(G2084), .C2(new_n778), .ZN(new_n780));
  INV_X1    g355(.A(new_n742), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n781), .A2(G19), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n556), .B2(new_n781), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(G1341), .Z(new_n784));
  NAND2_X1  g359(.A1(new_n734), .A2(G26), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT28), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n481), .A2(G140), .ZN(new_n787));
  OAI21_X1  g362(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n788));
  INV_X1    g363(.A(G116), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(G2105), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n790), .A2(KEYINPUT92), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(KEYINPUT92), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n791), .A2(new_n792), .B1(G128), .B2(new_n483), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n787), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n786), .B1(new_n794), .B2(G29), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G2067), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n734), .A2(G27), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G164), .B2(new_n734), .ZN(new_n798));
  INV_X1    g373(.A(G2078), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n784), .A2(new_n796), .A3(new_n800), .ZN(new_n801));
  NOR4_X1   g376(.A1(new_n752), .A2(new_n766), .A3(new_n780), .A4(new_n801), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n733), .A2(new_n741), .A3(new_n746), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n747), .A2(G6), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n585), .A2(new_n587), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n805), .B2(new_n747), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT32), .B(G1981), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n747), .A2(G23), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G288), .B2(G16), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT33), .B(G1976), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT90), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n810), .A2(new_n812), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n808), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n781), .A2(G22), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(G166), .B2(new_n781), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(G1971), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT91), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT34), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  NOR2_X1   g398(.A1(G25), .A2(G29), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n483), .A2(G119), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT87), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  OR2_X1    g402(.A1(G95), .A2(G2105), .ZN(new_n828));
  OAI211_X1 g403(.A(new_n828), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n829));
  INV_X1    g404(.A(G131), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n478), .A2(new_n480), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n827), .B(new_n829), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT88), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n824), .B1(new_n833), .B2(G29), .ZN(new_n834));
  XOR2_X1   g409(.A(KEYINPUT35), .B(G1991), .Z(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n834), .B(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n781), .A2(G24), .ZN(new_n838));
  INV_X1    g413(.A(G290), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n838), .B1(new_n839), .B2(new_n781), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(G1986), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n822), .A2(new_n823), .A3(new_n842), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n843), .A2(KEYINPUT36), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(KEYINPUT36), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n803), .B1(new_n844), .B2(new_n845), .ZN(G311));
  INV_X1    g421(.A(new_n803), .ZN(new_n847));
  INV_X1    g422(.A(new_n845), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n843), .A2(KEYINPUT36), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(G150));
  NAND2_X1  g425(.A1(G80), .A2(G543), .ZN(new_n851));
  INV_X1    g426(.A(G67), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n851), .B1(new_n504), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(G651), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n541), .A2(G93), .ZN(new_n855));
  INV_X1    g430(.A(G55), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n854), .B(new_n855), .C1(new_n856), .C2(new_n530), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(G860), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT37), .Z(new_n859));
  NOR2_X1   g434(.A1(new_n611), .A2(new_n619), .ZN(new_n860));
  XOR2_X1   g435(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT101), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n857), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n857), .A2(new_n863), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n864), .A2(new_n556), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n555), .A2(new_n857), .A3(new_n863), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n862), .B(new_n868), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n869), .A2(KEYINPUT39), .ZN(new_n870));
  INV_X1    g445(.A(G860), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(new_n869), .B2(KEYINPUT39), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n859), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT102), .ZN(G145));
  XNOR2_X1  g449(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(G160), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n635), .B(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(G162), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n832), .B(KEYINPUT88), .Z(new_n880));
  NAND2_X1  g455(.A1(new_n483), .A2(G130), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n466), .A2(G118), .ZN(new_n882));
  OAI21_X1  g457(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n883));
  INV_X1    g458(.A(G142), .ZN(new_n884));
  OAI221_X1 g459(.A(new_n881), .B1(new_n882), .B2(new_n883), .C1(new_n831), .C2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n641), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n880), .B(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT103), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n833), .A2(new_n886), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n833), .A2(new_n886), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT103), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n497), .A2(new_n499), .ZN(new_n894));
  AND2_X1   g469(.A1(KEYINPUT68), .A2(G114), .ZN(new_n895));
  NOR2_X1   g470(.A1(KEYINPUT68), .A2(G114), .ZN(new_n896));
  OAI21_X1  g471(.A(G2105), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n494), .ZN(new_n898));
  AOI22_X1  g473(.A1(G126), .A2(new_n483), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n894), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n794), .B(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n759), .A2(new_n721), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n759), .ZN(new_n905));
  OAI211_X1 g480(.A(new_n902), .B(new_n904), .C1(new_n722), .C2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n721), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT93), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT93), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n721), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n905), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n901), .B1(new_n911), .B2(new_n903), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n906), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n888), .A2(new_n893), .A3(new_n913), .A4(KEYINPUT104), .ZN(new_n914));
  INV_X1    g489(.A(new_n913), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n891), .A2(new_n892), .ZN(new_n916));
  AOI21_X1  g491(.A(KEYINPUT103), .B1(new_n889), .B2(new_n890), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n914), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n888), .A2(new_n893), .A3(new_n913), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT104), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n879), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(G37), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n879), .B1(new_n913), .B2(new_n891), .ZN(new_n925));
  INV_X1    g500(.A(new_n920), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n876), .B1(new_n923), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n927), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n878), .B(new_n488), .ZN(new_n930));
  INV_X1    g505(.A(new_n922), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n914), .A2(new_n918), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n929), .A2(new_n933), .A3(new_n875), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n928), .A2(new_n934), .ZN(G395));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT78), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n622), .B(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n938), .A2(new_n867), .A3(new_n866), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n623), .A2(new_n868), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT106), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n618), .A2(new_n574), .A3(new_n575), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n567), .A2(KEYINPUT74), .A3(new_n571), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT74), .B1(new_n567), .B2(new_n571), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n611), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n941), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n942), .A2(new_n945), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n947), .A2(KEYINPUT106), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n939), .B(new_n940), .C1(new_n946), .C2(new_n948), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n939), .A2(new_n940), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n942), .A2(new_n945), .A3(KEYINPUT41), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n945), .A2(new_n952), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n611), .B(KEYINPUT107), .C1(new_n943), .C2(new_n944), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n953), .A2(new_n942), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT41), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n951), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n949), .B1(new_n950), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(G166), .A2(G288), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(G303), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(G290), .A2(new_n805), .ZN(new_n963));
  NAND3_X1  g538(.A1(G305), .A2(new_n595), .A3(new_n596), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n959), .A2(new_n961), .A3(new_n963), .A4(new_n964), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n968), .A2(KEYINPUT42), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT108), .ZN(new_n970));
  AND4_X1   g545(.A1(new_n959), .A2(new_n961), .A3(new_n963), .A4(new_n964), .ZN(new_n971));
  AOI22_X1  g546(.A1(new_n959), .A2(new_n961), .B1(new_n963), .B2(new_n964), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n966), .A2(KEYINPUT108), .A3(new_n967), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n969), .B1(new_n975), .B2(KEYINPUT42), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n958), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n976), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n978), .B(new_n949), .C1(new_n950), .C2(new_n957), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(G868), .ZN(new_n981));
  INV_X1    g556(.A(G868), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n857), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n936), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n983), .ZN(new_n985));
  AOI211_X1 g560(.A(KEYINPUT109), .B(new_n985), .C1(new_n980), .C2(G868), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n984), .A2(new_n986), .ZN(G295));
  NAND2_X1  g562(.A1(new_n981), .A2(new_n983), .ZN(G331));
  INV_X1    g563(.A(KEYINPUT44), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n955), .A2(new_n956), .ZN(new_n990));
  INV_X1    g565(.A(new_n951), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT111), .ZN(new_n993));
  OAI211_X1 g568(.A(KEYINPUT110), .B(G168), .C1(new_n545), .C2(new_n546), .ZN(new_n994));
  OR2_X1    g569(.A1(new_n543), .A2(KEYINPUT72), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n521), .A2(new_n522), .ZN(new_n996));
  NAND2_X1  g571(.A1(G63), .A2(G651), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n519), .B1(new_n998), .B2(new_n507), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n999), .B(KEYINPUT110), .C1(new_n531), .C2(new_n530), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT110), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1001), .B1(new_n524), .B2(new_n532), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n995), .A2(new_n1000), .A3(new_n544), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n994), .A2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n1004), .B(new_n868), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n992), .A2(new_n993), .A3(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1004), .A2(new_n868), .ZN(new_n1007));
  AOI22_X1  g582(.A1(new_n994), .A2(new_n1003), .B1(new_n866), .B2(new_n867), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(KEYINPUT111), .B1(new_n957), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n947), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1006), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n975), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT43), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1006), .A2(new_n1010), .A3(new_n975), .A4(new_n1011), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1014), .A2(new_n1015), .A3(new_n924), .A4(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n948), .A2(new_n946), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n975), .B1(new_n1018), .B2(new_n1009), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n953), .A2(KEYINPUT41), .A3(new_n942), .A4(new_n954), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n947), .A2(new_n956), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1005), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(G37), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1016), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT43), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n989), .B1(new_n1017), .B2(new_n1025), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n1016), .A2(new_n1023), .A3(new_n1015), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1014), .A2(new_n924), .A3(new_n1016), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1027), .B1(new_n1028), .B2(KEYINPUT43), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1026), .B1(new_n989), .B2(new_n1029), .ZN(G397));
  INV_X1    g605(.A(KEYINPUT112), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT45), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1032), .B1(G164), .B2(G1384), .ZN(new_n1033));
  INV_X1    g608(.A(G125), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n476), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n471), .ZN(new_n1036));
  OAI21_X1  g611(.A(G2105), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n477), .A2(G137), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1037), .A2(G40), .A3(new_n461), .A4(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1031), .B1(new_n1033), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G1384), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n900), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(G40), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n469), .A2(new_n472), .A3(new_n1043), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1042), .A2(new_n1044), .A3(KEYINPUT112), .A4(new_n1032), .ZN(new_n1045));
  AND2_X1   g620(.A1(new_n1040), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G1996), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n1048), .B(KEYINPUT46), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n794), .A2(G2067), .ZN(new_n1050));
  INV_X1    g625(.A(G2067), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n787), .A2(new_n1051), .A3(new_n793), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1046), .B1(new_n721), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1049), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT47), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1049), .A2(KEYINPUT47), .A3(new_n1054), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1057), .A2(KEYINPUT127), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT127), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1046), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1053), .B1(G1996), .B2(new_n721), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n722), .A2(new_n1047), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n833), .A2(new_n835), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1064), .B1(KEYINPUT126), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1066), .B1(KEYINPUT126), .B2(new_n1065), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1061), .B1(new_n1067), .B2(new_n1052), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1046), .A2(new_n703), .A3(new_n839), .ZN(new_n1069));
  XOR2_X1   g644(.A(new_n1069), .B(KEYINPUT48), .Z(new_n1070));
  XNOR2_X1  g645(.A(new_n833), .B(new_n835), .ZN(new_n1071));
  OR2_X1    g646(.A1(new_n1071), .A2(new_n1064), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1070), .B1(new_n1046), .B2(new_n1072), .ZN(new_n1073));
  NOR4_X1   g648(.A1(new_n1059), .A2(new_n1060), .A3(new_n1068), .A4(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT114), .ZN(new_n1075));
  OAI21_X1  g650(.A(G1981), .B1(new_n585), .B2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1076), .A2(new_n805), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1076), .A2(new_n805), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1078), .A2(KEYINPUT49), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT49), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1079), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1081), .B1(new_n1082), .B2(new_n1077), .ZN(new_n1083));
  INV_X1    g658(.A(G8), .ZN(new_n1084));
  AOI21_X1  g659(.A(G1384), .B1(new_n894), .B2(new_n899), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1084), .B1(new_n1044), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1080), .A2(new_n1083), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n960), .A2(G1976), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(new_n1086), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT52), .ZN(new_n1090));
  INV_X1    g665(.A(G1976), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT52), .B1(G288), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1086), .A2(new_n1088), .A3(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1087), .A2(new_n1090), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT115), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1087), .A2(new_n1090), .A3(KEYINPUT115), .A4(new_n1093), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(G303), .A2(G8), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT55), .ZN(new_n1100));
  XNOR2_X1  g675(.A(new_n1099), .B(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1085), .A2(KEYINPUT45), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1033), .A2(new_n1102), .A3(KEYINPUT113), .ZN(new_n1103));
  OR3_X1    g678(.A1(new_n1085), .A2(KEYINPUT113), .A3(KEYINPUT45), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1039), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1105), .A2(G1971), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1039), .B1(new_n1042), .B2(KEYINPUT50), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT50), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1085), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1110), .A2(G2090), .ZN(new_n1111));
  OAI211_X1 g686(.A(G8), .B(new_n1101), .C1(new_n1106), .C2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(G8), .B1(new_n1106), .B2(new_n1111), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1101), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1033), .A2(new_n1044), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1102), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n762), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(G2084), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1107), .A2(new_n1119), .A3(new_n1109), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1121), .A2(G8), .A3(G168), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT63), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1098), .A2(new_n1112), .A3(new_n1115), .A4(new_n1124), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n1087), .A2(new_n1090), .A3(new_n1093), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1112), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1044), .B1(new_n1085), .B2(new_n1108), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT116), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1044), .B(KEYINPUT116), .C1(new_n1108), .C2(new_n1085), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1130), .A2(new_n1109), .A3(new_n1131), .ZN(new_n1132));
  OAI22_X1  g707(.A1(new_n1132), .A2(G2090), .B1(new_n1105), .B2(G1971), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1101), .B1(new_n1133), .B2(G8), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1127), .A2(new_n1134), .A3(new_n1122), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1125), .B1(new_n1135), .B2(KEYINPUT63), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT62), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1039), .B1(new_n1042), .B2(new_n1032), .ZN(new_n1139));
  AOI21_X1  g714(.A(G1966), .B1(new_n1139), .B2(new_n1102), .ZN(new_n1140));
  NOR3_X1   g715(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1141));
  NOR3_X1   g716(.A1(new_n1128), .A2(new_n1141), .A3(G2084), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1138), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1118), .A2(new_n1120), .A3(KEYINPUT123), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(G168), .A2(new_n1084), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1143), .A2(G168), .A3(new_n1144), .ZN(new_n1148));
  AND2_X1   g723(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1121), .A2(G8), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1146), .A2(KEYINPUT51), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1137), .B(new_n1147), .C1(new_n1150), .C2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(KEYINPUT53), .B1(new_n1105), .B2(new_n799), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT53), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1157), .A2(G2078), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(G1961), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1110), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(G171), .B1(new_n1155), .B2(new_n1162), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n1127), .A2(new_n1163), .A3(new_n1134), .ZN(new_n1164));
  AOI22_X1  g739(.A1(new_n1148), .A2(new_n1149), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1166));
  OAI21_X1  g741(.A(KEYINPUT62), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1154), .A2(new_n1164), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1112), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1087), .A2(new_n1091), .A3(new_n960), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1170), .B1(G1981), .B2(G305), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1169), .B1(new_n1086), .B2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1136), .A2(new_n1168), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(KEYINPUT57), .B1(new_n571), .B2(KEYINPUT117), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n572), .B(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1176));
  XNOR2_X1  g751(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(G2072), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1176), .A2(new_n1044), .A3(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(G1956), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1131), .A2(new_n1109), .ZN(new_n1181));
  OAI21_X1  g756(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1182));
  AOI21_X1  g757(.A(KEYINPUT116), .B1(new_n1182), .B2(new_n1044), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1180), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1175), .B1(new_n1179), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT119), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  AOI211_X1 g762(.A(KEYINPUT119), .B(new_n1175), .C1(new_n1179), .C2(new_n1184), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1179), .A2(new_n1184), .A3(new_n1175), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1189), .A2(KEYINPUT61), .ZN(new_n1190));
  NOR3_X1   g765(.A1(new_n1187), .A2(new_n1188), .A3(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT61), .ZN(new_n1192));
  AND3_X1   g767(.A1(new_n1179), .A2(new_n1184), .A3(new_n1175), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1192), .B1(new_n1193), .B2(new_n1185), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1044), .A2(new_n1085), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n1128), .A2(new_n1141), .ZN(new_n1196));
  OAI221_X1 g771(.A(new_n611), .B1(new_n1195), .B2(G2067), .C1(new_n1196), .C2(G1348), .ZN(new_n1197));
  AOI21_X1  g772(.A(G1348), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n1195), .A2(G2067), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n618), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1201));
  NOR2_X1   g776(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n611), .A2(KEYINPUT60), .ZN(new_n1203));
  AOI22_X1  g778(.A1(new_n1201), .A2(KEYINPUT60), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1194), .A2(new_n1204), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n1191), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g781(.A(KEYINPUT59), .ZN(new_n1207));
  NOR2_X1   g782(.A1(new_n1207), .A2(KEYINPUT121), .ZN(new_n1208));
  INV_X1    g783(.A(new_n1208), .ZN(new_n1209));
  NOR2_X1   g784(.A1(new_n1039), .A2(G1996), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1176), .A2(new_n1210), .ZN(new_n1211));
  XOR2_X1   g786(.A(KEYINPUT58), .B(G1341), .Z(new_n1212));
  NAND2_X1  g787(.A1(new_n1195), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1211), .A2(KEYINPUT120), .A3(new_n1213), .ZN(new_n1214));
  INV_X1    g789(.A(KEYINPUT120), .ZN(new_n1215));
  INV_X1    g790(.A(new_n1210), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1216), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1217));
  INV_X1    g792(.A(new_n1213), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n1215), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g794(.A1(new_n1214), .A2(new_n556), .A3(new_n1219), .ZN(new_n1220));
  INV_X1    g795(.A(KEYINPUT122), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1207), .A2(KEYINPUT121), .ZN(new_n1222));
  AND3_X1   g797(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  AOI21_X1  g798(.A(new_n1221), .B1(new_n1220), .B2(new_n1222), .ZN(new_n1224));
  OAI21_X1  g799(.A(new_n1209), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1220), .A2(new_n1222), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1226), .A2(KEYINPUT122), .ZN(new_n1227));
  NAND3_X1  g802(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1228));
  NAND3_X1  g803(.A1(new_n1227), .A2(new_n1208), .A3(new_n1228), .ZN(new_n1229));
  NAND3_X1  g804(.A1(new_n1206), .A2(new_n1225), .A3(new_n1229), .ZN(new_n1230));
  NOR2_X1   g805(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1231));
  NAND2_X1  g806(.A1(new_n1231), .A2(new_n1200), .ZN(new_n1232));
  NAND2_X1  g807(.A1(new_n1232), .A2(new_n1189), .ZN(new_n1233));
  NAND2_X1  g808(.A1(new_n1230), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1105), .A2(new_n799), .ZN(new_n1235));
  NAND2_X1  g810(.A1(new_n1235), .A2(new_n1157), .ZN(new_n1236));
  NAND4_X1  g811(.A1(new_n1236), .A2(G301), .A3(new_n1161), .A4(new_n1159), .ZN(new_n1237));
  INV_X1    g812(.A(KEYINPUT124), .ZN(new_n1238));
  NAND2_X1  g813(.A1(new_n1161), .A2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g814(.A1(new_n1110), .A2(KEYINPUT124), .A3(new_n1160), .ZN(new_n1240));
  NAND2_X1  g815(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  AND3_X1   g816(.A1(new_n1241), .A2(new_n1236), .A3(new_n1159), .ZN(new_n1242));
  OAI211_X1 g817(.A(KEYINPUT54), .B(new_n1237), .C1(new_n1242), .C2(G301), .ZN(new_n1243));
  NOR2_X1   g818(.A1(new_n1127), .A2(new_n1134), .ZN(new_n1244));
  OAI211_X1 g819(.A(new_n1243), .B(new_n1244), .C1(new_n1166), .C2(new_n1165), .ZN(new_n1245));
  AOI22_X1  g820(.A1(new_n1239), .A2(new_n1240), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1246));
  NAND4_X1  g821(.A1(new_n1246), .A2(KEYINPUT125), .A3(G301), .A4(new_n1236), .ZN(new_n1247));
  INV_X1    g822(.A(KEYINPUT54), .ZN(new_n1248));
  NAND2_X1  g823(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g824(.A(KEYINPUT125), .B1(new_n1242), .B2(G301), .ZN(new_n1250));
  AOI21_X1  g825(.A(new_n1249), .B1(new_n1250), .B2(new_n1163), .ZN(new_n1251));
  NOR2_X1   g826(.A1(new_n1245), .A2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g827(.A(new_n1173), .B1(new_n1234), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g828(.A(new_n1072), .ZN(new_n1254));
  XNOR2_X1  g829(.A(G290), .B(new_n703), .ZN(new_n1255));
  AOI21_X1  g830(.A(new_n1061), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  OAI21_X1  g831(.A(new_n1074), .B1(new_n1253), .B2(new_n1256), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g832(.A(G319), .B1(new_n660), .B2(new_n661), .ZN(new_n1259));
  AOI21_X1  g833(.A(new_n1259), .B1(new_n681), .B2(new_n684), .ZN(new_n1260));
  AND3_X1   g834(.A1(new_n710), .A2(new_n714), .A3(new_n1260), .ZN(new_n1261));
  OAI21_X1  g835(.A(new_n1261), .B1(new_n923), .B2(new_n927), .ZN(new_n1262));
  NOR2_X1   g836(.A1(new_n1262), .A2(new_n1029), .ZN(G308));
  NAND2_X1  g837(.A1(new_n929), .A2(new_n933), .ZN(new_n1264));
  AND2_X1   g838(.A1(new_n1028), .A2(KEYINPUT43), .ZN(new_n1265));
  OAI211_X1 g839(.A(new_n1264), .B(new_n1261), .C1(new_n1265), .C2(new_n1027), .ZN(G225));
endmodule


