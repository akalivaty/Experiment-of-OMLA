

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753;

  XNOR2_X1 U370 ( .A(n456), .B(n553), .ZN(n576) );
  NOR2_X1 U371 ( .A1(G953), .A2(G237), .ZN(n535) );
  XNOR2_X2 U372 ( .A(n437), .B(KEYINPUT19), .ZN(n593) );
  NOR2_X1 U373 ( .A1(n440), .A2(n438), .ZN(n627) );
  NOR2_X1 U374 ( .A1(n680), .A2(n679), .ZN(n462) );
  INV_X1 U375 ( .A(n693), .ZN(n596) );
  INV_X4 U376 ( .A(G143), .ZN(n460) );
  NOR2_X1 U377 ( .A1(n373), .A2(KEYINPUT2), .ZN(n668) );
  XNOR2_X1 U378 ( .A(n627), .B(n626), .ZN(n373) );
  NOR2_X1 U379 ( .A1(n584), .A2(n350), .ZN(n585) );
  XNOR2_X1 U380 ( .A(n622), .B(KEYINPUT32), .ZN(n753) );
  NAND2_X1 U381 ( .A1(n574), .A2(n556), .ZN(n657) );
  NAND2_X1 U382 ( .A1(n433), .A2(n450), .ZN(n449) );
  AND2_X2 U383 ( .A1(n376), .A2(n373), .ZN(n672) );
  XNOR2_X1 U384 ( .A(n668), .B(KEYINPUT85), .ZN(n669) );
  NAND2_X1 U385 ( .A1(n650), .A2(n753), .ZN(n445) );
  XNOR2_X1 U386 ( .A(n364), .B(KEYINPUT42), .ZN(n752) );
  XNOR2_X1 U387 ( .A(n453), .B(n358), .ZN(n374) );
  XNOR2_X1 U388 ( .A(n462), .B(n557), .ZN(n700) );
  NOR2_X1 U389 ( .A1(n424), .A2(n421), .ZN(n566) );
  INV_X1 U390 ( .A(n657), .ZN(n468) );
  XNOR2_X1 U391 ( .A(n578), .B(n382), .ZN(n677) );
  XNOR2_X1 U392 ( .A(n510), .B(n411), .ZN(n526) );
  XOR2_X2 U393 ( .A(G146), .B(G125), .Z(n501) );
  XNOR2_X1 U394 ( .A(G137), .B(G140), .ZN(n408) );
  XNOR2_X2 U395 ( .A(n467), .B(n355), .ZN(n558) );
  OR2_X2 U396 ( .A1(n711), .A2(G902), .ZN(n467) );
  XNOR2_X1 U397 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n626) );
  NAND2_X1 U398 ( .A1(n625), .A2(n439), .ZN(n438) );
  NAND2_X1 U399 ( .A1(n542), .A2(n543), .ZN(n560) );
  XNOR2_X1 U400 ( .A(n375), .B(n381), .ZN(n546) );
  XNOR2_X1 U401 ( .A(n488), .B(n730), .ZN(n375) );
  XNOR2_X1 U402 ( .A(n479), .B(n731), .ZN(n465) );
  NAND2_X1 U403 ( .A1(n559), .A2(KEYINPUT28), .ZN(n423) );
  AND2_X1 U404 ( .A1(n558), .A2(n427), .ZN(n422) );
  XNOR2_X1 U405 ( .A(n523), .B(n408), .ZN(n741) );
  INV_X1 U406 ( .A(n377), .ZN(n376) );
  XNOR2_X1 U407 ( .A(n432), .B(KEYINPUT39), .ZN(n469) );
  NAND2_X1 U408 ( .A1(n576), .A2(n555), .ZN(n432) );
  AND2_X1 U409 ( .A1(n451), .A2(n434), .ZN(n400) );
  INV_X1 U410 ( .A(n372), .ZN(n451) );
  XNOR2_X1 U411 ( .A(n466), .B(n360), .ZN(n586) );
  XNOR2_X1 U412 ( .A(n446), .B(n482), .ZN(n538) );
  XOR2_X1 U413 ( .A(KEYINPUT3), .B(G119), .Z(n482) );
  XNOR2_X1 U414 ( .A(n481), .B(n480), .ZN(n446) );
  INV_X1 U415 ( .A(KEYINPUT90), .ZN(n480) );
  XNOR2_X1 U416 ( .A(n558), .B(KEYINPUT1), .ZN(n690) );
  INV_X1 U417 ( .A(KEYINPUT111), .ZN(n393) );
  INV_X1 U418 ( .A(n690), .ZN(n606) );
  INV_X1 U419 ( .A(KEYINPUT34), .ZN(n389) );
  NAND2_X1 U420 ( .A1(n546), .A2(n547), .ZN(n407) );
  NAND2_X1 U421 ( .A1(n422), .A2(n423), .ZN(n421) );
  XNOR2_X1 U422 ( .A(n504), .B(n503), .ZN(n574) );
  XNOR2_X1 U423 ( .A(KEYINPUT13), .B(G475), .ZN(n503) );
  NAND2_X1 U424 ( .A1(n526), .A2(G221), .ZN(n410) );
  XNOR2_X1 U425 ( .A(n475), .B(KEYINPUT89), .ZN(n725) );
  NAND2_X1 U426 ( .A1(n672), .A2(KEYINPUT2), .ZN(n673) );
  AND2_X1 U427 ( .A1(n402), .A2(n401), .ZN(n397) );
  NAND2_X1 U428 ( .A1(G953), .A2(n434), .ZN(n401) );
  NAND2_X1 U429 ( .A1(n372), .A2(n348), .ZN(n402) );
  INV_X1 U430 ( .A(n452), .ZN(n450) );
  XNOR2_X1 U431 ( .A(KEYINPUT70), .B(G113), .ZN(n481) );
  XNOR2_X1 U432 ( .A(n430), .B(n501), .ZN(n484) );
  XNOR2_X1 U433 ( .A(n483), .B(n431), .ZN(n430) );
  INV_X1 U434 ( .A(KEYINPUT91), .ZN(n431) );
  NAND2_X1 U435 ( .A1(n740), .A2(G101), .ZN(n386) );
  XNOR2_X1 U436 ( .A(G116), .B(G137), .ZN(n531) );
  XOR2_X1 U437 ( .A(KEYINPUT97), .B(KEYINPUT5), .Z(n532) );
  XNOR2_X1 U438 ( .A(G131), .B(G134), .ZN(n739) );
  XOR2_X1 U439 ( .A(KEYINPUT101), .B(KEYINPUT12), .Z(n494) );
  XNOR2_X1 U440 ( .A(G143), .B(G104), .ZN(n496) );
  XOR2_X1 U441 ( .A(G140), .B(G131), .Z(n492) );
  XNOR2_X1 U442 ( .A(G113), .B(G122), .ZN(n491) );
  XNOR2_X1 U443 ( .A(n501), .B(KEYINPUT10), .ZN(n523) );
  XNOR2_X1 U444 ( .A(n408), .B(n354), .ZN(n405) );
  XNOR2_X1 U445 ( .A(n490), .B(n489), .ZN(n458) );
  INV_X1 U446 ( .A(KEYINPUT76), .ZN(n489) );
  XNOR2_X1 U447 ( .A(n739), .B(G146), .ZN(n536) );
  NAND2_X1 U448 ( .A1(n677), .A2(n676), .ZN(n680) );
  INV_X1 U449 ( .A(KEYINPUT38), .ZN(n382) );
  OR2_X1 U450 ( .A1(G902), .A2(G237), .ZN(n548) );
  XNOR2_X1 U451 ( .A(G902), .B(KEYINPUT15), .ZN(n547) );
  AND2_X1 U452 ( .A1(n391), .A2(n415), .ZN(n530) );
  NAND2_X1 U453 ( .A1(G234), .A2(G237), .ZN(n518) );
  XNOR2_X1 U454 ( .A(n476), .B(G110), .ZN(n731) );
  XNOR2_X1 U455 ( .A(G104), .B(KEYINPUT73), .ZN(n476) );
  XNOR2_X1 U456 ( .A(n447), .B(n538), .ZN(n730) );
  XNOR2_X1 U457 ( .A(n380), .B(n379), .ZN(n413) );
  XNOR2_X1 U458 ( .A(G119), .B(KEYINPUT71), .ZN(n380) );
  XNOR2_X1 U459 ( .A(KEYINPUT94), .B(KEYINPUT24), .ZN(n379) );
  INV_X1 U460 ( .A(KEYINPUT8), .ZN(n411) );
  XOR2_X1 U461 ( .A(KEYINPUT103), .B(KEYINPUT7), .Z(n506) );
  XNOR2_X1 U462 ( .A(G134), .B(KEYINPUT9), .ZN(n505) );
  XNOR2_X1 U463 ( .A(n385), .B(n384), .ZN(n508) );
  INV_X1 U464 ( .A(G122), .ZN(n384) );
  XNOR2_X1 U465 ( .A(G107), .B(G116), .ZN(n385) );
  XNOR2_X1 U466 ( .A(n488), .B(n457), .ZN(n711) );
  XNOR2_X1 U467 ( .A(n406), .B(n404), .ZN(n457) );
  XNOR2_X1 U468 ( .A(n458), .B(n731), .ZN(n406) );
  XNOR2_X1 U469 ( .A(n405), .B(n536), .ZN(n404) );
  NAND2_X1 U470 ( .A1(n371), .A2(n349), .ZN(n372) );
  AND2_X1 U471 ( .A1(n452), .A2(KEYINPUT2), .ZN(n370) );
  AND2_X1 U472 ( .A1(n471), .A2(KEYINPUT120), .ZN(n452) );
  AND2_X1 U473 ( .A1(n604), .A2(n415), .ZN(n454) );
  XOR2_X1 U474 ( .A(KEYINPUT6), .B(n693), .Z(n616) );
  XNOR2_X1 U475 ( .A(n487), .B(n486), .ZN(n628) );
  NAND2_X1 U476 ( .A1(n363), .A2(n361), .ZN(n429) );
  NAND2_X1 U477 ( .A1(n549), .A2(n383), .ZN(n550) );
  OR2_X1 U478 ( .A1(n700), .A2(n461), .ZN(n364) );
  INV_X1 U479 ( .A(n566), .ZN(n461) );
  INV_X1 U480 ( .A(n660), .ZN(n428) );
  NOR2_X1 U481 ( .A1(n392), .A2(n606), .ZN(n663) );
  XNOR2_X1 U482 ( .A(n615), .B(KEYINPUT35), .ZN(n751) );
  XNOR2_X1 U483 ( .A(n390), .B(n389), .ZN(n613) );
  NAND2_X1 U484 ( .A1(n419), .A2(n418), .ZN(n417) );
  INV_X1 U485 ( .A(n725), .ZN(n418) );
  XNOR2_X1 U486 ( .A(n420), .B(n359), .ZN(n419) );
  XNOR2_X1 U487 ( .A(n721), .B(n435), .ZN(n724) );
  AND2_X1 U488 ( .A1(n448), .A2(n348), .ZN(n396) );
  AND2_X1 U489 ( .A1(KEYINPUT53), .A2(n710), .ZN(n348) );
  OR2_X1 U490 ( .A1(n471), .A2(KEYINPUT120), .ZN(n349) );
  INV_X2 U491 ( .A(G953), .ZN(n710) );
  INV_X1 U492 ( .A(n687), .ZN(n415) );
  OR2_X1 U493 ( .A1(n654), .A2(n583), .ZN(n350) );
  XOR2_X1 U494 ( .A(n675), .B(KEYINPUT119), .Z(n351) );
  AND2_X1 U495 ( .A1(n749), .A2(n665), .ZN(n352) );
  AND2_X1 U496 ( .A1(n585), .A2(n587), .ZN(n353) );
  XOR2_X1 U497 ( .A(G107), .B(KEYINPUT93), .Z(n354) );
  XOR2_X1 U498 ( .A(KEYINPUT69), .B(G469), .Z(n355) );
  XOR2_X1 U499 ( .A(n529), .B(n528), .Z(n356) );
  NAND2_X1 U500 ( .A1(n673), .A2(n470), .ZN(n357) );
  XOR2_X1 U501 ( .A(KEYINPUT66), .B(KEYINPUT22), .Z(n358) );
  XNOR2_X1 U502 ( .A(n643), .B(KEYINPUT113), .ZN(n359) );
  INV_X1 U503 ( .A(KEYINPUT120), .ZN(n470) );
  XOR2_X1 U504 ( .A(KEYINPUT46), .B(KEYINPUT64), .Z(n360) );
  AND2_X1 U505 ( .A1(n632), .A2(G210), .ZN(n361) );
  INV_X1 U506 ( .A(KEYINPUT53), .ZN(n434) );
  AND2_X1 U507 ( .A1(n632), .A2(G472), .ZN(n362) );
  NAND2_X1 U508 ( .A1(n363), .A2(n633), .ZN(n637) );
  NAND2_X1 U509 ( .A1(n363), .A2(n362), .ZN(n420) );
  AND2_X2 U510 ( .A1(n363), .A2(n632), .ZN(n720) );
  XNOR2_X2 U511 ( .A(n672), .B(n459), .ZN(n363) );
  NAND2_X1 U512 ( .A1(n455), .A2(n752), .ZN(n466) );
  XNOR2_X2 U513 ( .A(n365), .B(KEYINPUT40), .ZN(n455) );
  NAND2_X1 U514 ( .A1(n469), .A2(n468), .ZN(n365) );
  XNOR2_X1 U515 ( .A(n366), .B(n464), .ZN(n463) );
  NAND2_X1 U516 ( .A1(n368), .A2(n367), .ZN(n366) );
  NAND2_X1 U517 ( .A1(n353), .A2(n586), .ZN(n367) );
  NAND2_X1 U518 ( .A1(n369), .A2(KEYINPUT88), .ZN(n368) );
  NAND2_X1 U519 ( .A1(n586), .A2(n585), .ZN(n369) );
  NAND2_X1 U520 ( .A1(n370), .A2(n672), .ZN(n371) );
  NAND2_X1 U521 ( .A1(n373), .A2(n710), .ZN(n729) );
  NAND2_X1 U522 ( .A1(n374), .A2(n606), .ZN(n624) );
  NAND2_X1 U523 ( .A1(n374), .A2(n621), .ZN(n622) );
  XNOR2_X2 U524 ( .A(n534), .B(KEYINPUT72), .ZN(n488) );
  AND2_X2 U525 ( .A1(n377), .A2(n459), .ZN(n667) );
  XNOR2_X1 U526 ( .A(n377), .B(n744), .ZN(n743) );
  NAND2_X2 U527 ( .A1(n463), .A2(n352), .ZN(n377) );
  NAND2_X1 U528 ( .A1(n378), .A2(n558), .ZN(n388) );
  NOR2_X2 U529 ( .A1(n623), .A2(n687), .ZN(n378) );
  NAND2_X1 U530 ( .A1(n690), .A2(n378), .ZN(n610) );
  NOR2_X1 U531 ( .A1(n690), .A2(n378), .ZN(n691) );
  XNOR2_X1 U532 ( .A(n485), .B(n465), .ZN(n381) );
  INV_X1 U533 ( .A(n578), .ZN(n383) );
  NAND2_X2 U534 ( .A1(n387), .A2(n386), .ZN(n534) );
  OR2_X2 U535 ( .A1(n740), .A2(G101), .ZN(n387) );
  XNOR2_X2 U536 ( .A(n388), .B(KEYINPUT96), .ZN(n597) );
  XNOR2_X1 U537 ( .A(n671), .B(KEYINPUT83), .ZN(n674) );
  NAND2_X1 U538 ( .A1(n605), .A2(n454), .ZN(n453) );
  NAND2_X1 U539 ( .A1(n612), .A2(n605), .ZN(n390) );
  BUF_X2 U540 ( .A(n623), .Z(n391) );
  OR2_X2 U541 ( .A1(n723), .A2(G902), .ZN(n416) );
  AND2_X1 U542 ( .A1(n399), .A2(n397), .ZN(n395) );
  XNOR2_X1 U543 ( .A(n564), .B(n563), .ZN(n392) );
  XNOR2_X1 U544 ( .A(n560), .B(n393), .ZN(n561) );
  XNOR2_X2 U545 ( .A(n509), .B(KEYINPUT4), .ZN(n740) );
  XNOR2_X2 U546 ( .A(n394), .B(n541), .ZN(n693) );
  NOR2_X1 U547 ( .A1(n642), .A2(G902), .ZN(n394) );
  XNOR2_X1 U548 ( .A(n417), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U549 ( .A1(n395), .A2(n398), .ZN(G75) );
  NAND2_X1 U550 ( .A1(n396), .A2(n449), .ZN(n398) );
  NAND2_X1 U551 ( .A1(n449), .A2(n448), .ZN(n403) );
  NAND2_X1 U552 ( .A1(n403), .A2(n400), .ZN(n399) );
  NOR2_X2 U553 ( .A1(n638), .A2(n725), .ZN(n641) );
  XNOR2_X2 U554 ( .A(n407), .B(n472), .ZN(n578) );
  XNOR2_X1 U555 ( .A(n508), .B(KEYINPUT16), .ZN(n447) );
  XNOR2_X1 U556 ( .A(n409), .B(n741), .ZN(n723) );
  XNOR2_X1 U557 ( .A(n412), .B(n410), .ZN(n409) );
  XNOR2_X1 U558 ( .A(n414), .B(n413), .ZN(n412) );
  XNOR2_X1 U559 ( .A(n525), .B(n524), .ZN(n414) );
  XNOR2_X2 U560 ( .A(n416), .B(n356), .ZN(n623) );
  NAND2_X1 U561 ( .A1(n566), .A2(n593), .ZN(n567) );
  NOR2_X1 U562 ( .A1(n559), .A2(n425), .ZN(n424) );
  NAND2_X1 U563 ( .A1(n596), .A2(n426), .ZN(n425) );
  INV_X1 U564 ( .A(KEYINPUT28), .ZN(n426) );
  NAND2_X1 U565 ( .A1(n693), .A2(KEYINPUT28), .ZN(n427) );
  NAND2_X1 U566 ( .A1(n469), .A2(n428), .ZN(n665) );
  XNOR2_X1 U567 ( .A(n429), .B(n628), .ZN(n629) );
  NOR2_X1 U568 ( .A1(n751), .A2(KEYINPUT44), .ZN(n443) );
  NAND2_X1 U569 ( .A1(n442), .A2(n441), .ZN(n440) );
  XNOR2_X1 U570 ( .A(n611), .B(KEYINPUT33), .ZN(n685) );
  INV_X1 U571 ( .A(n674), .ZN(n433) );
  XNOR2_X1 U572 ( .A(n723), .B(n722), .ZN(n435) );
  XNOR2_X1 U573 ( .A(n436), .B(n631), .ZN(G51) );
  NOR2_X2 U574 ( .A1(n629), .A2(n725), .ZN(n436) );
  NOR2_X1 U575 ( .A1(n561), .A2(n437), .ZN(n564) );
  NAND2_X1 U576 ( .A1(n578), .A2(n676), .ZN(n437) );
  NAND2_X1 U577 ( .A1(n751), .A2(KEYINPUT44), .ZN(n439) );
  NAND2_X1 U578 ( .A1(n445), .A2(KEYINPUT44), .ZN(n441) );
  NAND2_X1 U579 ( .A1(n444), .A2(n443), .ZN(n442) );
  INV_X1 U580 ( .A(n445), .ZN(n444) );
  NAND2_X1 U581 ( .A1(n674), .A2(n357), .ZN(n448) );
  XNOR2_X2 U582 ( .A(n595), .B(n594), .ZN(n605) );
  XNOR2_X1 U583 ( .A(n455), .B(G131), .ZN(G33) );
  NAND2_X1 U584 ( .A1(n552), .A2(n551), .ZN(n456) );
  INV_X1 U585 ( .A(KEYINPUT2), .ZN(n459) );
  XNOR2_X2 U586 ( .A(n460), .B(G128), .ZN(n509) );
  INV_X1 U587 ( .A(KEYINPUT48), .ZN(n464) );
  NOR2_X1 U588 ( .A1(n709), .A2(n351), .ZN(n471) );
  AND2_X1 U589 ( .A1(n548), .A2(G210), .ZN(n472) );
  AND2_X1 U590 ( .A1(n535), .A2(G210), .ZN(n473) );
  NAND2_X1 U591 ( .A1(n391), .A2(n693), .ZN(n474) );
  INV_X1 U592 ( .A(KEYINPUT86), .ZN(n666) );
  INV_X1 U593 ( .A(KEYINPUT11), .ZN(n495) );
  XNOR2_X1 U594 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U595 ( .A(n536), .B(n473), .ZN(n537) );
  INV_X1 U596 ( .A(KEYINPUT25), .ZN(n528) );
  INV_X1 U597 ( .A(KEYINPUT112), .ZN(n562) );
  XNOR2_X1 U598 ( .A(n562), .B(KEYINPUT36), .ZN(n563) );
  INV_X1 U599 ( .A(KEYINPUT60), .ZN(n639) );
  XNOR2_X1 U600 ( .A(n639), .B(KEYINPUT67), .ZN(n640) );
  INV_X1 U601 ( .A(G952), .ZN(n706) );
  NAND2_X1 U602 ( .A1(n706), .A2(G953), .ZN(n475) );
  XOR2_X1 U603 ( .A(KEYINPUT54), .B(KEYINPUT121), .Z(n487) );
  XOR2_X1 U604 ( .A(KEYINPUT78), .B(KEYINPUT17), .Z(n478) );
  XNOR2_X1 U605 ( .A(KEYINPUT92), .B(KEYINPUT77), .ZN(n477) );
  XNOR2_X1 U606 ( .A(n478), .B(n477), .ZN(n479) );
  NAND2_X1 U607 ( .A1(G224), .A2(n710), .ZN(n483) );
  XOR2_X1 U608 ( .A(n484), .B(KEYINPUT18), .Z(n485) );
  XNOR2_X1 U609 ( .A(n546), .B(KEYINPUT55), .ZN(n486) );
  INV_X1 U610 ( .A(n547), .ZN(n632) );
  NAND2_X1 U611 ( .A1(G227), .A2(n710), .ZN(n490) );
  XNOR2_X1 U612 ( .A(n492), .B(n491), .ZN(n500) );
  NAND2_X1 U613 ( .A1(n535), .A2(G214), .ZN(n493) );
  XNOR2_X1 U614 ( .A(n494), .B(n493), .ZN(n498) );
  XNOR2_X1 U615 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U616 ( .A(n500), .B(n499), .ZN(n502) );
  XNOR2_X1 U617 ( .A(n523), .B(n502), .ZN(n635) );
  NOR2_X1 U618 ( .A1(G902), .A2(n635), .ZN(n504) );
  XNOR2_X1 U619 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U620 ( .A(n508), .B(n507), .Z(n514) );
  XOR2_X1 U621 ( .A(n509), .B(KEYINPUT102), .Z(n512) );
  NAND2_X1 U622 ( .A1(G234), .A2(n710), .ZN(n510) );
  NAND2_X1 U623 ( .A1(G217), .A2(n526), .ZN(n511) );
  XNOR2_X1 U624 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U625 ( .A(n514), .B(n513), .ZN(n718) );
  NOR2_X1 U626 ( .A1(G902), .A2(n718), .ZN(n515) );
  XNOR2_X1 U627 ( .A(n515), .B(KEYINPUT104), .ZN(n516) );
  XNOR2_X1 U628 ( .A(n516), .B(G478), .ZN(n556) );
  NOR2_X1 U629 ( .A1(G953), .A2(n706), .ZN(n590) );
  NAND2_X1 U630 ( .A1(G953), .A2(G902), .ZN(n588) );
  NOR2_X1 U631 ( .A1(G900), .A2(n588), .ZN(n517) );
  NOR2_X1 U632 ( .A1(n590), .A2(n517), .ZN(n519) );
  XOR2_X1 U633 ( .A(KEYINPUT14), .B(n518), .Z(n705) );
  NOR2_X1 U634 ( .A1(n519), .A2(n705), .ZN(n551) );
  XOR2_X1 U635 ( .A(KEYINPUT95), .B(KEYINPUT21), .Z(n522) );
  NAND2_X1 U636 ( .A1(G234), .A2(n547), .ZN(n520) );
  XNOR2_X1 U637 ( .A(KEYINPUT20), .B(n520), .ZN(n527) );
  NAND2_X1 U638 ( .A1(n527), .A2(G221), .ZN(n521) );
  XNOR2_X1 U639 ( .A(n522), .B(n521), .ZN(n687) );
  XNOR2_X1 U640 ( .A(G128), .B(G110), .ZN(n524) );
  XOR2_X1 U641 ( .A(KEYINPUT75), .B(KEYINPUT23), .Z(n525) );
  NAND2_X1 U642 ( .A1(G217), .A2(n527), .ZN(n529) );
  NAND2_X1 U643 ( .A1(n551), .A2(n530), .ZN(n559) );
  NOR2_X1 U644 ( .A1(n657), .A2(n559), .ZN(n543) );
  XNOR2_X1 U645 ( .A(KEYINPUT98), .B(G472), .ZN(n541) );
  XNOR2_X1 U646 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U647 ( .A(n534), .B(n533), .ZN(n540) );
  XNOR2_X1 U648 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U649 ( .A(n540), .B(n539), .ZN(n642) );
  INV_X1 U650 ( .A(n616), .ZN(n542) );
  NOR2_X1 U651 ( .A1(n690), .A2(n560), .ZN(n544) );
  NAND2_X1 U652 ( .A1(G214), .A2(n548), .ZN(n676) );
  NAND2_X1 U653 ( .A1(n544), .A2(n676), .ZN(n545) );
  XNOR2_X1 U654 ( .A(n545), .B(KEYINPUT43), .ZN(n549) );
  XNOR2_X1 U655 ( .A(KEYINPUT108), .B(n550), .ZN(n749) );
  XNOR2_X1 U656 ( .A(n597), .B(KEYINPUT109), .ZN(n552) );
  INV_X1 U657 ( .A(KEYINPUT74), .ZN(n553) );
  NAND2_X1 U658 ( .A1(n676), .A2(n596), .ZN(n554) );
  XOR2_X1 U659 ( .A(KEYINPUT30), .B(n554), .Z(n575) );
  AND2_X1 U660 ( .A1(n677), .A2(n575), .ZN(n555) );
  OR2_X1 U661 ( .A1(n574), .A2(n556), .ZN(n660) );
  INV_X1 U662 ( .A(n556), .ZN(n573) );
  NOR2_X1 U663 ( .A1(n573), .A2(n574), .ZN(n604) );
  INV_X1 U664 ( .A(n604), .ZN(n679) );
  XNOR2_X1 U665 ( .A(KEYINPUT41), .B(KEYINPUT110), .ZN(n557) );
  NOR2_X1 U666 ( .A1(KEYINPUT47), .A2(KEYINPUT84), .ZN(n565) );
  NOR2_X1 U667 ( .A1(n663), .A2(n565), .ZN(n572) );
  XNOR2_X1 U668 ( .A(KEYINPUT82), .B(n567), .ZN(n655) );
  NAND2_X1 U669 ( .A1(KEYINPUT84), .A2(n655), .ZN(n569) );
  AND2_X1 U670 ( .A1(n657), .A2(n660), .ZN(n568) );
  XOR2_X1 U671 ( .A(KEYINPUT105), .B(n568), .Z(n681) );
  INV_X1 U672 ( .A(n681), .ZN(n602) );
  NAND2_X1 U673 ( .A1(n569), .A2(n602), .ZN(n570) );
  NAND2_X1 U674 ( .A1(n570), .A2(KEYINPUT47), .ZN(n571) );
  NAND2_X1 U675 ( .A1(n572), .A2(n571), .ZN(n584) );
  NAND2_X1 U676 ( .A1(n574), .A2(n573), .ZN(n609) );
  AND2_X1 U677 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U678 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U679 ( .A1(n609), .A2(n579), .ZN(n654) );
  INV_X1 U680 ( .A(KEYINPUT84), .ZN(n581) );
  NOR2_X1 U681 ( .A1(KEYINPUT47), .A2(n681), .ZN(n580) );
  NOR2_X1 U682 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U683 ( .A1(n655), .A2(n582), .ZN(n583) );
  INV_X1 U684 ( .A(KEYINPUT88), .ZN(n587) );
  NOR2_X1 U685 ( .A1(G898), .A2(n588), .ZN(n589) );
  NOR2_X1 U686 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U687 ( .A1(n705), .A2(n591), .ZN(n592) );
  NAND2_X1 U688 ( .A1(n593), .A2(n592), .ZN(n595) );
  XOR2_X1 U689 ( .A(KEYINPUT68), .B(KEYINPUT0), .Z(n594) );
  NOR2_X1 U690 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U691 ( .A1(n605), .A2(n598), .ZN(n646) );
  XOR2_X1 U692 ( .A(KEYINPUT31), .B(KEYINPUT100), .Z(n601) );
  OR2_X1 U693 ( .A1(n693), .A2(n610), .ZN(n599) );
  XNOR2_X1 U694 ( .A(n599), .B(KEYINPUT99), .ZN(n697) );
  NAND2_X1 U695 ( .A1(n697), .A2(n605), .ZN(n600) );
  XNOR2_X1 U696 ( .A(n601), .B(n600), .ZN(n661) );
  NAND2_X1 U697 ( .A1(n646), .A2(n661), .ZN(n603) );
  NAND2_X1 U698 ( .A1(n603), .A2(n602), .ZN(n608) );
  XNOR2_X1 U699 ( .A(n391), .B(KEYINPUT106), .ZN(n686) );
  NOR2_X1 U700 ( .A1(n686), .A2(n624), .ZN(n607) );
  NAND2_X1 U701 ( .A1(n616), .A2(n607), .ZN(n644) );
  AND2_X1 U702 ( .A1(n608), .A2(n644), .ZN(n625) );
  XNOR2_X1 U703 ( .A(n609), .B(KEYINPUT79), .ZN(n614) );
  NOR2_X1 U704 ( .A1(n610), .A2(n616), .ZN(n611) );
  INV_X1 U705 ( .A(n685), .ZN(n612) );
  NAND2_X1 U706 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U707 ( .A(n616), .B(KEYINPUT81), .ZN(n619) );
  AND2_X1 U708 ( .A1(n690), .A2(n686), .ZN(n617) );
  XNOR2_X1 U709 ( .A(n617), .B(KEYINPUT107), .ZN(n618) );
  NOR2_X1 U710 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U711 ( .A(KEYINPUT80), .B(n620), .ZN(n621) );
  OR2_X1 U712 ( .A1(n624), .A2(n474), .ZN(n650) );
  INV_X1 U713 ( .A(KEYINPUT87), .ZN(n630) );
  XNOR2_X1 U714 ( .A(n630), .B(KEYINPUT56), .ZN(n631) );
  AND2_X1 U715 ( .A1(n632), .A2(G475), .ZN(n633) );
  INV_X1 U716 ( .A(KEYINPUT59), .ZN(n634) );
  XNOR2_X1 U717 ( .A(n635), .B(n634), .ZN(n636) );
  XNOR2_X1 U718 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U719 ( .A(n641), .B(n640), .ZN(G60) );
  XNOR2_X1 U720 ( .A(n642), .B(KEYINPUT62), .ZN(n643) );
  XNOR2_X1 U721 ( .A(G101), .B(n644), .ZN(G3) );
  NOR2_X1 U722 ( .A1(n657), .A2(n646), .ZN(n645) );
  XOR2_X1 U723 ( .A(G104), .B(n645), .Z(G6) );
  NOR2_X1 U724 ( .A1(n660), .A2(n646), .ZN(n648) );
  XNOR2_X1 U725 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n647) );
  XNOR2_X1 U726 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U727 ( .A(G107), .B(n649), .ZN(G9) );
  XNOR2_X1 U728 ( .A(G110), .B(n650), .ZN(G12) );
  NOR2_X1 U729 ( .A1(n655), .A2(n660), .ZN(n652) );
  XNOR2_X1 U730 ( .A(KEYINPUT29), .B(KEYINPUT114), .ZN(n651) );
  XNOR2_X1 U731 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U732 ( .A(G128), .B(n653), .ZN(G30) );
  XOR2_X1 U733 ( .A(G143), .B(n654), .Z(G45) );
  NOR2_X1 U734 ( .A1(n655), .A2(n657), .ZN(n656) );
  XOR2_X1 U735 ( .A(G146), .B(n656), .Z(G48) );
  NOR2_X1 U736 ( .A1(n661), .A2(n657), .ZN(n659) );
  XNOR2_X1 U737 ( .A(G113), .B(KEYINPUT115), .ZN(n658) );
  XNOR2_X1 U738 ( .A(n659), .B(n658), .ZN(G15) );
  NOR2_X1 U739 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U740 ( .A(G116), .B(n662), .Z(G18) );
  XNOR2_X1 U741 ( .A(n663), .B(G125), .ZN(n664) );
  XNOR2_X1 U742 ( .A(n664), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U743 ( .A(G134), .B(n665), .ZN(G36) );
  XNOR2_X1 U744 ( .A(n667), .B(n666), .ZN(n670) );
  NAND2_X1 U745 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U746 ( .A1(n700), .A2(n685), .ZN(n675) );
  XNOR2_X1 U747 ( .A(KEYINPUT52), .B(KEYINPUT118), .ZN(n704) );
  NOR2_X1 U748 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U749 ( .A1(n679), .A2(n678), .ZN(n683) );
  NOR2_X1 U750 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U751 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U752 ( .A1(n685), .A2(n684), .ZN(n702) );
  XOR2_X1 U753 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n689) );
  NAND2_X1 U754 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U755 ( .A(n689), .B(n688), .ZN(n695) );
  XOR2_X1 U756 ( .A(KEYINPUT50), .B(n691), .Z(n692) );
  NAND2_X1 U757 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U758 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U759 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U760 ( .A(KEYINPUT51), .B(n698), .Z(n699) );
  NOR2_X1 U761 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U762 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U763 ( .A(n704), .B(n703), .ZN(n708) );
  OR2_X1 U764 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U765 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U766 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n713) );
  XNOR2_X1 U767 ( .A(n711), .B(KEYINPUT122), .ZN(n712) );
  XNOR2_X1 U768 ( .A(n713), .B(n712), .ZN(n715) );
  NAND2_X1 U769 ( .A1(n720), .A2(G469), .ZN(n714) );
  XNOR2_X1 U770 ( .A(n715), .B(n714), .ZN(n716) );
  NOR2_X1 U771 ( .A1(n725), .A2(n716), .ZN(G54) );
  NAND2_X1 U772 ( .A1(G478), .A2(n720), .ZN(n717) );
  XNOR2_X1 U773 ( .A(n718), .B(n717), .ZN(n719) );
  NOR2_X1 U774 ( .A1(n725), .A2(n719), .ZN(G63) );
  XOR2_X1 U775 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n722) );
  NAND2_X1 U776 ( .A1(n720), .A2(G217), .ZN(n721) );
  NOR2_X1 U777 ( .A1(n725), .A2(n724), .ZN(G66) );
  NAND2_X1 U778 ( .A1(G953), .A2(G224), .ZN(n726) );
  XNOR2_X1 U779 ( .A(KEYINPUT61), .B(n726), .ZN(n727) );
  NAND2_X1 U780 ( .A1(n727), .A2(G898), .ZN(n728) );
  NAND2_X1 U781 ( .A1(n729), .A2(n728), .ZN(n737) );
  XNOR2_X1 U782 ( .A(n730), .B(KEYINPUT126), .ZN(n733) );
  XNOR2_X1 U783 ( .A(G101), .B(n731), .ZN(n732) );
  XNOR2_X1 U784 ( .A(n733), .B(n732), .ZN(n735) );
  NOR2_X1 U785 ( .A1(G898), .A2(n710), .ZN(n734) );
  NOR2_X1 U786 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U787 ( .A(n737), .B(n736), .ZN(n738) );
  XOR2_X1 U788 ( .A(KEYINPUT125), .B(n738), .Z(G69) );
  XNOR2_X1 U789 ( .A(n740), .B(n739), .ZN(n742) );
  XOR2_X1 U790 ( .A(n742), .B(n741), .Z(n744) );
  NAND2_X1 U791 ( .A1(n743), .A2(n710), .ZN(n748) );
  XNOR2_X1 U792 ( .A(G227), .B(n744), .ZN(n745) );
  NAND2_X1 U793 ( .A1(n745), .A2(G900), .ZN(n746) );
  NAND2_X1 U794 ( .A1(n746), .A2(G953), .ZN(n747) );
  NAND2_X1 U795 ( .A1(n748), .A2(n747), .ZN(G72) );
  XNOR2_X1 U796 ( .A(G140), .B(n749), .ZN(n750) );
  XNOR2_X1 U797 ( .A(n750), .B(KEYINPUT116), .ZN(G42) );
  XOR2_X1 U798 ( .A(n751), .B(G122), .Z(G24) );
  XNOR2_X1 U799 ( .A(G137), .B(n752), .ZN(G39) );
  XNOR2_X1 U800 ( .A(G119), .B(n753), .ZN(G21) );
endmodule

