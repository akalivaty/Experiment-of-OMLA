

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757;

  AND2_X2 U364 ( .A1(n383), .A2(n382), .ZN(n393) );
  OR2_X2 U365 ( .A1(n632), .A2(G902), .ZN(n420) );
  XNOR2_X2 U366 ( .A(n408), .B(n407), .ZN(n505) );
  XNOR2_X2 U367 ( .A(KEYINPUT66), .B(G143), .ZN(n408) );
  OR2_X1 U368 ( .A1(n515), .A2(n514), .ZN(n517) );
  INV_X2 U369 ( .A(G953), .ZN(n742) );
  INV_X1 U370 ( .A(n524), .ZN(n341) );
  XNOR2_X1 U371 ( .A(n517), .B(n516), .ZN(n524) );
  XNOR2_X1 U372 ( .A(n677), .B(n421), .ZN(n588) );
  BUF_X1 U373 ( .A(n675), .Z(n362) );
  XNOR2_X1 U374 ( .A(n448), .B(n447), .ZN(n562) );
  XOR2_X1 U375 ( .A(G107), .B(G122), .Z(n497) );
  XNOR2_X1 U376 ( .A(KEYINPUT48), .B(KEYINPUT85), .ZN(n607) );
  NAND2_X1 U377 ( .A1(n365), .A2(n363), .ZN(n342) );
  NAND2_X1 U378 ( .A1(n365), .A2(n363), .ZN(n646) );
  XNOR2_X2 U379 ( .A(n356), .B(n574), .ZN(n750) );
  NOR2_X2 U380 ( .A1(n599), .A2(n573), .ZN(n356) );
  XNOR2_X1 U381 ( .A(KEYINPUT15), .B(G902), .ZN(n618) );
  NOR2_X1 U382 ( .A1(G902), .A2(G237), .ZN(n461) );
  NOR2_X1 U383 ( .A1(n679), .A2(n513), .ZN(n674) );
  INV_X1 U384 ( .A(KEYINPUT30), .ZN(n395) );
  XOR2_X1 U385 ( .A(G137), .B(KEYINPUT71), .Z(n409) );
  NAND2_X1 U386 ( .A1(n742), .A2(G224), .ZN(n376) );
  INV_X1 U387 ( .A(n618), .ZN(n367) );
  INV_X1 U388 ( .A(n712), .ZN(n359) );
  XNOR2_X1 U389 ( .A(n464), .B(n463), .ZN(n570) );
  XNOR2_X1 U390 ( .A(n562), .B(KEYINPUT1), .ZN(n675) );
  XNOR2_X1 U391 ( .A(n495), .B(n494), .ZN(n537) );
  XNOR2_X1 U392 ( .A(n493), .B(G475), .ZN(n494) );
  XNOR2_X1 U393 ( .A(n434), .B(n433), .ZN(n679) );
  NOR2_X1 U394 ( .A1(G953), .A2(G237), .ZN(n481) );
  XOR2_X1 U395 ( .A(G101), .B(G119), .Z(n413) );
  XNOR2_X1 U396 ( .A(n412), .B(n411), .ZN(n414) );
  INV_X1 U397 ( .A(KEYINPUT3), .ZN(n411) );
  XOR2_X1 U398 ( .A(G110), .B(G104), .Z(n450) );
  XNOR2_X1 U399 ( .A(n455), .B(n402), .ZN(n480) );
  XNOR2_X1 U400 ( .A(KEYINPUT10), .B(KEYINPUT70), .ZN(n402) );
  BUF_X1 U401 ( .A(n570), .Z(n612) );
  XNOR2_X1 U402 ( .A(n509), .B(n508), .ZN(n539) );
  INV_X1 U403 ( .A(G902), .ZN(n507) );
  INV_X1 U404 ( .A(n362), .ZN(n375) );
  NAND2_X1 U405 ( .A1(n343), .A2(n351), .ZN(n358) );
  AND2_X1 U406 ( .A1(n720), .A2(n742), .ZN(n361) );
  NAND2_X1 U407 ( .A1(G234), .A2(G237), .ZN(n469) );
  INV_X1 U408 ( .A(KEYINPUT76), .ZN(n390) );
  XNOR2_X1 U409 ( .A(G116), .B(G113), .ZN(n412) );
  XOR2_X1 U410 ( .A(G131), .B(G140), .Z(n479) );
  XNOR2_X1 U411 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U412 ( .A(G101), .B(G107), .ZN(n439) );
  XNOR2_X1 U413 ( .A(n354), .B(n353), .ZN(n695) );
  INV_X1 U414 ( .A(KEYINPUT109), .ZN(n353) );
  NAND2_X1 U415 ( .A1(n691), .A2(n690), .ZN(n354) );
  XNOR2_X1 U416 ( .A(n612), .B(n594), .ZN(n598) );
  XNOR2_X1 U417 ( .A(n397), .B(n396), .ZN(n586) );
  INV_X1 U418 ( .A(KEYINPUT72), .ZN(n396) );
  NOR2_X1 U419 ( .A1(n680), .A2(n399), .ZN(n398) );
  NOR2_X1 U420 ( .A1(n399), .A2(KEYINPUT76), .ZN(n392) );
  NOR2_X1 U421 ( .A1(n389), .A2(n388), .ZN(n387) );
  NOR2_X1 U422 ( .A1(n690), .A2(n395), .ZN(n388) );
  NOR2_X1 U423 ( .A1(n567), .A2(n390), .ZN(n389) );
  OR2_X1 U424 ( .A1(n569), .A2(n395), .ZN(n383) );
  AND2_X1 U425 ( .A1(n690), .A2(n395), .ZN(n394) );
  OR2_X1 U426 ( .A1(n570), .A2(n467), .ZN(n468) );
  AND2_X1 U427 ( .A1(n562), .A2(n674), .ZN(n568) );
  XNOR2_X1 U428 ( .A(G128), .B(G137), .ZN(n423) );
  XNOR2_X1 U429 ( .A(G119), .B(G110), .ZN(n426) );
  INV_X1 U430 ( .A(G128), .ZN(n407) );
  XNOR2_X1 U431 ( .A(G116), .B(KEYINPUT7), .ZN(n496) );
  XOR2_X1 U432 ( .A(KEYINPUT97), .B(KEYINPUT95), .Z(n483) );
  XNOR2_X1 U433 ( .A(G113), .B(G104), .ZN(n485) );
  XNOR2_X1 U434 ( .A(n357), .B(G122), .ZN(n488) );
  XNOR2_X1 U435 ( .A(n505), .B(n406), .ZN(n458) );
  XOR2_X1 U436 ( .A(KEYINPUT65), .B(KEYINPUT4), .Z(n406) );
  XNOR2_X1 U437 ( .A(n422), .B(G125), .ZN(n455) );
  NAND2_X1 U438 ( .A1(n379), .A2(n378), .ZN(n380) );
  NAND2_X1 U439 ( .A1(n376), .A2(KEYINPUT78), .ZN(n379) );
  NOR2_X1 U440 ( .A1(G953), .A2(KEYINPUT78), .ZN(n377) );
  XNOR2_X1 U441 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n454) );
  NAND2_X1 U442 ( .A1(n364), .A2(n344), .ZN(n363) );
  NAND2_X1 U443 ( .A1(n359), .A2(n350), .ZN(n365) );
  NAND2_X1 U444 ( .A1(n715), .A2(n714), .ZN(n712) );
  BUF_X1 U445 ( .A(n714), .Z(n728) );
  OR2_X1 U446 ( .A1(n524), .A2(n374), .ZN(n373) );
  NOR2_X1 U447 ( .A1(n372), .A2(n345), .ZN(n371) );
  NOR2_X1 U448 ( .A1(n375), .A2(n525), .ZN(n372) );
  BUF_X1 U449 ( .A(n515), .Z(n534) );
  XNOR2_X1 U450 ( .A(n381), .B(n418), .ZN(n632) );
  XNOR2_X1 U451 ( .A(n355), .B(n453), .ZN(n733) );
  XNOR2_X1 U452 ( .A(n403), .B(n400), .ZN(n724) );
  XNOR2_X1 U453 ( .A(n480), .B(n401), .ZN(n400) );
  XNOR2_X1 U454 ( .A(n429), .B(n348), .ZN(n403) );
  XNOR2_X1 U455 ( .A(n424), .B(n423), .ZN(n401) );
  BUF_X1 U456 ( .A(n342), .Z(n723) );
  NOR2_X1 U457 ( .A1(n609), .A2(n612), .ZN(n590) );
  BUF_X1 U458 ( .A(G143), .Z(n357) );
  INV_X1 U459 ( .A(n579), .ZN(n662) );
  NAND2_X1 U460 ( .A1(n369), .A2(n368), .ZN(n636) );
  NAND2_X1 U461 ( .A1(n370), .A2(KEYINPUT104), .ZN(n368) );
  AND2_X1 U462 ( .A1(n373), .A2(n371), .ZN(n369) );
  INV_X1 U463 ( .A(n341), .ZN(n370) );
  XNOR2_X1 U464 ( .A(KEYINPUT105), .B(n601), .ZN(n664) );
  XNOR2_X1 U465 ( .A(n545), .B(KEYINPUT102), .ZN(n756) );
  AND2_X1 U466 ( .A1(n719), .A2(n361), .ZN(n722) );
  NAND2_X1 U467 ( .A1(n713), .A2(KEYINPUT2), .ZN(n343) );
  AND2_X1 U468 ( .A1(n367), .A2(KEYINPUT2), .ZN(n344) );
  INV_X1 U469 ( .A(n567), .ZN(n399) );
  OR2_X1 U470 ( .A1(n569), .A2(n542), .ZN(n345) );
  AND2_X1 U471 ( .A1(n636), .A2(n639), .ZN(n346) );
  OR2_X1 U472 ( .A1(n712), .A2(KEYINPUT2), .ZN(n347) );
  XOR2_X1 U473 ( .A(n426), .B(n425), .Z(n348) );
  XOR2_X1 U474 ( .A(n632), .B(n631), .Z(n349) );
  AND2_X1 U475 ( .A1(n367), .A2(n366), .ZN(n350) );
  OR2_X1 U476 ( .A1(KEYINPUT2), .A2(KEYINPUT83), .ZN(n351) );
  INV_X1 U477 ( .A(KEYINPUT2), .ZN(n366) );
  XNOR2_X1 U478 ( .A(n352), .B(KEYINPUT42), .ZN(n597) );
  NOR2_X1 U479 ( .A1(n689), .A2(n596), .ZN(n352) );
  XNOR2_X1 U480 ( .A(n452), .B(n451), .ZN(n355) );
  NAND2_X1 U481 ( .A1(n358), .A2(n347), .ZN(n718) );
  XNOR2_X1 U482 ( .A(n750), .B(n575), .ZN(n576) );
  NOR2_X1 U483 ( .A1(n386), .A2(n385), .ZN(n384) );
  NAND2_X1 U484 ( .A1(n360), .A2(n634), .ZN(n635) );
  XNOR2_X1 U485 ( .A(n633), .B(n349), .ZN(n360) );
  NAND2_X1 U486 ( .A1(n646), .A2(G210), .ZN(n650) );
  NAND2_X1 U487 ( .A1(n714), .A2(n715), .ZN(n364) );
  XNOR2_X2 U488 ( .A(n556), .B(n555), .ZN(n714) );
  NAND2_X1 U489 ( .A1(n341), .A2(n375), .ZN(n544) );
  NAND2_X1 U490 ( .A1(n375), .A2(n525), .ZN(n374) );
  NAND2_X1 U491 ( .A1(n377), .A2(G224), .ZN(n378) );
  XNOR2_X1 U492 ( .A(n380), .B(n454), .ZN(n456) );
  XNOR2_X1 U493 ( .A(n381), .B(n444), .ZN(n619) );
  XNOR2_X2 U494 ( .A(n740), .B(G146), .ZN(n381) );
  NAND2_X1 U495 ( .A1(n569), .A2(n394), .ZN(n382) );
  XNOR2_X2 U496 ( .A(n526), .B(KEYINPUT103), .ZN(n569) );
  NAND2_X1 U497 ( .A1(n393), .A2(n384), .ZN(n599) );
  NOR2_X1 U498 ( .A1(n568), .A2(n390), .ZN(n385) );
  NAND2_X1 U499 ( .A1(n391), .A2(n387), .ZN(n386) );
  NAND2_X1 U500 ( .A1(n568), .A2(n392), .ZN(n391) );
  AND2_X1 U501 ( .A1(n569), .A2(n586), .ZN(n561) );
  NAND2_X1 U502 ( .A1(n679), .A2(n398), .ZN(n397) );
  XNOR2_X2 U503 ( .A(n468), .B(KEYINPUT19), .ZN(n564) );
  AND2_X1 U504 ( .A1(n628), .A2(n634), .ZN(G63) );
  AND2_X1 U505 ( .A1(n625), .A2(n634), .ZN(G54) );
  INV_X1 U506 ( .A(KEYINPUT82), .ZN(n575) );
  INV_X1 U507 ( .A(KEYINPUT74), .ZN(n584) );
  INV_X1 U508 ( .A(KEYINPUT90), .ZN(n438) );
  XNOR2_X1 U509 ( .A(n441), .B(n440), .ZN(n443) );
  INV_X1 U510 ( .A(KEYINPUT86), .ZN(n549) );
  XNOR2_X1 U511 ( .A(n485), .B(n484), .ZN(n486) );
  INV_X1 U512 ( .A(G469), .ZN(n445) );
  INV_X1 U513 ( .A(KEYINPUT24), .ZN(n425) );
  XNOR2_X1 U514 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U515 ( .A(n414), .B(n413), .ZN(n453) );
  INV_X1 U516 ( .A(n727), .ZN(n634) );
  INV_X1 U517 ( .A(n756), .ZN(n757) );
  XNOR2_X1 U518 ( .A(n409), .B(G134), .ZN(n410) );
  XNOR2_X2 U519 ( .A(n458), .B(n410), .ZN(n740) );
  XOR2_X1 U520 ( .A(G131), .B(KEYINPUT5), .Z(n416) );
  NAND2_X1 U521 ( .A1(n481), .A2(G210), .ZN(n415) );
  XNOR2_X1 U522 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U523 ( .A(n453), .B(n417), .ZN(n418) );
  INV_X1 U524 ( .A(G472), .ZN(n419) );
  XNOR2_X2 U525 ( .A(n420), .B(n419), .ZN(n526) );
  BUF_X2 U526 ( .A(n526), .Z(n677) );
  INV_X1 U527 ( .A(KEYINPUT6), .ZN(n421) );
  INV_X1 U528 ( .A(G146), .ZN(n422) );
  XOR2_X1 U529 ( .A(KEYINPUT23), .B(G140), .Z(n424) );
  NAND2_X1 U530 ( .A1(n742), .A2(G234), .ZN(n428) );
  XNOR2_X1 U531 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n427) );
  XNOR2_X1 U532 ( .A(n428), .B(n427), .ZN(n502) );
  NAND2_X1 U533 ( .A1(G221), .A2(n502), .ZN(n429) );
  NOR2_X1 U534 ( .A1(n724), .A2(G902), .ZN(n434) );
  NAND2_X1 U535 ( .A1(G234), .A2(n618), .ZN(n430) );
  XNOR2_X1 U536 ( .A(KEYINPUT20), .B(n430), .ZN(n435) );
  NAND2_X1 U537 ( .A1(G217), .A2(n435), .ZN(n432) );
  XNOR2_X1 U538 ( .A(KEYINPUT77), .B(KEYINPUT25), .ZN(n431) );
  XNOR2_X1 U539 ( .A(n432), .B(n431), .ZN(n433) );
  NAND2_X1 U540 ( .A1(G221), .A2(n435), .ZN(n436) );
  XNOR2_X1 U541 ( .A(n436), .B(KEYINPUT21), .ZN(n680) );
  INV_X1 U542 ( .A(KEYINPUT91), .ZN(n437) );
  XNOR2_X1 U543 ( .A(n680), .B(n437), .ZN(n513) );
  XOR2_X1 U544 ( .A(n479), .B(n450), .Z(n441) );
  NAND2_X1 U545 ( .A1(G227), .A2(n742), .ZN(n442) );
  XNOR2_X1 U546 ( .A(n443), .B(n442), .ZN(n444) );
  NOR2_X1 U547 ( .A1(n619), .A2(G902), .ZN(n448) );
  INV_X1 U548 ( .A(KEYINPUT73), .ZN(n446) );
  NAND2_X1 U549 ( .A1(n674), .A2(n675), .ZN(n533) );
  NOR2_X1 U550 ( .A1(n588), .A2(n533), .ZN(n449) );
  XNOR2_X1 U551 ( .A(KEYINPUT33), .B(n449), .ZN(n699) );
  XNOR2_X1 U552 ( .A(n497), .B(KEYINPUT16), .ZN(n452) );
  INV_X1 U553 ( .A(n450), .ZN(n451) );
  XNOR2_X1 U554 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U555 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U556 ( .A(n733), .B(n459), .ZN(n648) );
  NAND2_X1 U557 ( .A1(n648), .A2(n618), .ZN(n464) );
  INV_X1 U558 ( .A(KEYINPUT75), .ZN(n460) );
  XNOR2_X1 U559 ( .A(n461), .B(n460), .ZN(n466) );
  INV_X1 U560 ( .A(G210), .ZN(n462) );
  OR2_X1 U561 ( .A1(n466), .A2(n462), .ZN(n463) );
  INV_X1 U562 ( .A(G214), .ZN(n465) );
  OR2_X1 U563 ( .A1(n466), .A2(n465), .ZN(n690) );
  INV_X1 U564 ( .A(n690), .ZN(n467) );
  XNOR2_X1 U565 ( .A(n469), .B(KEYINPUT14), .ZN(n471) );
  NAND2_X1 U566 ( .A1(G952), .A2(n471), .ZN(n706) );
  NOR2_X1 U567 ( .A1(n706), .A2(G953), .ZN(n470) );
  XNOR2_X1 U568 ( .A(n470), .B(KEYINPUT89), .ZN(n560) );
  NAND2_X1 U569 ( .A1(G902), .A2(n471), .ZN(n557) );
  INV_X1 U570 ( .A(n557), .ZN(n472) );
  NOR2_X1 U571 ( .A1(G898), .A2(n742), .ZN(n735) );
  NAND2_X1 U572 ( .A1(n472), .A2(n735), .ZN(n473) );
  NAND2_X1 U573 ( .A1(n560), .A2(n473), .ZN(n474) );
  NAND2_X1 U574 ( .A1(n564), .A2(n474), .ZN(n477) );
  INV_X1 U575 ( .A(KEYINPUT87), .ZN(n475) );
  XNOR2_X1 U576 ( .A(n475), .B(KEYINPUT0), .ZN(n476) );
  XNOR2_X1 U577 ( .A(n477), .B(n476), .ZN(n515) );
  NOR2_X1 U578 ( .A1(n699), .A2(n534), .ZN(n478) );
  XNOR2_X1 U579 ( .A(n478), .B(KEYINPUT34), .ZN(n511) );
  XNOR2_X1 U580 ( .A(n480), .B(n479), .ZN(n739) );
  NAND2_X1 U581 ( .A1(G214), .A2(n481), .ZN(n482) );
  XNOR2_X1 U582 ( .A(n483), .B(n482), .ZN(n487) );
  INV_X1 U583 ( .A(KEYINPUT12), .ZN(n484) );
  XNOR2_X1 U584 ( .A(n487), .B(n486), .ZN(n491) );
  XOR2_X1 U585 ( .A(KEYINPUT11), .B(KEYINPUT96), .Z(n489) );
  XNOR2_X1 U586 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U587 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U588 ( .A(n739), .B(n492), .ZN(n641) );
  NOR2_X1 U589 ( .A1(n641), .A2(G902), .ZN(n495) );
  INV_X1 U590 ( .A(KEYINPUT13), .ZN(n493) );
  XNOR2_X1 U591 ( .A(n497), .B(n496), .ZN(n501) );
  XOR2_X1 U592 ( .A(KEYINPUT100), .B(KEYINPUT9), .Z(n499) );
  XNOR2_X1 U593 ( .A(G134), .B(KEYINPUT99), .ZN(n498) );
  XNOR2_X1 U594 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U595 ( .A(n501), .B(n500), .Z(n504) );
  NAND2_X1 U596 ( .A1(G217), .A2(n502), .ZN(n503) );
  XNOR2_X1 U597 ( .A(n504), .B(n503), .ZN(n506) );
  XNOR2_X1 U598 ( .A(n505), .B(n506), .ZN(n626) );
  NAND2_X1 U599 ( .A1(n626), .A2(n507), .ZN(n509) );
  INV_X1 U600 ( .A(G478), .ZN(n508) );
  NOR2_X1 U601 ( .A1(n537), .A2(n539), .ZN(n572) );
  XOR2_X1 U602 ( .A(n572), .B(KEYINPUT79), .Z(n510) );
  NAND2_X1 U603 ( .A1(n511), .A2(n510), .ZN(n512) );
  XNOR2_X2 U604 ( .A(n512), .B(KEYINPUT35), .ZN(n754) );
  INV_X1 U605 ( .A(n754), .ZN(n527) );
  NAND2_X1 U606 ( .A1(n537), .A2(n539), .ZN(n693) );
  OR2_X1 U607 ( .A1(n693), .A2(n513), .ZN(n514) );
  XNOR2_X1 U608 ( .A(KEYINPUT68), .B(KEYINPUT22), .ZN(n516) );
  NAND2_X1 U609 ( .A1(n362), .A2(n679), .ZN(n519) );
  INV_X1 U610 ( .A(n588), .ZN(n518) );
  NOR2_X1 U611 ( .A1(n519), .A2(n518), .ZN(n520) );
  NAND2_X1 U612 ( .A1(n341), .A2(n520), .ZN(n523) );
  INV_X1 U613 ( .A(KEYINPUT67), .ZN(n521) );
  XNOR2_X1 U614 ( .A(n521), .B(KEYINPUT32), .ZN(n522) );
  XNOR2_X1 U615 ( .A(n523), .B(n522), .ZN(n639) );
  INV_X1 U616 ( .A(KEYINPUT104), .ZN(n525) );
  INV_X1 U617 ( .A(n679), .ZN(n542) );
  NAND2_X1 U618 ( .A1(n527), .A2(n346), .ZN(n528) );
  NAND2_X1 U619 ( .A1(n528), .A2(KEYINPUT44), .ZN(n548) );
  INV_X1 U620 ( .A(n568), .ZN(n529) );
  NOR2_X1 U621 ( .A1(n534), .A2(n529), .ZN(n530) );
  XNOR2_X1 U622 ( .A(n530), .B(KEYINPUT92), .ZN(n531) );
  NAND2_X1 U623 ( .A1(n531), .A2(n677), .ZN(n532) );
  XNOR2_X1 U624 ( .A(n532), .B(KEYINPUT93), .ZN(n654) );
  OR2_X1 U625 ( .A1(n677), .A2(n533), .ZN(n673) );
  OR2_X1 U626 ( .A1(n534), .A2(n673), .ZN(n536) );
  XNOR2_X1 U627 ( .A(KEYINPUT94), .B(KEYINPUT31), .ZN(n535) );
  XNOR2_X1 U628 ( .A(n536), .B(n535), .ZN(n667) );
  NOR2_X1 U629 ( .A1(n654), .A2(n667), .ZN(n541) );
  XOR2_X1 U630 ( .A(n537), .B(KEYINPUT98), .Z(n538) );
  NAND2_X1 U631 ( .A1(n539), .A2(n538), .ZN(n601) );
  NOR2_X1 U632 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U633 ( .A(KEYINPUT101), .B(n540), .Z(n666) );
  INV_X1 U634 ( .A(n666), .ZN(n614) );
  NAND2_X1 U635 ( .A1(n601), .A2(n614), .ZN(n694) );
  XNOR2_X1 U636 ( .A(n694), .B(KEYINPUT81), .ZN(n580) );
  NOR2_X1 U637 ( .A1(n541), .A2(n580), .ZN(n546) );
  NAND2_X1 U638 ( .A1(n588), .A2(n542), .ZN(n543) );
  NOR2_X1 U639 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U640 ( .A1(n546), .A2(n756), .ZN(n547) );
  NAND2_X1 U641 ( .A1(n548), .A2(n547), .ZN(n550) );
  XNOR2_X1 U642 ( .A(n550), .B(n549), .ZN(n553) );
  NOR2_X1 U643 ( .A1(n754), .A2(KEYINPUT44), .ZN(n551) );
  NAND2_X1 U644 ( .A1(n551), .A2(n346), .ZN(n552) );
  NAND2_X1 U645 ( .A1(n553), .A2(n552), .ZN(n556) );
  XNOR2_X1 U646 ( .A(KEYINPUT84), .B(KEYINPUT45), .ZN(n554) );
  XNOR2_X1 U647 ( .A(n554), .B(KEYINPUT64), .ZN(n555) );
  NOR2_X1 U648 ( .A1(G900), .A2(n557), .ZN(n558) );
  NAND2_X1 U649 ( .A1(G953), .A2(n558), .ZN(n559) );
  NAND2_X1 U650 ( .A1(n560), .A2(n559), .ZN(n567) );
  XNOR2_X1 U651 ( .A(KEYINPUT28), .B(n561), .ZN(n563) );
  NAND2_X1 U652 ( .A1(n563), .A2(n562), .ZN(n596) );
  INV_X1 U653 ( .A(n596), .ZN(n565) );
  NAND2_X1 U654 ( .A1(n565), .A2(n564), .ZN(n579) );
  NAND2_X1 U655 ( .A1(n662), .A2(n694), .ZN(n566) );
  NAND2_X1 U656 ( .A1(n566), .A2(KEYINPUT47), .ZN(n577) );
  INV_X1 U657 ( .A(KEYINPUT107), .ZN(n574) );
  INV_X1 U658 ( .A(n612), .ZN(n571) );
  NAND2_X1 U659 ( .A1(n572), .A2(n571), .ZN(n573) );
  NAND2_X1 U660 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U661 ( .A(n578), .B(KEYINPUT80), .ZN(n583) );
  OR2_X1 U662 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U663 ( .A1(n581), .A2(KEYINPUT47), .ZN(n582) );
  NOR2_X2 U664 ( .A1(n583), .A2(n582), .ZN(n585) );
  XNOR2_X1 U665 ( .A(n585), .B(n584), .ZN(n593) );
  NAND2_X1 U666 ( .A1(n664), .A2(n586), .ZN(n587) );
  NOR2_X1 U667 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U668 ( .A1(n589), .A2(n690), .ZN(n609) );
  XNOR2_X1 U669 ( .A(n590), .B(KEYINPUT36), .ZN(n591) );
  NAND2_X1 U670 ( .A1(n591), .A2(n362), .ZN(n592) );
  XNOR2_X1 U671 ( .A(n592), .B(KEYINPUT111), .ZN(n752) );
  NOR2_X1 U672 ( .A1(n593), .A2(n752), .ZN(n606) );
  INV_X1 U673 ( .A(KEYINPUT38), .ZN(n594) );
  INV_X1 U674 ( .A(n598), .ZN(n691) );
  NOR2_X1 U675 ( .A1(n695), .A2(n693), .ZN(n595) );
  XNOR2_X1 U676 ( .A(n595), .B(KEYINPUT41), .ZN(n689) );
  XNOR2_X1 U677 ( .A(KEYINPUT110), .B(n597), .ZN(n755) );
  NOR2_X1 U678 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U679 ( .A(n600), .B(KEYINPUT39), .ZN(n615) );
  NOR2_X1 U680 ( .A1(n601), .A2(n615), .ZN(n603) );
  XNOR2_X1 U681 ( .A(KEYINPUT40), .B(KEYINPUT108), .ZN(n602) );
  XNOR2_X1 U682 ( .A(n603), .B(n602), .ZN(n751) );
  NOR2_X1 U683 ( .A1(n755), .A2(n751), .ZN(n604) );
  XNOR2_X1 U684 ( .A(n604), .B(KEYINPUT46), .ZN(n605) );
  NAND2_X1 U685 ( .A1(n606), .A2(n605), .ZN(n608) );
  XNOR2_X1 U686 ( .A(n608), .B(n607), .ZN(n617) );
  OR2_X1 U687 ( .A1(n362), .A2(n609), .ZN(n611) );
  XNOR2_X1 U688 ( .A(KEYINPUT106), .B(KEYINPUT43), .ZN(n610) );
  XNOR2_X1 U689 ( .A(n611), .B(n610), .ZN(n613) );
  NAND2_X1 U690 ( .A1(n613), .A2(n612), .ZN(n637) );
  OR2_X1 U691 ( .A1(n615), .A2(n614), .ZN(n669) );
  AND2_X1 U692 ( .A1(n637), .A2(n669), .ZN(n616) );
  AND2_X2 U693 ( .A1(n617), .A2(n616), .ZN(n715) );
  NAND2_X1 U694 ( .A1(n723), .A2(G469), .ZN(n623) );
  XOR2_X1 U695 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n621) );
  XNOR2_X1 U696 ( .A(n619), .B(KEYINPUT123), .ZN(n620) );
  XNOR2_X1 U697 ( .A(n621), .B(n620), .ZN(n622) );
  XNOR2_X1 U698 ( .A(n623), .B(n622), .ZN(n625) );
  INV_X1 U699 ( .A(G952), .ZN(n624) );
  AND2_X1 U700 ( .A1(n624), .A2(G953), .ZN(n727) );
  NAND2_X1 U701 ( .A1(n723), .A2(G478), .ZN(n627) );
  XNOR2_X1 U702 ( .A(n627), .B(n626), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n342), .A2(G472), .ZN(n633) );
  XOR2_X1 U704 ( .A(KEYINPUT88), .B(KEYINPUT113), .Z(n630) );
  XNOR2_X1 U705 ( .A(KEYINPUT62), .B(KEYINPUT112), .ZN(n629) );
  XNOR2_X1 U706 ( .A(n630), .B(n629), .ZN(n631) );
  XNOR2_X1 U707 ( .A(n635), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U708 ( .A(n636), .B(G110), .ZN(G12) );
  XNOR2_X1 U709 ( .A(n637), .B(G140), .ZN(G42) );
  XOR2_X1 U710 ( .A(G119), .B(KEYINPUT127), .Z(n638) );
  XNOR2_X1 U711 ( .A(n639), .B(n638), .ZN(G21) );
  NAND2_X1 U712 ( .A1(n646), .A2(G475), .ZN(n643) );
  XOR2_X1 U713 ( .A(KEYINPUT124), .B(KEYINPUT59), .Z(n640) );
  XNOR2_X1 U714 ( .A(n641), .B(n640), .ZN(n642) );
  XNOR2_X1 U715 ( .A(n643), .B(n642), .ZN(n644) );
  NOR2_X2 U716 ( .A1(n644), .A2(n727), .ZN(n645) );
  XNOR2_X1 U717 ( .A(n645), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U718 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n647) );
  XNOR2_X1 U719 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U720 ( .A(n650), .B(n649), .ZN(n651) );
  NOR2_X2 U721 ( .A1(n651), .A2(n727), .ZN(n652) );
  XNOR2_X1 U722 ( .A(n652), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U723 ( .A1(n654), .A2(n664), .ZN(n653) );
  XNOR2_X1 U724 ( .A(n653), .B(G104), .ZN(G6) );
  XNOR2_X1 U725 ( .A(KEYINPUT26), .B(KEYINPUT114), .ZN(n658) );
  XOR2_X1 U726 ( .A(G107), .B(KEYINPUT27), .Z(n656) );
  NAND2_X1 U727 ( .A1(n654), .A2(n666), .ZN(n655) );
  XNOR2_X1 U728 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U729 ( .A(n658), .B(n657), .ZN(G9) );
  XOR2_X1 U730 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n660) );
  NAND2_X1 U731 ( .A1(n662), .A2(n666), .ZN(n659) );
  XNOR2_X1 U732 ( .A(n660), .B(n659), .ZN(n661) );
  XOR2_X1 U733 ( .A(G128), .B(n661), .Z(G30) );
  NAND2_X1 U734 ( .A1(n662), .A2(n664), .ZN(n663) );
  XNOR2_X1 U735 ( .A(n663), .B(G146), .ZN(G48) );
  NAND2_X1 U736 ( .A1(n667), .A2(n664), .ZN(n665) );
  XNOR2_X1 U737 ( .A(n665), .B(G113), .ZN(G15) );
  NAND2_X1 U738 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U739 ( .A(n668), .B(G116), .ZN(G18) );
  INV_X1 U740 ( .A(n669), .ZN(n670) );
  XOR2_X1 U741 ( .A(G134), .B(n670), .Z(n671) );
  XNOR2_X1 U742 ( .A(KEYINPUT116), .B(n671), .ZN(G36) );
  NOR2_X1 U743 ( .A1(n689), .A2(n699), .ZN(n672) );
  XOR2_X1 U744 ( .A(KEYINPUT120), .B(n672), .Z(n709) );
  INV_X1 U745 ( .A(n673), .ZN(n686) );
  OR2_X1 U746 ( .A1(n362), .A2(n674), .ZN(n676) );
  XNOR2_X1 U747 ( .A(n676), .B(KEYINPUT50), .ZN(n678) );
  NAND2_X1 U748 ( .A1(n678), .A2(n677), .ZN(n683) );
  NAND2_X1 U749 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U750 ( .A(KEYINPUT49), .B(n681), .ZN(n682) );
  NOR2_X1 U751 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U752 ( .A(KEYINPUT117), .B(n684), .Z(n685) );
  NOR2_X1 U753 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U754 ( .A(KEYINPUT51), .B(n687), .Z(n688) );
  NOR2_X1 U755 ( .A1(n689), .A2(n688), .ZN(n703) );
  NOR2_X1 U756 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U757 ( .A1(n693), .A2(n692), .ZN(n698) );
  INV_X1 U758 ( .A(n694), .ZN(n696) );
  NOR2_X1 U759 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U760 ( .A1(n698), .A2(n697), .ZN(n700) );
  NOR2_X1 U761 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U762 ( .A(n701), .B(KEYINPUT118), .ZN(n702) );
  NOR2_X1 U763 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U764 ( .A(n704), .B(KEYINPUT52), .ZN(n705) );
  NOR2_X1 U765 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U766 ( .A(KEYINPUT119), .B(n707), .ZN(n708) );
  NAND2_X1 U767 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U768 ( .A(n710), .B(KEYINPUT121), .ZN(n720) );
  INV_X1 U769 ( .A(KEYINPUT83), .ZN(n711) );
  NAND2_X1 U770 ( .A1(n712), .A2(n711), .ZN(n713) );
  INV_X1 U771 ( .A(n715), .ZN(n738) );
  NAND2_X1 U772 ( .A1(n728), .A2(n738), .ZN(n716) );
  NAND2_X1 U773 ( .A1(n716), .A2(KEYINPUT83), .ZN(n717) );
  NAND2_X1 U774 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U775 ( .A(KEYINPUT53), .B(KEYINPUT122), .ZN(n721) );
  XNOR2_X1 U776 ( .A(n722), .B(n721), .ZN(G75) );
  NAND2_X1 U777 ( .A1(n723), .A2(G217), .ZN(n725) );
  XNOR2_X1 U778 ( .A(n725), .B(n724), .ZN(n726) );
  NOR2_X1 U779 ( .A1(n727), .A2(n726), .ZN(G66) );
  NAND2_X1 U780 ( .A1(n728), .A2(n742), .ZN(n732) );
  NAND2_X1 U781 ( .A1(G953), .A2(G224), .ZN(n729) );
  XNOR2_X1 U782 ( .A(KEYINPUT61), .B(n729), .ZN(n730) );
  NAND2_X1 U783 ( .A1(n730), .A2(G898), .ZN(n731) );
  NAND2_X1 U784 ( .A1(n732), .A2(n731), .ZN(n737) );
  XNOR2_X1 U785 ( .A(KEYINPUT125), .B(n733), .ZN(n734) );
  NOR2_X1 U786 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U787 ( .A(n737), .B(n736), .ZN(G69) );
  INV_X1 U788 ( .A(n738), .ZN(n741) );
  XNOR2_X1 U789 ( .A(n740), .B(n739), .ZN(n744) );
  XOR2_X1 U790 ( .A(n741), .B(n744), .Z(n743) );
  NAND2_X1 U791 ( .A1(n743), .A2(n742), .ZN(n748) );
  XNOR2_X1 U792 ( .A(G227), .B(n744), .ZN(n745) );
  NAND2_X1 U793 ( .A1(n745), .A2(G900), .ZN(n746) );
  NAND2_X1 U794 ( .A1(n746), .A2(G953), .ZN(n747) );
  NAND2_X1 U795 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U796 ( .A(KEYINPUT126), .B(n749), .ZN(G72) );
  XOR2_X1 U797 ( .A(n750), .B(n357), .Z(G45) );
  XOR2_X1 U798 ( .A(G131), .B(n751), .Z(G33) );
  XNOR2_X1 U799 ( .A(n752), .B(G125), .ZN(n753) );
  XNOR2_X1 U800 ( .A(n753), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U801 ( .A(n754), .B(G122), .Z(G24) );
  XOR2_X1 U802 ( .A(G137), .B(n755), .Z(G39) );
  XNOR2_X1 U803 ( .A(G101), .B(n757), .ZN(G3) );
endmodule

