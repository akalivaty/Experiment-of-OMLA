//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 1 0 1 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 0 0 0 0 1 1 1 0 1 0 0 0 0 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:02 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n537, new_n539, new_n540, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n559,
    new_n560, new_n561, new_n562, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n597, new_n598, new_n601, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1141, new_n1142,
    new_n1143, new_n1144;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT66), .Z(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(new_n451), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n456), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(new_n452), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  OR2_X1    g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n469), .A2(G137), .B1(G101), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n466), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  NAND2_X1  g049(.A1(new_n469), .A2(G136), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n476), .B1(new_n467), .B2(new_n468), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  MUX2_X1   g053(.A(G100), .B(G112), .S(G2105), .Z(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2104), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n475), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  AND2_X1   g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NOR2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  OAI211_X1 g059(.A(G138), .B(new_n476), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT4), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n462), .A2(new_n487), .A3(G138), .A4(new_n476), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(G114), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G102), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(G2105), .ZN(new_n492));
  AOI22_X1  g067(.A1(new_n477), .A2(G126), .B1(G2104), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G164));
  NAND2_X1  g070(.A1(KEYINPUT67), .A2(G543), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT5), .ZN(new_n497));
  XNOR2_X1  g072(.A(new_n496), .B(new_n497), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n498), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n499));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g076(.A(KEYINPUT6), .B(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G88), .ZN(new_n504));
  INV_X1    g079(.A(G50), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n502), .A2(G543), .ZN(new_n506));
  OAI22_X1  g081(.A1(new_n503), .A2(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n501), .A2(new_n507), .ZN(G166));
  INV_X1    g083(.A(new_n503), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n509), .A2(G89), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n498), .A2(G63), .A3(G651), .ZN(new_n511));
  NAND3_X1  g086(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n512));
  XNOR2_X1  g087(.A(new_n512), .B(KEYINPUT7), .ZN(new_n513));
  INV_X1    g088(.A(G51), .ZN(new_n514));
  OAI211_X1 g089(.A(new_n511), .B(new_n513), .C1(new_n514), .C2(new_n506), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n510), .A2(new_n515), .ZN(G168));
  AOI22_X1  g091(.A1(new_n498), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n517), .A2(new_n500), .ZN(new_n518));
  INV_X1    g093(.A(G90), .ZN(new_n519));
  INV_X1    g094(.A(G52), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n503), .A2(new_n519), .B1(new_n520), .B2(new_n506), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n518), .A2(new_n521), .ZN(G171));
  INV_X1    g097(.A(new_n506), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT68), .B(G43), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G81), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n526), .B2(new_n503), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(KEYINPUT69), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT69), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n525), .B(new_n529), .C1(new_n526), .C2(new_n503), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n498), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n532), .A2(new_n500), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G860), .ZN(G153));
  AND3_X1   g111(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G36), .ZN(G176));
  NAND2_X1  g113(.A1(G1), .A2(G3), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT8), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n537), .A2(new_n540), .ZN(G188));
  NAND2_X1  g116(.A1(G78), .A2(G543), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n496), .B(KEYINPUT5), .ZN(new_n543));
  INV_X1    g118(.A(G65), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G651), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(KEYINPUT70), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(KEYINPUT70), .ZN(new_n548));
  INV_X1    g123(.A(G53), .ZN(new_n549));
  OR3_X1    g124(.A1(new_n506), .A2(KEYINPUT9), .A3(new_n549), .ZN(new_n550));
  OAI21_X1  g125(.A(KEYINPUT9), .B1(new_n506), .B2(new_n549), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n550), .A2(new_n551), .B1(new_n509), .B2(G91), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n547), .A2(new_n548), .A3(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT71), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g130(.A1(new_n547), .A2(KEYINPUT71), .A3(new_n552), .A4(new_n548), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(G299));
  INV_X1    g133(.A(KEYINPUT72), .ZN(new_n559));
  NAND2_X1  g134(.A1(G171), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT72), .B1(new_n518), .B2(new_n521), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(G301));
  INV_X1    g138(.A(G168), .ZN(G286));
  INV_X1    g139(.A(G166), .ZN(G303));
  NAND2_X1  g140(.A1(new_n509), .A2(G87), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n498), .B2(G74), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n523), .A2(G49), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G288));
  NAND2_X1  g144(.A1(new_n523), .A2(G48), .ZN(new_n570));
  INV_X1    g145(.A(G86), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n571), .B2(new_n503), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n498), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n573), .A2(new_n500), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G305));
  AOI22_X1  g151(.A1(new_n498), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n577), .A2(new_n500), .ZN(new_n578));
  INV_X1    g153(.A(G85), .ZN(new_n579));
  INV_X1    g154(.A(G47), .ZN(new_n580));
  OAI22_X1  g155(.A1(new_n503), .A2(new_n579), .B1(new_n580), .B2(new_n506), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(G301), .A2(G868), .ZN(new_n584));
  AND3_X1   g159(.A1(new_n498), .A2(G92), .A3(new_n502), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n585), .B(KEYINPUT10), .ZN(new_n586));
  XOR2_X1   g161(.A(new_n506), .B(KEYINPUT73), .Z(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G54), .ZN(new_n588));
  AND2_X1   g163(.A1(new_n498), .A2(G66), .ZN(new_n589));
  NAND2_X1  g164(.A1(G79), .A2(G543), .ZN(new_n590));
  XOR2_X1   g165(.A(new_n590), .B(KEYINPUT74), .Z(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n586), .A2(new_n588), .A3(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n584), .B1(G868), .B2(new_n594), .ZN(G284));
  OAI21_X1  g170(.A(new_n584), .B1(G868), .B2(new_n594), .ZN(G321));
  NAND2_X1  g171(.A1(G286), .A2(G868), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n557), .B(KEYINPUT75), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(G868), .ZN(G297));
  OAI21_X1  g174(.A(new_n597), .B1(new_n598), .B2(G868), .ZN(G280));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n594), .B1(new_n601), .B2(G860), .ZN(G148));
  NOR2_X1   g177(.A1(new_n534), .A2(G868), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n593), .A2(G559), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n603), .B1(G868), .B2(new_n604), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g181(.A1(new_n469), .A2(G2104), .ZN(new_n607));
  XOR2_X1   g182(.A(new_n607), .B(KEYINPUT12), .Z(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(KEYINPUT13), .Z(new_n609));
  INV_X1    g184(.A(G2100), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n609), .A2(new_n610), .ZN(new_n612));
  MUX2_X1   g187(.A(G99), .B(G111), .S(G2105), .Z(new_n613));
  AOI22_X1  g188(.A1(G123), .A2(new_n477), .B1(new_n613), .B2(G2104), .ZN(new_n614));
  INV_X1    g189(.A(G135), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n462), .A2(new_n476), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(G2096), .Z(new_n618));
  NAND3_X1  g193(.A1(new_n611), .A2(new_n612), .A3(new_n618), .ZN(G156));
  XNOR2_X1  g194(.A(KEYINPUT15), .B(G2435), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2438), .ZN(new_n621));
  XNOR2_X1  g196(.A(G2427), .B(G2430), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(KEYINPUT14), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT76), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(new_n621), .B2(new_n622), .ZN(new_n626));
  XOR2_X1   g201(.A(G2451), .B(G2454), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT16), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n626), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(G2443), .B(G2446), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(G1341), .B(G1348), .ZN(new_n632));
  AND2_X1   g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(G14), .B1(new_n631), .B2(new_n632), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n633), .A2(new_n634), .ZN(G401));
  XNOR2_X1  g210(.A(G2072), .B(G2078), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT77), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT17), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2067), .B(G2678), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2084), .B(G2090), .ZN(new_n640));
  NOR3_X1   g215(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n640), .B1(new_n637), .B2(new_n639), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(new_n638), .B2(new_n639), .ZN(new_n643));
  INV_X1    g218(.A(new_n639), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n644), .A2(new_n640), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n637), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT18), .ZN(new_n647));
  NOR3_X1   g222(.A1(new_n641), .A2(new_n643), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2096), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2100), .ZN(G227));
  XOR2_X1   g225(.A(G1971), .B(G1976), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT19), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1956), .B(G2474), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1961), .B(G1966), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT20), .ZN(new_n657));
  AND2_X1   g232(.A1(new_n653), .A2(new_n654), .ZN(new_n658));
  NOR3_X1   g233(.A1(new_n652), .A2(new_n655), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n659), .B1(new_n652), .B2(new_n658), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT78), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n661), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT79), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1991), .B(G1996), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1981), .B(G1986), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n665), .B(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(G229));
  NOR2_X1   g245(.A1(G6), .A2(G16), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n671), .B1(new_n575), .B2(G16), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT82), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT32), .B(G1981), .Z(new_n674));
  OR2_X1    g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n673), .A2(new_n674), .ZN(new_n676));
  NOR2_X1   g251(.A1(G16), .A2(G23), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT83), .Z(new_n678));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n678), .B1(G288), .B2(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT33), .B(G1976), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(G22), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT84), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(G166), .B2(new_n679), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT85), .B(G1971), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NAND4_X1  g262(.A1(new_n675), .A2(new_n676), .A3(new_n682), .A4(new_n687), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n688), .A2(KEYINPUT34), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(KEYINPUT34), .ZN(new_n690));
  INV_X1    g265(.A(G29), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G25), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT80), .Z(new_n693));
  MUX2_X1   g268(.A(G95), .B(G107), .S(G2105), .Z(new_n694));
  AOI22_X1  g269(.A1(G119), .A2(new_n477), .B1(new_n694), .B2(G2104), .ZN(new_n695));
  INV_X1    g270(.A(G131), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(new_n616), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT81), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n693), .B1(new_n699), .B2(G29), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT35), .B(G1991), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(G16), .A2(G24), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n582), .B2(G16), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(G1986), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n689), .A2(new_n690), .A3(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT86), .B(KEYINPUT36), .Z(new_n708));
  OR2_X1    g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n691), .A2(G32), .ZN(new_n711));
  NAND3_X1  g286(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT89), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT26), .Z(new_n714));
  NAND2_X1  g289(.A1(new_n477), .A2(G129), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n469), .A2(G141), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n471), .A2(G105), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n711), .B1(new_n719), .B2(new_n691), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT27), .B(G1996), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT90), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT91), .ZN(new_n725));
  NOR2_X1   g300(.A1(G4), .A2(G16), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n594), .B2(G16), .ZN(new_n727));
  OAI22_X1  g302(.A1(new_n724), .A2(new_n725), .B1(new_n727), .B2(G1348), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G1348), .B2(new_n727), .ZN(new_n729));
  NOR2_X1   g304(.A1(G16), .A2(G19), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n535), .B2(G16), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(G1341), .Z(new_n732));
  NAND2_X1  g307(.A1(new_n691), .A2(G26), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT28), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n469), .A2(G140), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT87), .Z(new_n736));
  MUX2_X1   g311(.A(G104), .B(G116), .S(G2105), .Z(new_n737));
  AOI22_X1  g312(.A1(G128), .A2(new_n477), .B1(new_n737), .B2(G2104), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n734), .B1(new_n739), .B2(new_n691), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G2067), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n725), .B2(new_n724), .ZN(new_n742));
  NOR2_X1   g317(.A1(G27), .A2(G29), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G164), .B2(G29), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT94), .B(G2078), .Z(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT31), .B(G11), .Z(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT93), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT30), .B(G28), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n748), .B1(new_n691), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(KEYINPUT24), .A2(G34), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(KEYINPUT24), .A2(G34), .ZN(new_n753));
  AOI21_X1  g328(.A(G29), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G160), .B2(G29), .ZN(new_n755));
  OAI221_X1 g330(.A(new_n750), .B1(new_n691), .B2(new_n617), .C1(new_n755), .C2(G2084), .ZN(new_n756));
  AOI211_X1 g331(.A(new_n746), .B(new_n756), .C1(G2084), .C2(new_n755), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n729), .A2(new_n732), .A3(new_n742), .A4(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(G168), .A2(new_n679), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n679), .B2(G21), .ZN(new_n760));
  INV_X1    g335(.A(G1966), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT92), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n691), .A2(G33), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n471), .A2(G103), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(KEYINPUT25), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT25), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n471), .A2(new_n767), .A3(G103), .ZN(new_n768));
  INV_X1    g343(.A(G139), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n766), .B(new_n768), .C1(new_n616), .C2(new_n769), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT88), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n462), .A2(G127), .ZN(new_n772));
  INV_X1    g347(.A(G115), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(new_n470), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n771), .B1(G2105), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n764), .B1(new_n775), .B2(new_n691), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(G2072), .Z(new_n777));
  NAND2_X1  g352(.A1(new_n679), .A2(G5), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G171), .B2(new_n679), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n760), .A2(new_n761), .B1(new_n779), .B2(G1961), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n779), .A2(G1961), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n722), .B2(new_n720), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n691), .A2(G35), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT95), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G162), .B2(new_n691), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G2090), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n763), .A2(new_n777), .A3(new_n783), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n679), .A2(G20), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT23), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n557), .B2(new_n679), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G1956), .ZN(new_n794));
  NOR3_X1   g369(.A1(new_n758), .A2(new_n790), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n709), .A2(new_n710), .A3(new_n795), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT97), .Z(G311));
  XNOR2_X1  g372(.A(new_n796), .B(KEYINPUT98), .ZN(G150));
  AOI22_X1  g373(.A1(new_n498), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n799), .A2(new_n500), .ZN(new_n800));
  INV_X1    g375(.A(G93), .ZN(new_n801));
  INV_X1    g376(.A(G55), .ZN(new_n802));
  OAI22_X1  g377(.A1(new_n503), .A2(new_n801), .B1(new_n802), .B2(new_n506), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(G860), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT37), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n804), .B(KEYINPUT99), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n535), .A2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT99), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n804), .B(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(new_n534), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT38), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n594), .A2(G559), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(KEYINPUT39), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT100), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n805), .B1(new_n816), .B2(KEYINPUT39), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n807), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT101), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OAI211_X1 g398(.A(KEYINPUT101), .B(new_n807), .C1(new_n819), .C2(new_n820), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(G145));
  XNOR2_X1  g400(.A(new_n775), .B(new_n719), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT102), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n487), .B1(new_n469), .B2(G138), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n485), .A2(KEYINPUT4), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n486), .A2(new_n488), .A3(KEYINPUT102), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n830), .A2(new_n493), .A3(new_n831), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n739), .B(new_n832), .Z(new_n833));
  XNOR2_X1  g408(.A(new_n826), .B(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n699), .B(new_n608), .ZN(new_n835));
  MUX2_X1   g410(.A(G106), .B(G118), .S(G2105), .Z(new_n836));
  AOI22_X1  g411(.A1(G130), .A2(new_n477), .B1(new_n836), .B2(G2104), .ZN(new_n837));
  INV_X1    g412(.A(G142), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n837), .B1(new_n838), .B2(new_n616), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n835), .B(new_n839), .Z(new_n840));
  AND2_X1   g415(.A1(new_n834), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n841), .A2(KEYINPUT104), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n834), .A2(new_n840), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n473), .B(new_n481), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n617), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT105), .Z(new_n846));
  NOR3_X1   g421(.A1(new_n842), .A2(new_n843), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n841), .A2(KEYINPUT104), .ZN(new_n848));
  AOI21_X1  g423(.A(G37), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n845), .B1(new_n841), .B2(new_n843), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT103), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT40), .ZN(G395));
  NOR3_X1   g428(.A1(new_n800), .A2(new_n803), .A3(G868), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n813), .B(new_n604), .Z(new_n855));
  NAND2_X1  g430(.A1(G299), .A2(new_n593), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT41), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n593), .B1(new_n555), .B2(new_n556), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n856), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n557), .A2(new_n594), .ZN(new_n861));
  OAI21_X1  g436(.A(KEYINPUT41), .B1(new_n861), .B2(new_n858), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n855), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n861), .A2(new_n858), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n864), .B1(new_n866), .B2(new_n855), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n582), .B(G288), .Z(new_n868));
  XNOR2_X1  g443(.A(new_n575), .B(G166), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT106), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n870), .B1(new_n871), .B2(KEYINPUT42), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n867), .B(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n871), .A2(KEYINPUT42), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n873), .B(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n854), .B1(new_n875), .B2(G868), .ZN(G295));
  AOI21_X1  g451(.A(new_n854), .B1(new_n875), .B2(G868), .ZN(G331));
  NAND3_X1  g452(.A1(new_n560), .A2(G168), .A3(new_n561), .ZN(new_n878));
  NAND2_X1  g453(.A1(G286), .A2(G171), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n813), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT107), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n809), .A2(new_n812), .A3(new_n879), .A4(new_n878), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n813), .A2(KEYINPUT107), .A3(new_n880), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n881), .A2(new_n883), .ZN(new_n887));
  AOI22_X1  g462(.A1(new_n886), .A2(new_n865), .B1(new_n863), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(G37), .B1(new_n888), .B2(new_n870), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT108), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n860), .A2(new_n890), .A3(new_n862), .ZN(new_n891));
  OAI211_X1 g466(.A(KEYINPUT108), .B(KEYINPUT41), .C1(new_n861), .C2(new_n858), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n891), .A2(new_n884), .A3(new_n885), .A4(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n865), .A2(new_n881), .A3(new_n883), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n870), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n889), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n888), .A2(new_n870), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n901), .A2(KEYINPUT43), .A3(new_n889), .ZN(new_n902));
  AOI21_X1  g477(.A(KEYINPUT44), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n889), .A2(new_n897), .A3(KEYINPUT109), .ZN(new_n904));
  AOI21_X1  g479(.A(KEYINPUT109), .B1(new_n889), .B2(new_n897), .ZN(new_n905));
  OAI21_X1  g480(.A(KEYINPUT43), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n901), .A2(new_n899), .A3(new_n889), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n903), .B1(new_n908), .B2(KEYINPUT44), .ZN(G397));
  XNOR2_X1  g484(.A(KEYINPUT110), .B(G1384), .ZN(new_n910));
  AOI21_X1  g485(.A(KEYINPUT45), .B1(new_n832), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n466), .A2(G40), .A3(new_n472), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(G1996), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT112), .ZN(new_n917));
  INV_X1    g492(.A(new_n719), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(G2067), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n739), .B(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n921), .B1(G1996), .B2(new_n918), .ZN(new_n922));
  INV_X1    g497(.A(new_n914), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n919), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(G290), .A2(G1986), .ZN(new_n927));
  XOR2_X1   g502(.A(new_n927), .B(KEYINPUT111), .Z(new_n928));
  NAND2_X1  g503(.A1(G290), .A2(G1986), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n923), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n699), .B(new_n701), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n931), .A2(new_n923), .ZN(new_n932));
  NOR3_X1   g507(.A1(new_n926), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(KEYINPUT116), .B(G8), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n492), .A2(G2104), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n462), .A2(G2105), .ZN(new_n936));
  INV_X1    g511(.A(G126), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n938), .B1(new_n489), .B2(new_n827), .ZN(new_n939));
  AOI21_X1  g514(.A(G1384), .B1(new_n939), .B2(new_n831), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n940), .A2(new_n913), .ZN(new_n941));
  INV_X1    g516(.A(G288), .ZN(new_n942));
  AOI211_X1 g517(.A(new_n934), .B(new_n941), .C1(G1976), .C2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT52), .ZN(new_n944));
  OR2_X1    g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n943), .B(new_n944), .C1(G1976), .C2(new_n942), .ZN(new_n946));
  OR2_X1    g521(.A1(G305), .A2(G1981), .ZN(new_n947));
  XNOR2_X1  g522(.A(KEYINPUT117), .B(G86), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n570), .B1(new_n503), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(G1981), .B1(new_n949), .B2(new_n574), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT49), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n941), .A2(new_n934), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n947), .A2(KEYINPUT49), .A3(new_n950), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n945), .A2(new_n946), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(G303), .A2(G8), .ZN(new_n958));
  XOR2_X1   g533(.A(new_n958), .B(KEYINPUT55), .Z(new_n959));
  NAND3_X1  g534(.A1(new_n832), .A2(KEYINPUT45), .A3(new_n910), .ZN(new_n960));
  INV_X1    g535(.A(G1384), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n494), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n912), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n960), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G1971), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G2090), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n912), .B1(new_n962), .B2(KEYINPUT50), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT113), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT50), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n970), .B1(new_n940), .B2(new_n971), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n832), .A2(new_n970), .A3(new_n971), .A4(new_n961), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n968), .B(new_n969), .C1(new_n972), .C2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n967), .B1(new_n975), .B2(KEYINPUT114), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT114), .ZN(new_n977));
  INV_X1    g552(.A(new_n969), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n832), .A2(new_n971), .A3(new_n961), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT113), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n978), .B1(new_n980), .B2(new_n973), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n977), .B1(new_n981), .B2(new_n968), .ZN(new_n982));
  OAI211_X1 g557(.A(G8), .B(new_n959), .C1(new_n976), .C2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT115), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n975), .A2(KEYINPUT114), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n981), .A2(new_n977), .A3(new_n968), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n985), .A2(new_n986), .A3(new_n967), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT115), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n987), .A2(new_n988), .A3(G8), .A4(new_n959), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n957), .A2(new_n984), .A3(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(G288), .A2(G1976), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n956), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n947), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n954), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n990), .A2(new_n994), .A3(KEYINPUT118), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT118), .B1(new_n990), .B2(new_n994), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(G1384), .B1(new_n489), .B2(new_n493), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT119), .B1(new_n998), .B2(new_n971), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n998), .A2(KEYINPUT119), .A3(new_n971), .ZN(new_n1000));
  OAI221_X1 g575(.A(new_n913), .B1(new_n940), .B2(new_n971), .C1(new_n999), .C2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G1956), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT122), .ZN(new_n1003));
  XNOR2_X1  g578(.A(KEYINPUT56), .B(G2072), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n960), .A2(new_n964), .A3(new_n1004), .ZN(new_n1005));
  AOI22_X1  g580(.A1(new_n1001), .A2(new_n1002), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n960), .A2(new_n964), .A3(KEYINPUT122), .A4(new_n1004), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n553), .B(KEYINPUT57), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1006), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT123), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n980), .A2(new_n973), .ZN(new_n1012));
  AOI21_X1  g587(.A(G1348), .B1(new_n1012), .B2(new_n969), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n941), .A2(new_n920), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1011), .B(new_n594), .C1(new_n1013), .C2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n913), .B1(new_n1000), .B2(new_n999), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n940), .A2(new_n971), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1002), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1005), .A2(new_n1003), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1019), .A2(new_n1007), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n1008), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1016), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1014), .B1(new_n981), .B2(G1348), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1011), .B1(new_n1024), .B2(new_n594), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1010), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT124), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT124), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1028), .B(new_n1010), .C1(new_n1023), .C2(new_n1025), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT125), .ZN(new_n1030));
  OAI211_X1 g605(.A(KEYINPUT60), .B(new_n1014), .C1(new_n981), .C2(G1348), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1030), .B1(new_n1031), .B2(new_n594), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1031), .A2(new_n594), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1031), .A2(new_n1030), .A3(new_n594), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT60), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n1034), .A2(new_n1035), .B1(new_n1036), .B2(new_n1024), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT61), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1009), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1021), .A2(new_n1008), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1038), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1010), .A2(new_n1022), .A3(KEYINPUT61), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n960), .A2(new_n964), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(new_n915), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n940), .A2(new_n913), .ZN(new_n1045));
  XOR2_X1   g620(.A(KEYINPUT58), .B(G1341), .Z(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n534), .B1(new_n1044), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT59), .ZN(new_n1049));
  XNOR2_X1  g624(.A(new_n1048), .B(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1041), .A2(new_n1042), .A3(new_n1050), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1027), .B(new_n1029), .C1(new_n1037), .C2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n981), .A2(G1961), .ZN(new_n1054));
  INV_X1    g629(.A(G2078), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT53), .B1(new_n1043), .B2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT45), .B1(new_n832), .B2(new_n961), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT120), .B1(new_n1058), .B2(new_n912), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT120), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1060), .B(new_n913), .C1(new_n940), .C2(KEYINPUT45), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n998), .A2(KEYINPUT45), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1059), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1055), .A2(KEYINPUT53), .ZN(new_n1064));
  OR2_X1    g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(G301), .B1(new_n1057), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT53), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1067), .B1(new_n965), .B2(G2078), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n913), .A2(KEYINPUT126), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT126), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1064), .B1(new_n912), .B2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n960), .A2(new_n1069), .A3(new_n1071), .ZN(new_n1072));
  OAI221_X1 g647(.A(new_n1068), .B1(new_n911), .B2(new_n1072), .C1(new_n981), .C2(G1961), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1073), .A2(new_n562), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1053), .B1(new_n1066), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1053), .B1(new_n1073), .B2(G171), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1057), .A2(new_n1065), .A3(G301), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G2084), .ZN(new_n1080));
  AOI22_X1  g655(.A1(new_n1063), .A2(new_n761), .B1(new_n981), .B2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(G168), .A2(new_n934), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G8), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1063), .A2(new_n761), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n981), .A2(new_n1080), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT51), .B1(new_n1088), .B2(new_n1082), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1082), .A2(KEYINPUT51), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(new_n1081), .B2(new_n934), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1084), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1079), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1066), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT62), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1094), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1083), .B1(new_n1081), .B2(new_n1085), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1098));
  INV_X1    g673(.A(new_n934), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  AOI22_X1  g675(.A1(KEYINPUT51), .A2(new_n1097), .B1(new_n1100), .B2(new_n1090), .ZN(new_n1101));
  OAI21_X1  g676(.A(KEYINPUT62), .B1(new_n1101), .B2(new_n1084), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1052), .A2(new_n1093), .B1(new_n1096), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n984), .A2(new_n989), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1104), .A2(new_n957), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n967), .B1(new_n1001), .B2(G2090), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1106), .A2(new_n1099), .ZN(new_n1107));
  OR2_X1    g682(.A1(new_n1107), .A2(new_n959), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n997), .B1(new_n1103), .B2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1100), .A2(G286), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1104), .A2(new_n1111), .A3(new_n957), .A4(new_n1108), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT63), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1112), .A2(KEYINPUT121), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n959), .B1(new_n987), .B2(G8), .ZN(new_n1115));
  NOR4_X1   g690(.A1(new_n1115), .A2(new_n1100), .A3(new_n1113), .A4(G286), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1105), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT121), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n933), .B1(new_n1110), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n917), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1122), .A2(KEYINPUT46), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(KEYINPUT46), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n914), .B1(new_n921), .B2(new_n918), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n1126), .B(KEYINPUT47), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n701), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n699), .A2(new_n1129), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n925), .A2(new_n1130), .B1(new_n920), .B2(new_n739), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1128), .B1(new_n1131), .B2(new_n923), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n928), .A2(new_n923), .ZN(new_n1133));
  XOR2_X1   g708(.A(new_n1133), .B(KEYINPUT48), .Z(new_n1134));
  OAI211_X1 g709(.A(new_n1134), .B(new_n925), .C1(new_n923), .C2(new_n931), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1127), .A2(new_n1132), .A3(new_n1135), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1131), .A2(new_n1128), .A3(new_n923), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1121), .A2(new_n1138), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g714(.A1(new_n849), .A2(new_n851), .ZN(new_n1141));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n902), .ZN(new_n1142));
  NOR2_X1   g716(.A1(G227), .A2(new_n460), .ZN(new_n1143));
  OAI211_X1 g717(.A(new_n1143), .B(new_n669), .C1(new_n633), .C2(new_n634), .ZN(new_n1144));
  NOR3_X1   g718(.A1(new_n1141), .A2(new_n1142), .A3(new_n1144), .ZN(G308));
  OR3_X1    g719(.A1(new_n1141), .A2(new_n1142), .A3(new_n1144), .ZN(G225));
endmodule


