

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580;

  XNOR2_X1 U322 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U323 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n290) );
  INV_X1 U324 ( .A(KEYINPUT110), .ZN(n378) );
  XNOR2_X1 U325 ( .A(n390), .B(n332), .ZN(n333) );
  XNOR2_X1 U326 ( .A(n406), .B(n290), .ZN(n564) );
  XOR2_X1 U327 ( .A(KEYINPUT36), .B(n557), .Z(n578) );
  XOR2_X1 U328 ( .A(n343), .B(n342), .Z(n557) );
  XNOR2_X1 U329 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U330 ( .A(n453), .B(n452), .ZN(G1349GAT) );
  XOR2_X1 U331 ( .A(G127GAT), .B(G134GAT), .Z(n292) );
  XNOR2_X1 U332 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n291) );
  XNOR2_X1 U333 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U334 ( .A(G113GAT), .B(n293), .Z(n441) );
  XOR2_X1 U335 ( .A(KEYINPUT82), .B(KEYINPUT17), .Z(n295) );
  XNOR2_X1 U336 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n294) );
  XNOR2_X1 U337 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U338 ( .A(G169GAT), .B(n296), .Z(n401) );
  XOR2_X1 U339 ( .A(G99GAT), .B(G190GAT), .Z(n298) );
  XNOR2_X1 U340 ( .A(G15GAT), .B(G183GAT), .ZN(n297) );
  XNOR2_X1 U341 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U342 ( .A(n401), .B(n299), .Z(n301) );
  NAND2_X1 U343 ( .A1(G227GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U344 ( .A(n301), .B(n300), .ZN(n309) );
  XOR2_X1 U345 ( .A(KEYINPUT80), .B(G71GAT), .Z(n303) );
  XNOR2_X1 U346 ( .A(KEYINPUT20), .B(G176GAT), .ZN(n302) );
  XNOR2_X1 U347 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U348 ( .A(KEYINPUT81), .B(KEYINPUT83), .Z(n305) );
  XNOR2_X1 U349 ( .A(G43GAT), .B(KEYINPUT65), .ZN(n304) );
  XNOR2_X1 U350 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U351 ( .A(n307), .B(n306), .Z(n308) );
  XNOR2_X1 U352 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U353 ( .A(n441), .B(n310), .ZN(n454) );
  XOR2_X1 U354 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n446) );
  XOR2_X1 U355 ( .A(G22GAT), .B(G197GAT), .Z(n312) );
  XNOR2_X1 U356 ( .A(G169GAT), .B(G113GAT), .ZN(n311) );
  XNOR2_X1 U357 ( .A(n312), .B(n311), .ZN(n327) );
  XOR2_X1 U358 ( .A(G15GAT), .B(G1GAT), .Z(n355) );
  XOR2_X1 U359 ( .A(G29GAT), .B(G43GAT), .Z(n314) );
  XNOR2_X1 U360 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n313) );
  XNOR2_X1 U361 ( .A(n314), .B(n313), .ZN(n334) );
  XOR2_X1 U362 ( .A(n355), .B(n334), .Z(n316) );
  XNOR2_X1 U363 ( .A(G36GAT), .B(G50GAT), .ZN(n315) );
  XNOR2_X1 U364 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U365 ( .A(KEYINPUT69), .B(KEYINPUT68), .Z(n318) );
  NAND2_X1 U366 ( .A1(G229GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U367 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U368 ( .A(n320), .B(n319), .Z(n325) );
  XOR2_X1 U369 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n322) );
  XNOR2_X1 U370 ( .A(G141GAT), .B(G8GAT), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U372 ( .A(n323), .B(KEYINPUT30), .ZN(n324) );
  XNOR2_X1 U373 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U374 ( .A(n327), .B(n326), .ZN(n551) );
  XOR2_X1 U375 ( .A(KEYINPUT9), .B(KEYINPUT78), .Z(n329) );
  XNOR2_X1 U376 ( .A(KEYINPUT10), .B(KEYINPUT79), .ZN(n328) );
  XNOR2_X1 U377 ( .A(n329), .B(n328), .ZN(n343) );
  XOR2_X1 U378 ( .A(KEYINPUT11), .B(G92GAT), .Z(n331) );
  XNOR2_X1 U379 ( .A(G134GAT), .B(G106GAT), .ZN(n330) );
  XNOR2_X1 U380 ( .A(n331), .B(n330), .ZN(n336) );
  XOR2_X1 U381 ( .A(G36GAT), .B(G190GAT), .Z(n390) );
  AND2_X1 U382 ( .A1(G232GAT), .A2(G233GAT), .ZN(n332) );
  XOR2_X1 U383 ( .A(n336), .B(n335), .Z(n341) );
  XOR2_X1 U384 ( .A(G162GAT), .B(KEYINPUT77), .Z(n338) );
  XNOR2_X1 U385 ( .A(G50GAT), .B(G218GAT), .ZN(n337) );
  XNOR2_X1 U386 ( .A(n338), .B(n337), .ZN(n413) );
  XNOR2_X1 U387 ( .A(G99GAT), .B(G85GAT), .ZN(n339) );
  XNOR2_X1 U388 ( .A(n339), .B(KEYINPUT74), .ZN(n367) );
  XNOR2_X1 U389 ( .A(n413), .B(n367), .ZN(n340) );
  XNOR2_X1 U390 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U391 ( .A(G22GAT), .B(G155GAT), .Z(n410) );
  XOR2_X1 U392 ( .A(KEYINPUT15), .B(G64GAT), .Z(n345) );
  XNOR2_X1 U393 ( .A(G127GAT), .B(G211GAT), .ZN(n344) );
  XNOR2_X1 U394 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U395 ( .A(n410), .B(n346), .Z(n348) );
  NAND2_X1 U396 ( .A1(G231GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U397 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U398 ( .A(n349), .B(KEYINPUT12), .Z(n353) );
  XOR2_X1 U399 ( .A(G57GAT), .B(KEYINPUT13), .Z(n351) );
  XNOR2_X1 U400 ( .A(G71GAT), .B(G78GAT), .ZN(n350) );
  XNOR2_X1 U401 ( .A(n351), .B(n350), .ZN(n363) );
  XNOR2_X1 U402 ( .A(n363), .B(KEYINPUT14), .ZN(n352) );
  XNOR2_X1 U403 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U404 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U405 ( .A(G8GAT), .B(G183GAT), .Z(n389) );
  XNOR2_X1 U406 ( .A(n356), .B(n389), .ZN(n544) );
  INV_X1 U407 ( .A(n544), .ZN(n575) );
  NOR2_X1 U408 ( .A1(n578), .A2(n575), .ZN(n357) );
  XNOR2_X1 U409 ( .A(n357), .B(KEYINPUT45), .ZN(n376) );
  XOR2_X1 U410 ( .A(G148GAT), .B(G204GAT), .Z(n359) );
  XNOR2_X1 U411 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n358) );
  XNOR2_X1 U412 ( .A(n359), .B(n358), .ZN(n420) );
  XNOR2_X1 U413 ( .A(G176GAT), .B(G92GAT), .ZN(n360) );
  XNOR2_X1 U414 ( .A(n360), .B(G64GAT), .ZN(n393) );
  XNOR2_X1 U415 ( .A(n420), .B(n393), .ZN(n375) );
  XOR2_X1 U416 ( .A(KEYINPUT72), .B(KEYINPUT32), .Z(n362) );
  XNOR2_X1 U417 ( .A(G120GAT), .B(KEYINPUT75), .ZN(n361) );
  XNOR2_X1 U418 ( .A(n362), .B(n361), .ZN(n364) );
  XOR2_X1 U419 ( .A(n364), .B(n363), .Z(n373) );
  XOR2_X1 U420 ( .A(KEYINPUT33), .B(KEYINPUT71), .Z(n366) );
  XNOR2_X1 U421 ( .A(KEYINPUT70), .B(KEYINPUT76), .ZN(n365) );
  XNOR2_X1 U422 ( .A(n366), .B(n365), .ZN(n371) );
  XOR2_X1 U423 ( .A(n367), .B(KEYINPUT31), .Z(n369) );
  NAND2_X1 U424 ( .A1(G230GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U425 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U426 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U427 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U428 ( .A(n375), .B(n374), .ZN(n570) );
  NAND2_X1 U429 ( .A1(n376), .A2(n570), .ZN(n377) );
  NOR2_X1 U430 ( .A1(n551), .A2(n377), .ZN(n379) );
  XNOR2_X1 U431 ( .A(n379), .B(n378), .ZN(n387) );
  XOR2_X1 U432 ( .A(KEYINPUT46), .B(KEYINPUT109), .Z(n382) );
  XNOR2_X1 U433 ( .A(n570), .B(KEYINPUT41), .ZN(n380) );
  XNOR2_X1 U434 ( .A(n380), .B(KEYINPUT64), .ZN(n539) );
  NAND2_X1 U435 ( .A1(n539), .A2(n551), .ZN(n381) );
  XNOR2_X1 U436 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U437 ( .A(KEYINPUT108), .B(n575), .ZN(n554) );
  NAND2_X1 U438 ( .A1(n383), .A2(n554), .ZN(n384) );
  NOR2_X1 U439 ( .A1(n557), .A2(n384), .ZN(n385) );
  XNOR2_X1 U440 ( .A(KEYINPUT47), .B(n385), .ZN(n386) );
  NAND2_X1 U441 ( .A1(n387), .A2(n386), .ZN(n388) );
  XNOR2_X1 U442 ( .A(KEYINPUT48), .B(n388), .ZN(n518) );
  XOR2_X1 U443 ( .A(KEYINPUT94), .B(KEYINPUT96), .Z(n392) );
  XNOR2_X1 U444 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U445 ( .A(n392), .B(n391), .ZN(n397) );
  XOR2_X1 U446 ( .A(n393), .B(KEYINPUT95), .Z(n395) );
  NAND2_X1 U447 ( .A1(G226GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U448 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U449 ( .A(n397), .B(n396), .Z(n399) );
  XNOR2_X1 U450 ( .A(G204GAT), .B(G218GAT), .ZN(n398) );
  XNOR2_X1 U451 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U452 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U453 ( .A(KEYINPUT85), .B(KEYINPUT86), .Z(n403) );
  XNOR2_X1 U454 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n402) );
  XNOR2_X1 U455 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U456 ( .A(G197GAT), .B(n404), .ZN(n424) );
  XNOR2_X1 U457 ( .A(n405), .B(n424), .ZN(n507) );
  NAND2_X1 U458 ( .A1(n518), .A2(n507), .ZN(n406) );
  XOR2_X1 U459 ( .A(KEYINPUT24), .B(KEYINPUT89), .Z(n408) );
  XNOR2_X1 U460 ( .A(KEYINPUT23), .B(KEYINPUT88), .ZN(n407) );
  XNOR2_X1 U461 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U462 ( .A(n409), .B(KEYINPUT84), .Z(n412) );
  XNOR2_X1 U463 ( .A(n410), .B(G78GAT), .ZN(n411) );
  XNOR2_X1 U464 ( .A(n412), .B(n411), .ZN(n417) );
  XOR2_X1 U465 ( .A(n413), .B(KEYINPUT22), .Z(n415) );
  NAND2_X1 U466 ( .A1(G228GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U467 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U468 ( .A(n417), .B(n416), .Z(n422) );
  XOR2_X1 U469 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n419) );
  XNOR2_X1 U470 ( .A(G141GAT), .B(KEYINPUT87), .ZN(n418) );
  XNOR2_X1 U471 ( .A(n419), .B(n418), .ZN(n436) );
  XNOR2_X1 U472 ( .A(n436), .B(n420), .ZN(n421) );
  XNOR2_X1 U473 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U474 ( .A(n424), .B(n423), .Z(n460) );
  XOR2_X1 U475 ( .A(KEYINPUT6), .B(G57GAT), .Z(n426) );
  XNOR2_X1 U476 ( .A(G1GAT), .B(G148GAT), .ZN(n425) );
  XNOR2_X1 U477 ( .A(n426), .B(n425), .ZN(n430) );
  XOR2_X1 U478 ( .A(KEYINPUT4), .B(KEYINPUT1), .Z(n428) );
  XNOR2_X1 U479 ( .A(KEYINPUT90), .B(KEYINPUT91), .ZN(n427) );
  XNOR2_X1 U480 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U481 ( .A(n430), .B(n429), .Z(n435) );
  XOR2_X1 U482 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n432) );
  NAND2_X1 U483 ( .A1(G225GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U484 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U485 ( .A(KEYINPUT5), .B(n433), .ZN(n434) );
  XNOR2_X1 U486 ( .A(n435), .B(n434), .ZN(n440) );
  XOR2_X1 U487 ( .A(G85GAT), .B(G155GAT), .Z(n438) );
  XNOR2_X1 U488 ( .A(n436), .B(G162GAT), .ZN(n437) );
  XNOR2_X1 U489 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U490 ( .A(n440), .B(n439), .Z(n443) );
  XNOR2_X1 U491 ( .A(G29GAT), .B(n441), .ZN(n442) );
  XNOR2_X1 U492 ( .A(n443), .B(n442), .ZN(n505) );
  INV_X1 U493 ( .A(n505), .ZN(n563) );
  AND2_X1 U494 ( .A1(n460), .A2(n563), .ZN(n444) );
  NAND2_X1 U495 ( .A1(n564), .A2(n444), .ZN(n445) );
  XNOR2_X1 U496 ( .A(n446), .B(n445), .ZN(n447) );
  NOR2_X1 U497 ( .A1(n454), .A2(n447), .ZN(n449) );
  INV_X1 U498 ( .A(KEYINPUT121), .ZN(n448) );
  XNOR2_X1 U499 ( .A(n449), .B(n448), .ZN(n558) );
  XNOR2_X1 U500 ( .A(n539), .B(KEYINPUT102), .ZN(n524) );
  NAND2_X1 U501 ( .A1(n558), .A2(n524), .ZN(n453) );
  XOR2_X1 U502 ( .A(G176GAT), .B(KEYINPUT122), .Z(n451) );
  XNOR2_X1 U503 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n450) );
  NAND2_X1 U504 ( .A1(n570), .A2(n551), .ZN(n483) );
  XNOR2_X1 U505 ( .A(KEYINPUT27), .B(n507), .ZN(n463) );
  NAND2_X1 U506 ( .A1(n505), .A2(n463), .ZN(n516) );
  INV_X1 U507 ( .A(n454), .ZN(n520) );
  XNOR2_X1 U508 ( .A(KEYINPUT28), .B(KEYINPUT66), .ZN(n455) );
  XOR2_X1 U509 ( .A(n455), .B(n460), .Z(n519) );
  OR2_X1 U510 ( .A1(n520), .A2(n519), .ZN(n456) );
  NOR2_X1 U511 ( .A1(n516), .A2(n456), .ZN(n468) );
  NAND2_X1 U512 ( .A1(n520), .A2(n507), .ZN(n457) );
  XNOR2_X1 U513 ( .A(n457), .B(KEYINPUT98), .ZN(n458) );
  NAND2_X1 U514 ( .A1(n458), .A2(n460), .ZN(n459) );
  XNOR2_X1 U515 ( .A(n459), .B(KEYINPUT25), .ZN(n465) );
  NOR2_X1 U516 ( .A1(n520), .A2(n460), .ZN(n462) );
  XNOR2_X1 U517 ( .A(KEYINPUT97), .B(KEYINPUT26), .ZN(n461) );
  XNOR2_X1 U518 ( .A(n462), .B(n461), .ZN(n535) );
  INV_X1 U519 ( .A(n535), .ZN(n566) );
  AND2_X1 U520 ( .A1(n463), .A2(n566), .ZN(n464) );
  NOR2_X1 U521 ( .A1(n465), .A2(n464), .ZN(n466) );
  NOR2_X1 U522 ( .A1(n505), .A2(n466), .ZN(n467) );
  NOR2_X1 U523 ( .A1(n468), .A2(n467), .ZN(n479) );
  NOR2_X1 U524 ( .A1(n557), .A2(n575), .ZN(n469) );
  XOR2_X1 U525 ( .A(KEYINPUT16), .B(n469), .Z(n470) );
  OR2_X1 U526 ( .A1(n479), .A2(n470), .ZN(n493) );
  NOR2_X1 U527 ( .A1(n483), .A2(n493), .ZN(n477) );
  NAND2_X1 U528 ( .A1(n505), .A2(n477), .ZN(n471) );
  XNOR2_X1 U529 ( .A(KEYINPUT34), .B(n471), .ZN(n472) );
  XNOR2_X1 U530 ( .A(G1GAT), .B(n472), .ZN(G1324GAT) );
  XOR2_X1 U531 ( .A(G8GAT), .B(KEYINPUT99), .Z(n474) );
  NAND2_X1 U532 ( .A1(n477), .A2(n507), .ZN(n473) );
  XNOR2_X1 U533 ( .A(n474), .B(n473), .ZN(G1325GAT) );
  XOR2_X1 U534 ( .A(G15GAT), .B(KEYINPUT35), .Z(n476) );
  NAND2_X1 U535 ( .A1(n477), .A2(n520), .ZN(n475) );
  XNOR2_X1 U536 ( .A(n476), .B(n475), .ZN(G1326GAT) );
  NAND2_X1 U537 ( .A1(n477), .A2(n519), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n478), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U539 ( .A(G29GAT), .B(KEYINPUT39), .Z(n487) );
  XOR2_X1 U540 ( .A(KEYINPUT100), .B(KEYINPUT37), .Z(n482) );
  NOR2_X1 U541 ( .A1(n578), .A2(n479), .ZN(n480) );
  NAND2_X1 U542 ( .A1(n480), .A2(n575), .ZN(n481) );
  XNOR2_X1 U543 ( .A(n482), .B(n481), .ZN(n504) );
  NOR2_X1 U544 ( .A1(n483), .A2(n504), .ZN(n484) );
  XOR2_X1 U545 ( .A(KEYINPUT101), .B(n484), .Z(n485) );
  XNOR2_X1 U546 ( .A(KEYINPUT38), .B(n485), .ZN(n491) );
  NAND2_X1 U547 ( .A1(n505), .A2(n491), .ZN(n486) );
  XNOR2_X1 U548 ( .A(n487), .B(n486), .ZN(G1328GAT) );
  NAND2_X1 U549 ( .A1(n491), .A2(n507), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n488), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U551 ( .A1(n491), .A2(n520), .ZN(n489) );
  XNOR2_X1 U552 ( .A(n489), .B(KEYINPUT40), .ZN(n490) );
  XNOR2_X1 U553 ( .A(G43GAT), .B(n490), .ZN(G1330GAT) );
  NAND2_X1 U554 ( .A1(n519), .A2(n491), .ZN(n492) );
  XNOR2_X1 U555 ( .A(G50GAT), .B(n492), .ZN(G1331GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT42), .B(KEYINPUT104), .Z(n496) );
  INV_X1 U557 ( .A(n551), .ZN(n567) );
  NAND2_X1 U558 ( .A1(n524), .A2(n567), .ZN(n503) );
  OR2_X1 U559 ( .A1(n493), .A2(n503), .ZN(n494) );
  XNOR2_X1 U560 ( .A(n494), .B(KEYINPUT103), .ZN(n500) );
  NAND2_X1 U561 ( .A1(n500), .A2(n505), .ZN(n495) );
  XNOR2_X1 U562 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U563 ( .A(G57GAT), .B(n497), .Z(G1332GAT) );
  NAND2_X1 U564 ( .A1(n507), .A2(n500), .ZN(n498) );
  XNOR2_X1 U565 ( .A(n498), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U566 ( .A1(n520), .A2(n500), .ZN(n499) );
  XNOR2_X1 U567 ( .A(n499), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U568 ( .A(G78GAT), .B(KEYINPUT43), .Z(n502) );
  NAND2_X1 U569 ( .A1(n500), .A2(n519), .ZN(n501) );
  XNOR2_X1 U570 ( .A(n502), .B(n501), .ZN(G1335GAT) );
  NOR2_X1 U571 ( .A1(n504), .A2(n503), .ZN(n511) );
  NAND2_X1 U572 ( .A1(n505), .A2(n511), .ZN(n506) );
  XNOR2_X1 U573 ( .A(G85GAT), .B(n506), .ZN(G1336GAT) );
  XOR2_X1 U574 ( .A(G92GAT), .B(KEYINPUT105), .Z(n509) );
  NAND2_X1 U575 ( .A1(n511), .A2(n507), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n509), .B(n508), .ZN(G1337GAT) );
  NAND2_X1 U577 ( .A1(n520), .A2(n511), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n510), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U579 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n515) );
  XOR2_X1 U580 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n513) );
  NAND2_X1 U581 ( .A1(n511), .A2(n519), .ZN(n512) );
  XNOR2_X1 U582 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U583 ( .A(n515), .B(n514), .ZN(G1339GAT) );
  INV_X1 U584 ( .A(n516), .ZN(n517) );
  NAND2_X1 U585 ( .A1(n518), .A2(n517), .ZN(n536) );
  NOR2_X1 U586 ( .A1(n519), .A2(n536), .ZN(n521) );
  NAND2_X1 U587 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U588 ( .A(KEYINPUT111), .B(n522), .ZN(n530) );
  NAND2_X1 U589 ( .A1(n530), .A2(n551), .ZN(n523) );
  XNOR2_X1 U590 ( .A(G113GAT), .B(n523), .ZN(G1340GAT) );
  XOR2_X1 U591 ( .A(G120GAT), .B(KEYINPUT49), .Z(n526) );
  NAND2_X1 U592 ( .A1(n530), .A2(n524), .ZN(n525) );
  XNOR2_X1 U593 ( .A(n526), .B(n525), .ZN(G1341GAT) );
  INV_X1 U594 ( .A(n530), .ZN(n527) );
  NOR2_X1 U595 ( .A1(n554), .A2(n527), .ZN(n528) );
  XOR2_X1 U596 ( .A(KEYINPUT50), .B(n528), .Z(n529) );
  XNOR2_X1 U597 ( .A(G127GAT), .B(n529), .ZN(G1342GAT) );
  AND2_X1 U598 ( .A1(n530), .A2(n557), .ZN(n534) );
  XOR2_X1 U599 ( .A(KEYINPUT112), .B(KEYINPUT51), .Z(n532) );
  XNOR2_X1 U600 ( .A(G134GAT), .B(KEYINPUT113), .ZN(n531) );
  XNOR2_X1 U601 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U602 ( .A(n534), .B(n533), .ZN(G1343GAT) );
  NOR2_X1 U603 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n537), .B(KEYINPUT114), .ZN(n548) );
  NAND2_X1 U605 ( .A1(n551), .A2(n548), .ZN(n538) );
  XNOR2_X1 U606 ( .A(G141GAT), .B(n538), .ZN(G1344GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT52), .B(KEYINPUT53), .Z(n541) );
  NAND2_X1 U608 ( .A1(n539), .A2(n548), .ZN(n540) );
  XNOR2_X1 U609 ( .A(n541), .B(n540), .ZN(n543) );
  XOR2_X1 U610 ( .A(G148GAT), .B(KEYINPUT115), .Z(n542) );
  XNOR2_X1 U611 ( .A(n543), .B(n542), .ZN(G1345GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n546) );
  NAND2_X1 U613 ( .A1(n544), .A2(n548), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U615 ( .A(G155GAT), .B(n547), .ZN(G1346GAT) );
  NAND2_X1 U616 ( .A1(n548), .A2(n557), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n549), .B(KEYINPUT118), .ZN(n550) );
  XNOR2_X1 U618 ( .A(G162GAT), .B(n550), .ZN(G1347GAT) );
  NAND2_X1 U619 ( .A1(n551), .A2(n558), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n552), .B(G169GAT), .ZN(G1348GAT) );
  INV_X1 U621 ( .A(n558), .ZN(n553) );
  NOR2_X1 U622 ( .A1(n554), .A2(n553), .ZN(n556) );
  XNOR2_X1 U623 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(G1350GAT) );
  NAND2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(KEYINPUT58), .ZN(n560) );
  XNOR2_X1 U627 ( .A(G190GAT), .B(n560), .ZN(G1351GAT) );
  XNOR2_X1 U628 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n561), .B(KEYINPUT60), .ZN(n562) );
  XOR2_X1 U630 ( .A(KEYINPUT124), .B(n562), .Z(n569) );
  AND2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n565) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n577) );
  OR2_X1 U633 ( .A1(n577), .A2(n567), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(G1352GAT) );
  NOR2_X1 U635 ( .A1(n577), .A2(n570), .ZN(n574) );
  XOR2_X1 U636 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n572) );
  XNOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n577), .ZN(n576) );
  XOR2_X1 U641 ( .A(G211GAT), .B(n576), .Z(G1354GAT) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U643 ( .A(KEYINPUT62), .B(n579), .Z(n580) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(n580), .ZN(G1355GAT) );
endmodule

