//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 0 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1289, new_n1290, new_n1291,
    new_n1292, new_n1293, new_n1294, new_n1295, new_n1296, new_n1297,
    new_n1298, new_n1299, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  INV_X1    g0014(.A(new_n201), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n212), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  INV_X1    g0025(.A(G77), .ZN(new_n226));
  INV_X1    g0026(.A(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G107), .ZN(new_n228));
  INV_X1    g0028(.A(G264), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n225), .B1(new_n226), .B2(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n209), .B1(new_n224), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT64), .ZN(new_n232));
  INV_X1    g0032(.A(KEYINPUT1), .ZN(new_n233));
  OR2_X1    g0033(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n232), .A2(new_n233), .ZN(new_n235));
  NAND3_X1  g0035(.A1(new_n218), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n236), .B(KEYINPUT65), .Z(G361));
  XOR2_X1   g0037(.A(G250), .B(G257), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT66), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  INV_X1    g0042(.A(G232), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(KEYINPUT2), .B(G226), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n241), .B(new_n246), .ZN(G358));
  XNOR2_X1  g0047(.A(G50), .B(G68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n248), .B(new_n249), .Z(new_n250));
  XOR2_X1   g0050(.A(G87), .B(G97), .Z(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  OAI211_X1 g0055(.A(new_n206), .B(G45), .C1(new_n255), .C2(KEYINPUT5), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT78), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G45), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(G1), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT5), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G41), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n260), .A2(KEYINPUT78), .A3(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n261), .A2(G41), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G274), .ZN(new_n266));
  AND2_X1   g0066(.A1(G1), .A2(G13), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND4_X1  g0069(.A1(new_n258), .A2(new_n263), .A3(new_n265), .A4(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n267), .A2(new_n268), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n272), .B1(new_n256), .B2(new_n264), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n270), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT72), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT3), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(KEYINPUT72), .A2(KEYINPUT3), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(G33), .A3(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT3), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n229), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n279), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT80), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n276), .A2(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n281), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G303), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n279), .A2(G257), .A3(new_n282), .A4(new_n281), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n279), .A2(KEYINPUT80), .A3(new_n281), .A4(new_n283), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n286), .A2(new_n289), .A3(new_n290), .A4(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n274), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT21), .ZN(new_n295));
  NAND3_X1  g0095(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n296));
  INV_X1    g0096(.A(G116), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n296), .A2(new_n213), .B1(G20), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(G33), .A2(G283), .ZN(new_n299));
  INV_X1    g0099(.A(G97), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n299), .B(new_n207), .C1(G33), .C2(new_n300), .ZN(new_n301));
  AND3_X1   g0101(.A1(new_n298), .A2(KEYINPUT20), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(KEYINPUT20), .B1(new_n298), .B2(new_n301), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n297), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n296), .A2(new_n213), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n206), .A2(G33), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n309), .A2(new_n305), .A3(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n307), .B1(new_n311), .B2(new_n297), .ZN(new_n312));
  OAI21_X1  g0112(.A(G169), .B1(new_n304), .B2(new_n312), .ZN(new_n313));
  NOR3_X1   g0113(.A1(new_n294), .A2(new_n295), .A3(new_n313), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n270), .B(G179), .C1(new_n271), .C2(new_n273), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n315), .B1(new_n292), .B2(new_n293), .ZN(new_n316));
  OR2_X1    g0116(.A1(new_n304), .A2(new_n312), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT81), .B1(new_n314), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n292), .A2(new_n293), .ZN(new_n320));
  INV_X1    g0120(.A(new_n274), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n313), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n322), .A2(KEYINPUT21), .A3(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT81), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n316), .A2(new_n317), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n295), .B1(new_n294), .B2(new_n313), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n319), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n304), .A2(new_n312), .ZN(new_n330));
  INV_X1    g0130(.A(G200), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n330), .B1(new_n294), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT82), .ZN(new_n333));
  AND2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  XOR2_X1   g0134(.A(KEYINPUT74), .B(G190), .Z(new_n335));
  NAND2_X1  g0135(.A1(new_n294), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n336), .B1(new_n332), .B2(new_n333), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n329), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n206), .A2(G20), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G50), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n341), .B(KEYINPUT67), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n306), .A2(new_n308), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n342), .A2(new_n344), .B1(G50), .B2(new_n305), .ZN(new_n345));
  XNOR2_X1  g0145(.A(KEYINPUT8), .B(G58), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n280), .A2(G20), .ZN(new_n348));
  NOR2_X1   g0148(.A1(G20), .A2(G33), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n347), .A2(new_n348), .B1(G150), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n203), .A2(G20), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n309), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n345), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT69), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NOR3_X1   g0155(.A1(new_n345), .A2(KEYINPUT69), .A3(new_n352), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT9), .ZN(new_n358));
  XNOR2_X1  g0158(.A(KEYINPUT3), .B(G33), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n359), .A2(G222), .A3(new_n282), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(G1698), .ZN(new_n361));
  INV_X1    g0161(.A(G223), .ZN(new_n362));
  OAI221_X1 g0162(.A(new_n360), .B1(new_n226), .B2(new_n359), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n293), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n365));
  NOR3_X1   g0165(.A1(new_n293), .A2(new_n266), .A3(new_n365), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n272), .A2(new_n365), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n366), .B1(G226), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G200), .ZN(new_n370));
  AND2_X1   g0170(.A1(new_n358), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT10), .ZN(new_n372));
  INV_X1    g0172(.A(G190), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g0174(.A(new_n374), .B(KEYINPUT70), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT9), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n376), .B1(new_n355), .B2(new_n356), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n371), .A2(new_n372), .A3(new_n375), .A4(new_n377), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n375), .A2(new_n377), .A3(new_n358), .A4(new_n370), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT10), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n369), .A2(G179), .ZN(new_n382));
  INV_X1    g0182(.A(G169), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n353), .B1(new_n383), .B2(new_n369), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n382), .B1(new_n384), .B2(KEYINPUT68), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n385), .B1(KEYINPUT68), .B2(new_n384), .ZN(new_n386));
  OR3_X1    g0186(.A1(new_n305), .A2(KEYINPUT12), .A3(G68), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT12), .B1(new_n305), .B2(G68), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n340), .A2(G68), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n348), .A2(G77), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n207), .B2(G68), .ZN(new_n392));
  INV_X1    g0192(.A(new_n349), .ZN(new_n393));
  OAI22_X1  g0193(.A1(new_n392), .A2(KEYINPUT71), .B1(new_n202), .B2(new_n393), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n392), .A2(KEYINPUT71), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n308), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT11), .ZN(new_n397));
  OAI221_X1 g0197(.A(new_n389), .B1(new_n344), .B2(new_n390), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n396), .A2(new_n397), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT13), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n359), .A2(G232), .A3(G1698), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n359), .A2(G226), .A3(new_n282), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G97), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n293), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n366), .B1(G238), .B2(new_n367), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n402), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n407), .A2(new_n408), .A3(new_n402), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT14), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(new_n413), .A3(G169), .ZN(new_n414));
  INV_X1    g0214(.A(new_n411), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n415), .A2(new_n409), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(G179), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n413), .B1(new_n412), .B2(G169), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n401), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n412), .A2(G200), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n400), .B(new_n421), .C1(new_n373), .C2(new_n412), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n347), .A2(new_n349), .B1(G20), .B2(G77), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n222), .A2(KEYINPUT15), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT15), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(G87), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n348), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n309), .B1(new_n425), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n343), .A2(G77), .A3(new_n340), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(G77), .B2(new_n305), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  OAI22_X1  g0234(.A1(new_n361), .A2(new_n221), .B1(new_n228), .B2(new_n359), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n288), .A2(new_n243), .A3(G1698), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n293), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n366), .B1(G244), .B2(new_n367), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n434), .B1(new_n383), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n439), .ZN(new_n441));
  INV_X1    g0241(.A(G179), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n439), .A2(G200), .ZN(new_n446));
  AOI211_X1 g0246(.A(new_n431), .B(new_n433), .C1(new_n441), .C2(G190), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n381), .A2(new_n386), .A3(new_n424), .A4(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(G58), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n450), .A2(new_n220), .ZN(new_n451));
  OAI21_X1  g0251(.A(G20), .B1(new_n451), .B2(new_n201), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n349), .A2(G159), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n279), .A2(new_n281), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n207), .ZN(new_n457));
  OAI21_X1  g0257(.A(G68), .B1(new_n457), .B2(KEYINPUT7), .ZN(new_n458));
  AOI21_X1  g0258(.A(G20), .B1(new_n279), .B2(new_n281), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT7), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI211_X1 g0261(.A(KEYINPUT16), .B(new_n455), .C1(new_n458), .C2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT16), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n460), .A2(G20), .ZN(new_n464));
  AOI21_X1  g0264(.A(G33), .B1(new_n277), .B2(new_n278), .ZN(new_n465));
  INV_X1    g0265(.A(new_n287), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n460), .B1(new_n359), .B2(G20), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n220), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n463), .B1(new_n469), .B2(new_n454), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n462), .A2(new_n308), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n366), .B1(G232), .B2(new_n367), .ZN(new_n472));
  MUX2_X1   g0272(.A(G223), .B(G226), .S(G1698), .Z(new_n473));
  NAND3_X1  g0273(.A1(new_n473), .A2(new_n279), .A3(new_n281), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G87), .ZN(new_n475));
  AND2_X1   g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n472), .B(new_n335), .C1(new_n476), .C2(new_n272), .ZN(new_n477));
  INV_X1    g0277(.A(new_n366), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n367), .A2(G232), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n272), .B1(new_n474), .B2(new_n475), .ZN(new_n481));
  OAI21_X1  g0281(.A(G200), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n347), .A2(new_n340), .ZN(new_n484));
  OAI22_X1  g0284(.A1(new_n344), .A2(new_n484), .B1(new_n305), .B2(new_n347), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n471), .A2(new_n483), .A3(KEYINPUT75), .A4(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT17), .ZN(new_n488));
  XNOR2_X1  g0288(.A(new_n487), .B(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n471), .A2(new_n486), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n472), .B(G179), .C1(new_n476), .C2(new_n272), .ZN(new_n491));
  OAI21_X1  g0291(.A(G169), .B1(new_n480), .B2(new_n481), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(KEYINPUT18), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n490), .A2(new_n493), .A3(KEYINPUT18), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n494), .B1(new_n495), .B2(KEYINPUT73), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n490), .A2(new_n493), .A3(KEYINPUT18), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT73), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n489), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n449), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT79), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n306), .A2(new_n300), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n504), .B1(new_n311), .B2(new_n300), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT6), .ZN(new_n506));
  AND2_X1   g0306(.A1(G97), .A2(G107), .ZN(new_n507));
  NOR2_X1   g0307(.A1(G97), .A2(G107), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT76), .ZN(new_n510));
  NAND2_X1  g0310(.A1(KEYINPUT6), .A2(G97), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n510), .B1(new_n511), .B2(G107), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n228), .A2(KEYINPUT76), .A3(KEYINPUT6), .A4(G97), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n509), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G20), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n393), .A2(new_n226), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n228), .B1(new_n467), .B2(new_n468), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n308), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT77), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n464), .ZN(new_n523));
  AND2_X1   g0323(.A1(KEYINPUT72), .A2(KEYINPUT3), .ZN(new_n524));
  NOR2_X1   g0324(.A1(KEYINPUT72), .A2(KEYINPUT3), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n280), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n523), .B1(new_n526), .B2(new_n287), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT7), .B1(new_n288), .B2(new_n207), .ZN(new_n528));
  OAI21_X1  g0328(.A(G107), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n516), .B1(new_n514), .B2(G20), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n531), .A2(KEYINPUT77), .A3(new_n308), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n505), .B1(new_n522), .B2(new_n532), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n279), .A2(G244), .A3(new_n282), .A4(new_n281), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT4), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AND2_X1   g0336(.A1(KEYINPUT4), .A2(G244), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n281), .A2(new_n287), .A3(new_n537), .A4(new_n282), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n281), .A2(new_n287), .A3(G250), .A4(G1698), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n538), .A2(new_n539), .A3(new_n299), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n272), .B1(new_n536), .B2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n272), .B(G257), .C1(new_n256), .C2(new_n264), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n270), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n383), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n543), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n538), .A2(new_n539), .A3(new_n299), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n546), .B1(new_n535), .B2(new_n534), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n545), .B(new_n442), .C1(new_n547), .C2(new_n272), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n503), .B1(new_n533), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n505), .ZN(new_n551));
  AOI21_X1  g0351(.A(KEYINPUT77), .B1(new_n531), .B2(new_n308), .ZN(new_n552));
  AOI211_X1 g0352(.A(new_n521), .B(new_n309), .C1(new_n529), .C2(new_n530), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n544), .A2(new_n548), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n554), .A2(new_n555), .A3(KEYINPUT79), .ZN(new_n556));
  OAI21_X1  g0356(.A(G200), .B1(new_n541), .B2(new_n543), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n545), .B(G190), .C1(new_n547), .C2(new_n272), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n533), .A2(new_n559), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n550), .A2(new_n556), .A3(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(G238), .A2(G1698), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n562), .B1(new_n227), .B2(G1698), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n563), .A2(new_n279), .A3(new_n281), .ZN(new_n564));
  NAND2_X1  g0364(.A1(G33), .A2(G116), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n272), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n260), .A2(G250), .ZN(new_n567));
  NOR3_X1   g0367(.A1(new_n259), .A2(G1), .A3(G274), .ZN(new_n568));
  NOR3_X1   g0368(.A1(new_n567), .A2(new_n293), .A3(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n442), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n429), .A2(new_n305), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT19), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n348), .A2(new_n573), .A3(G97), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n508), .A2(new_n222), .B1(new_n405), .B2(new_n207), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n574), .B1(new_n575), .B2(new_n573), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n279), .A2(new_n207), .A3(G68), .A4(new_n281), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n572), .B1(new_n578), .B2(new_n308), .ZN(new_n579));
  INV_X1    g0379(.A(new_n311), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n429), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n383), .B1(new_n566), .B2(new_n569), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n571), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(G200), .B1(new_n566), .B2(new_n569), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n580), .A2(G87), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n579), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n570), .A2(G190), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n584), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  MUX2_X1   g0391(.A(G250), .B(G257), .S(G1698), .Z(new_n592));
  NAND3_X1  g0392(.A1(new_n592), .A2(new_n279), .A3(new_n281), .ZN(new_n593));
  NAND2_X1  g0393(.A1(G33), .A2(G294), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n272), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AND4_X1   g0395(.A1(new_n265), .A2(new_n258), .A3(new_n269), .A4(new_n263), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n272), .B(G264), .C1(new_n256), .C2(new_n264), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NOR4_X1   g0398(.A1(new_n595), .A2(new_n596), .A3(G179), .A4(new_n598), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n595), .A2(new_n596), .A3(new_n598), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n599), .B1(new_n601), .B2(new_n383), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT83), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT22), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n604), .A2(new_n207), .A3(G87), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n288), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  NOR3_X1   g0406(.A1(new_n222), .A2(KEYINPUT22), .A3(G20), .ZN(new_n607));
  AOI21_X1  g0407(.A(KEYINPUT83), .B1(new_n359), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n279), .A2(new_n207), .A3(G87), .A4(new_n281), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(KEYINPUT22), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n228), .A2(KEYINPUT23), .A3(G20), .ZN(new_n613));
  AOI21_X1  g0413(.A(KEYINPUT23), .B1(new_n228), .B2(G20), .ZN(new_n614));
  OAI22_X1  g0414(.A1(new_n613), .A2(new_n614), .B1(G20), .B2(new_n565), .ZN(new_n615));
  OAI21_X1  g0415(.A(KEYINPUT24), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n615), .B1(new_n609), .B2(new_n611), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT24), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n309), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n306), .A2(KEYINPUT25), .A3(new_n228), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT25), .B1(new_n306), .B2(new_n228), .ZN(new_n623));
  OAI22_X1  g0423(.A1(new_n622), .A2(new_n623), .B1(new_n311), .B2(new_n228), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n602), .B1(new_n620), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n600), .A2(new_n373), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n626), .B1(G200), .B2(new_n600), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n617), .A2(new_n618), .ZN(new_n628));
  AOI211_X1 g0428(.A(KEYINPUT24), .B(new_n615), .C1(new_n609), .C2(new_n611), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n308), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n624), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n627), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n591), .A2(new_n625), .A3(new_n632), .ZN(new_n633));
  AND4_X1   g0433(.A1(new_n339), .A2(new_n502), .A3(new_n561), .A4(new_n633), .ZN(G372));
  NOR2_X1   g0434(.A1(new_n495), .A2(new_n494), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n422), .A2(new_n445), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n420), .ZN(new_n637));
  XNOR2_X1  g0437(.A(new_n487), .B(KEYINPUT17), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n635), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n639), .A2(KEYINPUT85), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(KEYINPUT85), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(new_n381), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n386), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n502), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n554), .A2(new_n555), .A3(KEYINPUT79), .ZN(new_n646));
  AOI21_X1  g0446(.A(KEYINPUT79), .B1(new_n554), .B2(new_n555), .ZN(new_n647));
  OAI211_X1 g0447(.A(KEYINPUT26), .B(new_n591), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT26), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n571), .A2(new_n582), .A3(new_n583), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT84), .ZN(new_n651));
  INV_X1    g0451(.A(new_n588), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n651), .B1(new_n652), .B2(new_n585), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n585), .A2(new_n651), .A3(new_n579), .A4(new_n587), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n590), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n650), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n554), .A2(new_n555), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n649), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n648), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n653), .A2(new_n655), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n324), .A2(new_n326), .A3(new_n328), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n660), .B1(new_n661), .B2(new_n625), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n646), .A2(new_n647), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n560), .A2(new_n632), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n659), .A2(new_n665), .A3(new_n650), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n644), .B1(new_n645), .B2(new_n667), .ZN(G369));
  NAND3_X1  g0468(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(G213), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(G343), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n339), .B1(new_n330), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n324), .A2(new_n326), .A3(new_n328), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n677), .A2(new_n317), .A3(new_n674), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n678), .A2(KEYINPUT86), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(KEYINPUT86), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n676), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n681), .A2(G330), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n625), .A2(new_n632), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n674), .B1(new_n620), .B2(new_n624), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n625), .B2(new_n675), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n329), .A2(new_n675), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n683), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n600), .A2(new_n442), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(G169), .B2(new_n600), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(new_n630), .B2(new_n631), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n675), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n687), .A2(new_n694), .ZN(G399));
  AND2_X1   g0495(.A1(new_n654), .A2(new_n590), .ZN(new_n696));
  OAI21_X1  g0496(.A(KEYINPUT84), .B1(new_n586), .B2(new_n588), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n584), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n663), .A2(new_n664), .A3(new_n698), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n625), .A2(new_n319), .A3(new_n327), .A4(new_n328), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(KEYINPUT90), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n550), .A2(new_n556), .A3(new_n560), .A4(new_n632), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT90), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n704), .A2(new_n705), .A3(new_n698), .A4(new_n700), .ZN(new_n706));
  OAI211_X1 g0506(.A(new_n649), .B(new_n591), .C1(new_n646), .C2(new_n647), .ZN(new_n707));
  OAI21_X1  g0507(.A(KEYINPUT26), .B1(new_n656), .B2(new_n657), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n707), .A2(new_n650), .A3(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n702), .A2(new_n706), .A3(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(KEYINPUT29), .A3(new_n675), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n533), .A2(new_n549), .ZN(new_n712));
  AOI21_X1  g0512(.A(KEYINPUT26), .B1(new_n698), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n589), .A2(new_n590), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n650), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n715), .B1(new_n550), .B2(new_n556), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n713), .B1(KEYINPUT26), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n696), .A2(new_n697), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n692), .B2(new_n677), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n650), .B1(new_n703), .B2(new_n719), .ZN(new_n720));
  OAI211_X1 g0520(.A(KEYINPUT88), .B(new_n675), .C1(new_n717), .C2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(KEYINPUT88), .B1(new_n666), .B2(new_n675), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT29), .ZN(new_n725));
  AOI21_X1  g0525(.A(KEYINPUT89), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n675), .B1(new_n717), .B2(new_n720), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT88), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n729), .A2(KEYINPUT89), .A3(new_n725), .A4(new_n721), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n711), .B1(new_n726), .B2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT91), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n339), .A2(new_n561), .A3(new_n633), .A4(new_n675), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n536), .A2(new_n540), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n543), .B1(new_n735), .B2(new_n293), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n595), .A2(new_n598), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n316), .A2(new_n736), .A3(new_n570), .A4(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT30), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n600), .A2(new_n570), .A3(G179), .ZN(new_n741));
  INV_X1    g0541(.A(new_n736), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n741), .A2(new_n322), .A3(new_n742), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n737), .A2(new_n570), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n744), .A2(KEYINPUT30), .A3(new_n316), .A4(new_n736), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n740), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n746), .A2(KEYINPUT31), .A3(new_n674), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT31), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n743), .A2(new_n745), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n740), .A2(KEYINPUT87), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT87), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n738), .A2(new_n751), .A3(new_n739), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n749), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n748), .B1(new_n753), .B2(new_n675), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n734), .A2(new_n747), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G330), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n732), .A2(new_n733), .A3(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n711), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n729), .A2(new_n725), .A3(new_n721), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT89), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n758), .B1(new_n761), .B2(new_n730), .ZN(new_n762));
  INV_X1    g0562(.A(new_n756), .ZN(new_n763));
  OAI21_X1  g0563(.A(KEYINPUT91), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n757), .A2(new_n206), .A3(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n210), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G41), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n508), .A2(new_n222), .A3(new_n297), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n768), .A2(G1), .A3(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(new_n216), .B2(new_n768), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT28), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n765), .A2(new_n773), .ZN(G364));
  AND2_X1   g0574(.A1(new_n207), .A2(G13), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n206), .B1(new_n775), .B2(G45), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n767), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n682), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(G330), .B2(new_n681), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n210), .A2(new_n359), .ZN(new_n781));
  INV_X1    g0581(.A(G355), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n781), .A2(new_n782), .B1(G116), .B2(new_n210), .ZN(new_n783));
  INV_X1    g0583(.A(new_n456), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n766), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n786), .B1(new_n259), .B2(new_n217), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n250), .A2(new_n259), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n783), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G13), .A2(G33), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(G20), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n213), .B1(G20), .B2(new_n383), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n778), .B1(new_n789), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n207), .A2(G179), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n331), .A2(G190), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(G190), .A2(G200), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(G283), .A2(new_n800), .B1(new_n803), .B2(G329), .ZN(new_n804));
  INV_X1    g0604(.A(G303), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n797), .A2(G190), .A3(G200), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n804), .B(new_n288), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  NOR3_X1   g0607(.A1(new_n373), .A2(G179), .A3(G200), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n207), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n807), .B1(G294), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G311), .ZN(new_n812));
  NAND2_X1  g0612(.A1(G20), .A2(G179), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT92), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(new_n801), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n798), .ZN(new_n816));
  XOR2_X1   g0616(.A(KEYINPUT33), .B(G317), .Z(new_n817));
  OAI22_X1  g0617(.A1(new_n812), .A2(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n814), .A2(new_n331), .A3(new_n335), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n818), .B1(G322), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G326), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n814), .A2(G200), .A3(new_n335), .ZN(new_n823));
  XOR2_X1   g0623(.A(new_n823), .B(KEYINPUT94), .Z(new_n824));
  OAI211_X1 g0624(.A(new_n811), .B(new_n821), .C1(new_n822), .C2(new_n824), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n815), .A2(KEYINPUT93), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n815), .A2(KEYINPUT93), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(new_n226), .ZN(new_n829));
  INV_X1    g0629(.A(new_n823), .ZN(new_n830));
  AOI22_X1  g0630(.A1(G50), .A2(new_n830), .B1(new_n820), .B2(G58), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n806), .A2(new_n222), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n359), .B1(new_n799), .B2(new_n228), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n832), .B(new_n833), .C1(G97), .C2(new_n810), .ZN(new_n834));
  INV_X1    g0634(.A(new_n816), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n803), .A2(KEYINPUT32), .A3(G159), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT32), .ZN(new_n837));
  INV_X1    g0637(.A(G159), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n837), .B1(new_n802), .B2(new_n838), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n835), .A2(G68), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n831), .A2(new_n834), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n825), .B1(new_n829), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n796), .B1(new_n842), .B2(new_n793), .ZN(new_n843));
  INV_X1    g0643(.A(new_n792), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n843), .B1(new_n681), .B2(new_n844), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n780), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(G396));
  NOR2_X1   g0647(.A1(new_n444), .A2(new_n674), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n447), .A2(new_n446), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n434), .B2(new_n675), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n848), .B1(new_n850), .B2(new_n444), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n724), .A2(new_n852), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n675), .B(new_n851), .C1(new_n717), .C2(new_n720), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n778), .B1(new_n855), .B2(new_n756), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n756), .B2(new_n855), .ZN(new_n857));
  INV_X1    g0657(.A(new_n778), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n793), .A2(new_n790), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT95), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n858), .B1(new_n861), .B2(new_n226), .ZN(new_n862));
  INV_X1    g0662(.A(new_n806), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n863), .A2(G107), .B1(new_n803), .B2(G311), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n359), .B1(new_n800), .B2(G87), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n864), .B(new_n865), .C1(new_n300), .C2(new_n809), .ZN(new_n866));
  AOI22_X1  g0666(.A1(G294), .A2(new_n820), .B1(new_n830), .B2(G303), .ZN(new_n867));
  INV_X1    g0667(.A(G283), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n867), .B1(new_n868), .B2(new_n816), .ZN(new_n869));
  INV_X1    g0669(.A(new_n828), .ZN(new_n870));
  AOI211_X1 g0670(.A(new_n866), .B(new_n869), .C1(G116), .C2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n800), .A2(G68), .ZN(new_n872));
  INV_X1    g0672(.A(G132), .ZN(new_n873));
  OAI221_X1 g0673(.A(new_n872), .B1(new_n202), .B2(new_n806), .C1(new_n873), .C2(new_n802), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n784), .B1(new_n450), .B2(new_n809), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n820), .A2(G143), .B1(new_n835), .B2(G150), .ZN(new_n876));
  INV_X1    g0676(.A(G137), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n876), .B1(new_n877), .B2(new_n823), .C1(new_n828), .C2(new_n838), .ZN(new_n878));
  XOR2_X1   g0678(.A(KEYINPUT96), .B(KEYINPUT34), .Z(new_n879));
  XNOR2_X1  g0679(.A(new_n878), .B(new_n879), .ZN(new_n880));
  AOI211_X1 g0680(.A(new_n874), .B(new_n875), .C1(new_n880), .C2(KEYINPUT97), .ZN(new_n881));
  OR2_X1    g0681(.A1(new_n880), .A2(KEYINPUT97), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n871), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n793), .ZN(new_n884));
  OAI221_X1 g0684(.A(new_n862), .B1(new_n791), .B2(new_n851), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n857), .A2(new_n885), .ZN(G384));
  OR2_X1    g0686(.A1(new_n514), .A2(KEYINPUT35), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n514), .A2(KEYINPUT35), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n887), .A2(G116), .A3(new_n214), .A4(new_n888), .ZN(new_n889));
  XOR2_X1   g0689(.A(new_n889), .B(KEYINPUT36), .Z(new_n890));
  OR3_X1    g0690(.A1(new_n216), .A2(new_n226), .A3(new_n451), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n202), .A2(G68), .ZN(new_n892));
  AOI211_X1 g0692(.A(new_n206), .B(G13), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n711), .A2(new_n502), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n895), .B1(new_n761), .B2(new_n730), .ZN(new_n896));
  OR2_X1    g0696(.A1(new_n896), .A2(new_n643), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n471), .A2(new_n483), .A3(new_n486), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n457), .A2(KEYINPUT7), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n220), .B1(new_n459), .B2(new_n460), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n454), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n309), .B1(new_n901), .B2(KEYINPUT16), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n455), .B1(new_n458), .B2(new_n461), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n463), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n485), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n898), .B1(new_n905), .B2(new_n672), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n491), .A2(new_n492), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT37), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n490), .A2(new_n493), .ZN(new_n910));
  INV_X1    g0710(.A(new_n672), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n490), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT37), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n910), .A2(new_n912), .A3(new_n913), .A4(new_n898), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n909), .A2(new_n914), .ZN(new_n915));
  OR2_X1    g0715(.A1(new_n905), .A2(new_n672), .ZN(new_n916));
  OAI211_X1 g0716(.A(KEYINPUT38), .B(new_n915), .C1(new_n500), .C2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT38), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n490), .A2(KEYINPUT73), .A3(KEYINPUT18), .A4(new_n493), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT18), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n910), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n499), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n916), .B1(new_n922), .B2(new_n638), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n909), .A2(new_n914), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n918), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n917), .A2(new_n925), .A3(KEYINPUT39), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n910), .A2(new_n912), .A3(new_n898), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(KEYINPUT37), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n914), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n921), .A2(new_n497), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n912), .B1(new_n638), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n918), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(KEYINPUT39), .B1(new_n917), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n926), .A2(new_n934), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n418), .A2(new_n419), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n936), .A2(new_n401), .A3(new_n675), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n400), .A2(new_n675), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n423), .A2(new_n940), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n420), .B(new_n422), .C1(new_n400), .C2(new_n675), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n848), .B(KEYINPUT98), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n944), .B1(new_n854), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n917), .A2(new_n925), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n946), .A2(new_n947), .B1(new_n635), .B2(new_n672), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n939), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n897), .B(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n754), .A2(KEYINPUT99), .ZN(new_n951));
  OR3_X1    g0751(.A1(new_n753), .A2(new_n748), .A3(new_n675), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT99), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n953), .B(new_n748), .C1(new_n753), .C2(new_n675), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n951), .A2(new_n734), .A3(new_n952), .A4(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n852), .B1(new_n942), .B2(new_n941), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(KEYINPUT100), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT40), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(new_n917), .B2(new_n933), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT100), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n955), .A2(new_n956), .A3(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n958), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n917), .A2(new_n925), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n959), .B1(new_n964), .B2(new_n957), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n502), .A2(new_n955), .ZN(new_n967));
  OAI21_X1  g0767(.A(G330), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(new_n966), .B2(new_n967), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n950), .A2(new_n969), .B1(new_n206), .B2(new_n775), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n950), .A2(new_n969), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n894), .B1(new_n970), .B2(new_n971), .ZN(G367));
  INV_X1    g0772(.A(new_n429), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n794), .B1(new_n210), .B2(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(new_n241), .B2(new_n785), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n824), .A2(new_n812), .B1(new_n868), .B2(new_n828), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT46), .ZN(new_n977));
  NOR3_X1   g0777(.A1(new_n806), .A2(new_n977), .A3(new_n297), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n977), .B1(new_n806), .B2(new_n297), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n228), .B2(new_n809), .ZN(new_n980));
  INV_X1    g0780(.A(G317), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n799), .A2(new_n300), .B1(new_n802), .B2(new_n981), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n784), .B(new_n982), .C1(new_n835), .C2(G294), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n805), .B2(new_n819), .ZN(new_n984));
  NOR4_X1   g0784(.A1(new_n976), .A2(new_n978), .A3(new_n980), .A4(new_n984), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT105), .ZN(new_n986));
  INV_X1    g0786(.A(G150), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n819), .A2(new_n987), .B1(new_n816), .B2(new_n838), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n809), .A2(new_n220), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n359), .B1(new_n799), .B2(new_n226), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n806), .A2(new_n450), .B1(new_n802), .B2(new_n877), .ZN(new_n991));
  NOR4_X1   g0791(.A1(new_n988), .A2(new_n989), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(G143), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n992), .B1(new_n202), .B2(new_n828), .C1(new_n993), .C2(new_n824), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n986), .A2(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(KEYINPUT106), .B(KEYINPUT47), .Z(new_n996));
  XNOR2_X1  g0796(.A(new_n995), .B(new_n996), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n858), .B(new_n975), .C1(new_n997), .C2(new_n793), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n588), .A2(new_n674), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n584), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(new_n656), .B2(new_n999), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT101), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n998), .B1(new_n844), .B2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT107), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT44), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n561), .B1(new_n533), .B2(new_n675), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n712), .A2(new_n674), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1005), .B1(new_n694), .B2(new_n1008), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n689), .A2(new_n693), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1010), .A2(new_n1011), .A3(KEYINPUT44), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1009), .A2(KEYINPUT104), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(KEYINPUT44), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT104), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n694), .A2(KEYINPUT45), .A3(new_n1008), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT45), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  AND4_X1   g0820(.A1(new_n687), .A2(new_n1013), .A3(new_n1016), .A4(new_n1020), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1019), .A2(new_n1017), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n687), .B1(new_n1022), .B2(new_n1013), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n689), .B1(new_n686), .B2(new_n688), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n682), .B(new_n1025), .Z(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n757), .A2(new_n764), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n767), .B(KEYINPUT41), .Z(new_n1029));
  OAI21_X1  g0829(.A(new_n776), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OR3_X1    g0830(.A1(new_n1010), .A2(KEYINPUT42), .A3(new_n689), .ZN(new_n1031));
  OAI21_X1  g0831(.A(KEYINPUT42), .B1(new_n1010), .B2(new_n689), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n647), .B(new_n646), .C1(new_n1008), .C2(new_n692), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1031), .B(new_n1032), .C1(new_n674), .C2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1002), .A2(KEYINPUT43), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT102), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n687), .A2(new_n1010), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n1002), .A2(KEYINPUT43), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT103), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AND3_X1   g0841(.A1(new_n1037), .A2(new_n1038), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1038), .B1(new_n1037), .B2(new_n1041), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n1042), .A2(new_n1043), .B1(new_n1040), .B2(new_n1039), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1037), .A2(new_n1041), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1038), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1037), .A2(new_n1038), .A3(new_n1041), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  AND2_X1   g0850(.A1(new_n1044), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1004), .B1(new_n1030), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(G387));
  AOI21_X1  g0853(.A(new_n733), .B1(new_n732), .B2(new_n756), .ZN(new_n1054));
  NOR3_X1   g0854(.A1(new_n762), .A2(KEYINPUT91), .A3(new_n763), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1027), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT112), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n767), .B(KEYINPUT111), .Z(new_n1058));
  NAND3_X1  g0858(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1026), .B1(new_n757), .B2(new_n764), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1058), .ZN(new_n1061));
  OAI21_X1  g0861(.A(KEYINPUT112), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n757), .A2(new_n764), .A3(new_n1026), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1059), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n820), .A2(G317), .B1(new_n835), .B2(G311), .ZN(new_n1065));
  INV_X1    g0865(.A(G322), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1065), .B1(new_n828), .B2(new_n805), .C1(new_n824), .C2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT48), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n810), .A2(G283), .B1(new_n863), .B2(G294), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT49), .Z(new_n1073));
  OAI221_X1 g0873(.A(new_n456), .B1(new_n297), .B2(new_n799), .C1(new_n822), .C2(new_n802), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT110), .Z(new_n1075));
  NOR2_X1   g0875(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n830), .A2(G159), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT109), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(G97), .A2(new_n800), .B1(new_n803), .B2(G150), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n226), .B2(new_n806), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n809), .A2(new_n973), .ZN(new_n1081));
  NOR3_X1   g0881(.A1(new_n1080), .A2(new_n456), .A3(new_n1081), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n220), .A2(new_n815), .B1(new_n816), .B2(new_n346), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(G50), .B2(new_n820), .ZN(new_n1084));
  AND3_X1   g0884(.A1(new_n1078), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n793), .B1(new_n1076), .B2(new_n1085), .ZN(new_n1086));
  OR2_X1    g0886(.A1(new_n686), .A2(new_n844), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n781), .A2(new_n770), .B1(G107), .B2(new_n210), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n246), .A2(G45), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n346), .A2(G50), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT50), .ZN(new_n1091));
  AOI211_X1 g0891(.A(G45), .B(new_n769), .C1(G68), .C2(G77), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n786), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1088), .B1(new_n1089), .B2(new_n1093), .ZN(new_n1094));
  OR2_X1    g0894(.A1(new_n1094), .A2(KEYINPUT108), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n795), .B1(new_n1094), .B2(KEYINPUT108), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n858), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n1086), .A2(new_n1087), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n1027), .B2(new_n777), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1064), .A2(new_n1099), .ZN(G393));
  OAI221_X1 g0900(.A(new_n794), .B1(new_n300), .B2(new_n210), .C1(new_n786), .C2(new_n253), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n778), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(G68), .A2(new_n863), .B1(new_n800), .B2(G87), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1103), .B(new_n784), .C1(new_n993), .C2(new_n802), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT113), .Z(new_n1105));
  AOI22_X1  g0905(.A1(new_n835), .A2(G50), .B1(G77), .B2(new_n810), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1105), .B(new_n1106), .C1(new_n346), .C2(new_n828), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n987), .A2(new_n823), .B1(new_n819), .B2(new_n838), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT51), .Z(new_n1109));
  OAI22_X1  g0909(.A1(new_n812), .A2(new_n819), .B1(new_n823), .B2(new_n981), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT52), .Z(new_n1111));
  AOI22_X1  g0911(.A1(new_n863), .A2(G283), .B1(new_n803), .B2(G322), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1112), .B(new_n288), .C1(new_n228), .C2(new_n799), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n809), .A2(new_n297), .ZN(new_n1114));
  INV_X1    g0914(.A(G294), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n1115), .A2(new_n815), .B1(new_n816), .B2(new_n805), .ZN(new_n1116));
  OR3_X1    g0916(.A1(new_n1113), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n1107), .A2(new_n1109), .B1(new_n1111), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1102), .B1(new_n1118), .B2(new_n793), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n1008), .B2(new_n844), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1024), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1120), .B1(new_n1121), .B2(new_n776), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1061), .B1(new_n1060), .B2(new_n1024), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1056), .A2(new_n1121), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1122), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(G390));
  NAND2_X1  g0926(.A1(new_n955), .A2(G330), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n645), .A2(new_n1127), .ZN(new_n1128));
  NOR3_X1   g0928(.A1(new_n896), .A2(new_n643), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1127), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n755), .A2(G330), .A3(new_n851), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1130), .A2(new_n956), .B1(new_n944), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n854), .A2(new_n945), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n943), .B1(new_n1130), .B2(new_n851), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n710), .A2(new_n675), .A3(new_n851), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n755), .A2(G330), .A3(new_n851), .A4(new_n943), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1136), .A2(new_n1137), .A3(new_n945), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n1132), .A2(new_n1134), .B1(new_n1135), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1129), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1130), .A2(new_n956), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NOR3_X1   g0942(.A1(new_n923), .A2(new_n924), .A3(new_n918), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n490), .B(new_n911), .C1(new_n489), .C2(new_n635), .ZN(new_n1144));
  AOI21_X1  g0944(.A(KEYINPUT38), .B1(new_n1144), .B2(new_n929), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n937), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1136), .A2(new_n945), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1146), .B1(new_n1147), .B2(new_n943), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1133), .A2(new_n943), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT39), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n917), .A2(new_n925), .A3(KEYINPUT39), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n937), .A2(new_n1149), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1142), .B1(new_n1148), .B2(new_n1153), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n926), .A2(new_n934), .B1(new_n946), .B2(new_n938), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n944), .B1(new_n1136), .B2(new_n945), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1155), .B(new_n1137), .C1(new_n1156), .C2(new_n1146), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1140), .A2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1129), .A2(new_n1139), .A3(new_n1157), .A4(new_n1154), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1159), .A2(new_n1058), .A3(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1154), .A2(new_n1157), .A3(new_n777), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n858), .B1(new_n861), .B2(new_n346), .ZN(new_n1163));
  INV_X1    g0963(.A(G125), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n359), .B1(new_n802), .B2(new_n1164), .C1(new_n202), .C2(new_n799), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n806), .A2(new_n987), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT114), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1167), .A2(KEYINPUT53), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n1165), .B(new_n1168), .C1(G159), .C2(new_n810), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1167), .A2(KEYINPUT53), .ZN(new_n1170));
  XOR2_X1   g0970(.A(KEYINPUT54), .B(G143), .Z(new_n1171));
  NAND2_X1  g0971(.A1(new_n870), .A2(new_n1171), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n819), .A2(new_n873), .B1(new_n816), .B2(new_n877), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G128), .B2(new_n830), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1169), .A2(new_n1170), .A3(new_n1172), .A4(new_n1174), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n823), .A2(new_n868), .B1(new_n816), .B2(new_n228), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(G116), .B2(new_n820), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n872), .B1(new_n1115), .B2(new_n802), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n809), .A2(new_n226), .ZN(new_n1179));
  NOR4_X1   g0979(.A1(new_n1178), .A2(new_n359), .A3(new_n832), .A4(new_n1179), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1177), .B(new_n1180), .C1(new_n300), .C2(new_n828), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT115), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1175), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1163), .B1(new_n884), .B2(new_n1185), .C1(new_n935), .C2(new_n791), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1162), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT116), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1162), .A2(KEYINPUT116), .A3(new_n1186), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1189), .A2(KEYINPUT117), .A3(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(KEYINPUT117), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1161), .B1(new_n1192), .B2(new_n1193), .ZN(G378));
  NAND3_X1  g0994(.A1(new_n963), .A2(G330), .A3(new_n965), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n381), .A2(new_n386), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n357), .A2(new_n672), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1197), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1202), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1204), .A2(new_n1200), .A3(new_n1196), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1195), .A2(new_n1207), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1206), .A2(new_n963), .A3(G330), .A4(new_n965), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n949), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1208), .A2(new_n949), .A3(new_n1209), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1207), .A2(new_n790), .ZN(new_n1215));
  NOR3_X1   g1015(.A1(new_n793), .A2(G50), .A3(new_n790), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n784), .A2(G41), .ZN(new_n1217));
  AOI211_X1 g1017(.A(G50), .B(new_n1217), .C1(new_n280), .C2(new_n255), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n806), .A2(new_n226), .B1(new_n802), .B2(new_n868), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n989), .B(new_n1219), .C1(new_n835), .C2(G97), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1220), .B(new_n1217), .C1(new_n297), .C2(new_n823), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n799), .A2(new_n450), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT118), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1223), .B1(new_n228), .B2(new_n819), .C1(new_n973), .C2(new_n815), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1221), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  XOR2_X1   g1026(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n1227));
  AOI21_X1  g1027(.A(new_n1218), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(G128), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n1164), .A2(new_n823), .B1(new_n819), .B2(new_n1229), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n810), .A2(G150), .B1(new_n863), .B2(new_n1171), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n877), .B2(new_n815), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n1230), .B(new_n1232), .C1(G132), .C2(new_n835), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1234), .A2(KEYINPUT59), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n280), .B(new_n255), .C1(new_n799), .C2(new_n838), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(G124), .B2(new_n803), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT59), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1237), .B1(new_n1233), .B2(new_n1238), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1228), .B1(new_n1235), .B2(new_n1239), .C1(new_n1227), .C2(new_n1226), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n858), .B(new_n1216), .C1(new_n1240), .C2(new_n793), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n1214), .A2(new_n777), .B1(new_n1215), .B2(new_n1241), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n1213), .A2(new_n1212), .B1(new_n1160), .B2(new_n1129), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1058), .B1(new_n1243), .B2(KEYINPUT57), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1131), .A2(new_n944), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1134), .B1(new_n1141), .B2(new_n1246), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1245), .A2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1129), .B1(new_n1158), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(KEYINPUT57), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1208), .A2(new_n949), .A3(new_n1209), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n949), .B1(new_n1209), .B2(new_n1208), .ZN(new_n1252));
  OAI21_X1  g1052(.A(KEYINPUT120), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT120), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1213), .A2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1250), .B1(new_n1253), .B2(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1242), .B1(new_n1244), .B2(new_n1256), .ZN(G375));
  XOR2_X1   g1057(.A(new_n776), .B(KEYINPUT121), .Z(new_n1258));
  OAI21_X1  g1058(.A(KEYINPUT122), .B1(new_n1248), .B2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n858), .B1(new_n861), .B2(new_n220), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n806), .A2(new_n838), .B1(new_n802), .B2(new_n1229), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n456), .B(new_n1261), .C1(G50), .C2(new_n810), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1262), .B(new_n1223), .C1(new_n987), .C2(new_n815), .ZN(new_n1263));
  XOR2_X1   g1063(.A(new_n1263), .B(KEYINPUT123), .Z(new_n1264));
  AOI22_X1  g1064(.A1(new_n830), .A2(G132), .B1(new_n835), .B2(new_n1171), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1264), .B(new_n1265), .C1(new_n877), .C2(new_n819), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n823), .A2(new_n1115), .B1(new_n816), .B2(new_n297), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(G283), .B2(new_n820), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n806), .A2(new_n300), .B1(new_n802), .B2(new_n805), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n288), .B1(new_n799), .B2(new_n226), .ZN(new_n1270));
  NOR3_X1   g1070(.A1(new_n1081), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1268), .B(new_n1271), .C1(new_n228), .C2(new_n828), .ZN(new_n1272));
  AND2_X1   g1072(.A1(new_n1266), .A2(new_n1272), .ZN(new_n1273));
  OAI221_X1 g1073(.A(new_n1260), .B1(new_n1273), .B2(new_n884), .C1(new_n943), .C2(new_n791), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1259), .A2(new_n1274), .ZN(new_n1275));
  NOR3_X1   g1075(.A1(new_n1248), .A2(KEYINPUT122), .A3(new_n1258), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1029), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1140), .A2(new_n1278), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1129), .A2(new_n1139), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1277), .B1(new_n1279), .B2(new_n1280), .ZN(G381));
  NAND3_X1  g1081(.A1(new_n1064), .A2(new_n846), .A3(new_n1099), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(G375), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1161), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NOR3_X1   g1086(.A1(G390), .A2(G381), .A3(G384), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1283), .A2(new_n1052), .A3(new_n1286), .A4(new_n1287), .ZN(G407));
  NAND2_X1  g1088(.A1(new_n1214), .A2(new_n777), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1215), .A2(new_n1241), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1253), .A2(new_n1255), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT57), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1293), .B1(new_n1160), .B2(new_n1129), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1292), .A2(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1249), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1061), .B1(new_n1296), .B2(new_n1293), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1291), .B1(new_n1295), .B2(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1298), .A2(new_n673), .A3(new_n1286), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(G407), .A2(G213), .A3(new_n1299), .ZN(G409));
  OAI21_X1  g1100(.A(new_n1290), .B1(new_n1296), .B2(new_n1029), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1258), .B1(new_n1253), .B2(new_n1255), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1286), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT117), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1285), .A2(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1284), .B1(new_n1305), .B2(new_n1191), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1303), .B1(G375), .B2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(KEYINPUT124), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n673), .A2(G213), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1280), .A2(KEYINPUT60), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT60), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1311), .B1(new_n1129), .B2(new_n1139), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1310), .A2(new_n1058), .A3(new_n1140), .A4(new_n1312), .ZN(new_n1313));
  AND3_X1   g1113(.A1(new_n1313), .A2(new_n1277), .A3(G384), .ZN(new_n1314));
  AOI21_X1  g1114(.A(G384), .B1(new_n1313), .B2(new_n1277), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT124), .ZN(new_n1317));
  OAI211_X1 g1117(.A(new_n1303), .B(new_n1317), .C1(G375), .C2(new_n1306), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1308), .A2(new_n1309), .A3(new_n1316), .A4(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT63), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT125), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1064), .A2(new_n846), .A3(new_n1099), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n846), .B1(new_n1064), .B2(new_n1099), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1322), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(G393), .A2(G396), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1326), .A2(KEYINPUT125), .A3(new_n1282), .ZN(new_n1327));
  XNOR2_X1  g1127(.A(new_n1052), .B(new_n1125), .ZN(new_n1328));
  AND3_X1   g1128(.A1(new_n1325), .A2(new_n1327), .A3(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1328), .B1(new_n1325), .B2(new_n1327), .ZN(new_n1330));
  NOR3_X1   g1130(.A1(new_n1329), .A2(new_n1330), .A3(KEYINPUT61), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1308), .A2(new_n1309), .A3(new_n1318), .ZN(new_n1332));
  INV_X1    g1132(.A(G2897), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1309), .A2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1316), .A2(new_n1334), .ZN(new_n1335));
  OAI22_X1  g1135(.A1(new_n1314), .A2(new_n1315), .B1(new_n1333), .B2(new_n1309), .ZN(new_n1336));
  AND2_X1   g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1332), .A2(new_n1338), .ZN(new_n1339));
  AND2_X1   g1139(.A1(new_n1307), .A2(new_n1309), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1340), .A2(KEYINPUT63), .A3(new_n1316), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1321), .A2(new_n1331), .A3(new_n1339), .A4(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT61), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1343), .B1(new_n1340), .B2(new_n1337), .ZN(new_n1344));
  XNOR2_X1  g1144(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1319), .A2(new_n1345), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1340), .A2(KEYINPUT62), .A3(new_n1316), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1344), .B1(new_n1346), .B2(new_n1347), .ZN(new_n1348));
  NOR2_X1   g1148(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1342), .B1(new_n1348), .B2(new_n1349), .ZN(G405));
  INV_X1    g1150(.A(KEYINPUT127), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1298), .A2(G378), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(G375), .A2(new_n1286), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1352), .A2(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1354), .A2(new_n1316), .ZN(new_n1355));
  INV_X1    g1155(.A(new_n1316), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1352), .A2(new_n1353), .A3(new_n1356), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1355), .A2(new_n1357), .ZN(new_n1358));
  AND3_X1   g1158(.A1(new_n1349), .A2(new_n1351), .A3(new_n1358), .ZN(new_n1359));
  AOI21_X1  g1159(.A(new_n1351), .B1(new_n1349), .B2(new_n1358), .ZN(new_n1360));
  NOR2_X1   g1160(.A1(new_n1349), .A2(new_n1358), .ZN(new_n1361));
  NOR3_X1   g1161(.A1(new_n1359), .A2(new_n1360), .A3(new_n1361), .ZN(G402));
endmodule


