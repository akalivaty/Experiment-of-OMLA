

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U556 ( .A1(n656), .A2(n542), .ZN(n674) );
  XNOR2_X1 U557 ( .A(n747), .B(KEYINPUT31), .ZN(n748) );
  NAND2_X1 U558 ( .A1(n522), .A2(n523), .ZN(n747) );
  NOR2_X1 U559 ( .A1(n726), .A2(n725), .ZN(n729) );
  XNOR2_X1 U560 ( .A(n758), .B(n757), .ZN(n786) );
  OR2_X1 U561 ( .A1(n765), .A2(n764), .ZN(n787) );
  AND2_X1 U562 ( .A1(G40), .A2(G160), .ZN(n709) );
  NOR2_X1 U563 ( .A1(n602), .A2(n601), .ZN(n603) );
  OR2_X1 U564 ( .A1(G168), .A2(n745), .ZN(n522) );
  OR2_X1 U565 ( .A1(G171), .A2(n746), .ZN(n523) );
  OR2_X1 U566 ( .A1(n778), .A2(n777), .ZN(n524) );
  OR2_X1 U567 ( .A1(n791), .A2(n784), .ZN(n525) );
  AND2_X1 U568 ( .A1(n525), .A2(n1005), .ZN(n526) );
  INV_X1 U569 ( .A(G8), .ZN(n742) );
  OR2_X1 U570 ( .A1(n761), .A2(n742), .ZN(n743) );
  INV_X1 U571 ( .A(n750), .ZN(n736) );
  INV_X1 U572 ( .A(KEYINPUT28), .ZN(n730) );
  XNOR2_X1 U573 ( .A(n731), .B(n730), .ZN(n732) );
  INV_X1 U574 ( .A(KEYINPUT29), .ZN(n734) );
  XNOR2_X1 U575 ( .A(n735), .B(n734), .ZN(n741) );
  INV_X1 U576 ( .A(KEYINPUT64), .ZN(n775) );
  NAND2_X1 U577 ( .A1(n810), .A2(n709), .ZN(n750) );
  INV_X1 U578 ( .A(KEYINPUT71), .ZN(n592) );
  NAND2_X1 U579 ( .A1(G8), .A2(n750), .ZN(n791) );
  XNOR2_X1 U580 ( .A(n593), .B(n592), .ZN(n596) );
  INV_X1 U581 ( .A(KEYINPUT17), .ZN(n527) );
  NAND2_X1 U582 ( .A1(n903), .A2(G137), .ZN(n530) );
  NOR2_X2 U583 ( .A1(G651), .A2(n656), .ZN(n667) );
  INV_X1 U584 ( .A(G651), .ZN(n542) );
  INV_X1 U585 ( .A(n717), .ZN(n984) );
  XNOR2_X1 U586 ( .A(n614), .B(n613), .ZN(n717) );
  XNOR2_X1 U587 ( .A(n603), .B(KEYINPUT72), .ZN(n989) );
  NOR2_X1 U588 ( .A1(G2105), .A2(G2104), .ZN(n528) );
  XNOR2_X2 U589 ( .A(n528), .B(n527), .ZN(n903) );
  INV_X1 U590 ( .A(G2104), .ZN(n568) );
  AND2_X1 U591 ( .A1(G2105), .A2(G2104), .ZN(n898) );
  NAND2_X1 U592 ( .A1(G113), .A2(n898), .ZN(n529) );
  NAND2_X1 U593 ( .A1(n530), .A2(n529), .ZN(n531) );
  OR2_X1 U594 ( .A1(n531), .A2(KEYINPUT65), .ZN(n533) );
  NAND2_X1 U595 ( .A1(n531), .A2(KEYINPUT65), .ZN(n532) );
  NAND2_X1 U596 ( .A1(n533), .A2(n532), .ZN(n539) );
  AND2_X1 U597 ( .A1(n568), .A2(G2105), .ZN(n896) );
  AND2_X1 U598 ( .A1(G125), .A2(n896), .ZN(n537) );
  INV_X1 U599 ( .A(G2105), .ZN(n534) );
  AND2_X1 U600 ( .A1(n534), .A2(G2104), .ZN(n904) );
  NAND2_X1 U601 ( .A1(G101), .A2(n904), .ZN(n535) );
  XNOR2_X1 U602 ( .A(KEYINPUT23), .B(n535), .ZN(n536) );
  NOR2_X1 U603 ( .A1(n537), .A2(n536), .ZN(n538) );
  AND2_X1 U604 ( .A1(n539), .A2(n538), .ZN(G160) );
  NOR2_X1 U605 ( .A1(G651), .A2(G543), .ZN(n673) );
  NAND2_X1 U606 ( .A1(G85), .A2(n673), .ZN(n541) );
  XOR2_X1 U607 ( .A(G543), .B(KEYINPUT0), .Z(n656) );
  NAND2_X1 U608 ( .A1(G72), .A2(n674), .ZN(n540) );
  NAND2_X1 U609 ( .A1(n541), .A2(n540), .ZN(n548) );
  NAND2_X1 U610 ( .A1(G47), .A2(n667), .ZN(n546) );
  NOR2_X1 U611 ( .A1(G543), .A2(n542), .ZN(n543) );
  XOR2_X1 U612 ( .A(KEYINPUT66), .B(n543), .Z(n544) );
  XNOR2_X2 U613 ( .A(KEYINPUT1), .B(n544), .ZN(n669) );
  NAND2_X1 U614 ( .A1(G60), .A2(n669), .ZN(n545) );
  NAND2_X1 U615 ( .A1(n546), .A2(n545), .ZN(n547) );
  OR2_X1 U616 ( .A1(n548), .A2(n547), .ZN(G290) );
  NAND2_X1 U617 ( .A1(G52), .A2(n667), .ZN(n550) );
  NAND2_X1 U618 ( .A1(G64), .A2(n669), .ZN(n549) );
  NAND2_X1 U619 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U620 ( .A(KEYINPUT67), .B(n551), .Z(n556) );
  NAND2_X1 U621 ( .A1(G90), .A2(n673), .ZN(n553) );
  NAND2_X1 U622 ( .A1(G77), .A2(n674), .ZN(n552) );
  NAND2_X1 U623 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U624 ( .A(KEYINPUT9), .B(n554), .Z(n555) );
  NOR2_X1 U625 ( .A1(n556), .A2(n555), .ZN(G171) );
  XOR2_X1 U626 ( .A(G2443), .B(G2446), .Z(n558) );
  XNOR2_X1 U627 ( .A(G2427), .B(G2451), .ZN(n557) );
  XNOR2_X1 U628 ( .A(n558), .B(n557), .ZN(n564) );
  XOR2_X1 U629 ( .A(G2430), .B(G2454), .Z(n560) );
  XNOR2_X1 U630 ( .A(G1348), .B(G1341), .ZN(n559) );
  XNOR2_X1 U631 ( .A(n560), .B(n559), .ZN(n562) );
  XOR2_X1 U632 ( .A(G2435), .B(G2438), .Z(n561) );
  XNOR2_X1 U633 ( .A(n562), .B(n561), .ZN(n563) );
  XOR2_X1 U634 ( .A(n564), .B(n563), .Z(n565) );
  AND2_X1 U635 ( .A1(G14), .A2(n565), .ZN(G401) );
  XNOR2_X1 U636 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  AND2_X1 U637 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U638 ( .A(G132), .ZN(G219) );
  INV_X1 U639 ( .A(G82), .ZN(G220) );
  INV_X1 U640 ( .A(G120), .ZN(G236) );
  INV_X1 U641 ( .A(G69), .ZN(G235) );
  INV_X1 U642 ( .A(G57), .ZN(G237) );
  NAND2_X1 U643 ( .A1(G138), .A2(n903), .ZN(n567) );
  NAND2_X1 U644 ( .A1(G102), .A2(n904), .ZN(n566) );
  NAND2_X1 U645 ( .A1(n567), .A2(n566), .ZN(n576) );
  AND2_X1 U646 ( .A1(n568), .A2(G126), .ZN(n569) );
  NAND2_X1 U647 ( .A1(n569), .A2(G2105), .ZN(n570) );
  XNOR2_X1 U648 ( .A(n570), .B(KEYINPUT92), .ZN(n572) );
  NAND2_X1 U649 ( .A1(G114), .A2(n898), .ZN(n571) );
  NAND2_X1 U650 ( .A1(n572), .A2(n571), .ZN(n574) );
  INV_X1 U651 ( .A(KEYINPUT93), .ZN(n573) );
  XNOR2_X1 U652 ( .A(n574), .B(n573), .ZN(n575) );
  NOR2_X1 U653 ( .A1(n576), .A2(n575), .ZN(G164) );
  NAND2_X1 U654 ( .A1(G51), .A2(n667), .ZN(n578) );
  NAND2_X1 U655 ( .A1(G63), .A2(n669), .ZN(n577) );
  NAND2_X1 U656 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U657 ( .A(KEYINPUT6), .B(n579), .ZN(n587) );
  NAND2_X1 U658 ( .A1(G89), .A2(n673), .ZN(n580) );
  XNOR2_X1 U659 ( .A(n580), .B(KEYINPUT4), .ZN(n581) );
  XNOR2_X1 U660 ( .A(n581), .B(KEYINPUT78), .ZN(n583) );
  NAND2_X1 U661 ( .A1(G76), .A2(n674), .ZN(n582) );
  NAND2_X1 U662 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U663 ( .A(KEYINPUT79), .B(n584), .ZN(n585) );
  XNOR2_X1 U664 ( .A(KEYINPUT5), .B(n585), .ZN(n586) );
  NOR2_X1 U665 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U666 ( .A(KEYINPUT7), .B(n588), .Z(G168) );
  XOR2_X1 U667 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U668 ( .A(KEYINPUT70), .B(KEYINPUT11), .Z(n591) );
  NAND2_X1 U669 ( .A1(G7), .A2(G661), .ZN(n589) );
  XOR2_X1 U670 ( .A(n589), .B(KEYINPUT10), .Z(n934) );
  NAND2_X1 U671 ( .A1(G567), .A2(n934), .ZN(n590) );
  XNOR2_X1 U672 ( .A(n591), .B(n590), .ZN(G234) );
  NAND2_X1 U673 ( .A1(n674), .A2(G68), .ZN(n593) );
  NAND2_X1 U674 ( .A1(n673), .A2(G81), .ZN(n594) );
  XNOR2_X1 U675 ( .A(KEYINPUT12), .B(n594), .ZN(n595) );
  NAND2_X1 U676 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U677 ( .A(n597), .B(KEYINPUT13), .ZN(n599) );
  NAND2_X1 U678 ( .A1(G43), .A2(n667), .ZN(n598) );
  NAND2_X1 U679 ( .A1(n599), .A2(n598), .ZN(n602) );
  NAND2_X1 U680 ( .A1(n669), .A2(G56), .ZN(n600) );
  XOR2_X1 U681 ( .A(KEYINPUT14), .B(n600), .Z(n601) );
  NAND2_X1 U682 ( .A1(G860), .A2(n989), .ZN(G153) );
  XNOR2_X1 U683 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  NAND2_X1 U684 ( .A1(G868), .A2(G301), .ZN(n604) );
  XNOR2_X1 U685 ( .A(n604), .B(KEYINPUT74), .ZN(n616) );
  NAND2_X1 U686 ( .A1(n669), .A2(G66), .ZN(n611) );
  NAND2_X1 U687 ( .A1(G92), .A2(n673), .ZN(n606) );
  NAND2_X1 U688 ( .A1(G79), .A2(n674), .ZN(n605) );
  NAND2_X1 U689 ( .A1(n606), .A2(n605), .ZN(n609) );
  NAND2_X1 U690 ( .A1(G54), .A2(n667), .ZN(n607) );
  XNOR2_X1 U691 ( .A(KEYINPUT75), .B(n607), .ZN(n608) );
  NOR2_X1 U692 ( .A1(n609), .A2(n608), .ZN(n610) );
  NAND2_X1 U693 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U694 ( .A(n612), .B(KEYINPUT76), .ZN(n614) );
  XNOR2_X1 U695 ( .A(KEYINPUT15), .B(KEYINPUT77), .ZN(n613) );
  INV_X1 U696 ( .A(G868), .ZN(n688) );
  NAND2_X1 U697 ( .A1(n717), .A2(n688), .ZN(n615) );
  NAND2_X1 U698 ( .A1(n616), .A2(n615), .ZN(G284) );
  NAND2_X1 U699 ( .A1(G91), .A2(n673), .ZN(n617) );
  XOR2_X1 U700 ( .A(KEYINPUT68), .B(n617), .Z(n622) );
  NAND2_X1 U701 ( .A1(G53), .A2(n667), .ZN(n619) );
  NAND2_X1 U702 ( .A1(G65), .A2(n669), .ZN(n618) );
  NAND2_X1 U703 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U704 ( .A(KEYINPUT69), .B(n620), .Z(n621) );
  NOR2_X1 U705 ( .A1(n622), .A2(n621), .ZN(n624) );
  NAND2_X1 U706 ( .A1(n674), .A2(G78), .ZN(n623) );
  NAND2_X1 U707 ( .A1(n624), .A2(n623), .ZN(G299) );
  XOR2_X1 U708 ( .A(KEYINPUT80), .B(G868), .Z(n625) );
  NOR2_X1 U709 ( .A1(G286), .A2(n625), .ZN(n627) );
  NOR2_X1 U710 ( .A1(G868), .A2(G299), .ZN(n626) );
  NOR2_X1 U711 ( .A1(n627), .A2(n626), .ZN(G297) );
  INV_X1 U712 ( .A(G860), .ZN(n628) );
  NAND2_X1 U713 ( .A1(n628), .A2(G559), .ZN(n629) );
  NAND2_X1 U714 ( .A1(n629), .A2(n984), .ZN(n630) );
  XNOR2_X1 U715 ( .A(n630), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U716 ( .A1(n717), .A2(n688), .ZN(n631) );
  XNOR2_X1 U717 ( .A(n631), .B(KEYINPUT81), .ZN(n632) );
  NOR2_X1 U718 ( .A1(G559), .A2(n632), .ZN(n634) );
  AND2_X1 U719 ( .A1(n989), .A2(n688), .ZN(n633) );
  NOR2_X1 U720 ( .A1(n634), .A2(n633), .ZN(G282) );
  NAND2_X1 U721 ( .A1(n896), .A2(G123), .ZN(n635) );
  XNOR2_X1 U722 ( .A(n635), .B(KEYINPUT18), .ZN(n637) );
  NAND2_X1 U723 ( .A1(G111), .A2(n898), .ZN(n636) );
  NAND2_X1 U724 ( .A1(n637), .A2(n636), .ZN(n641) );
  NAND2_X1 U725 ( .A1(G135), .A2(n903), .ZN(n639) );
  NAND2_X1 U726 ( .A1(G99), .A2(n904), .ZN(n638) );
  NAND2_X1 U727 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U728 ( .A1(n641), .A2(n640), .ZN(n936) );
  XNOR2_X1 U729 ( .A(n936), .B(G2096), .ZN(n642) );
  INV_X1 U730 ( .A(G2100), .ZN(n854) );
  NAND2_X1 U731 ( .A1(n642), .A2(n854), .ZN(G156) );
  NAND2_X1 U732 ( .A1(G55), .A2(n667), .ZN(n644) );
  NAND2_X1 U733 ( .A1(G67), .A2(n669), .ZN(n643) );
  NAND2_X1 U734 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U735 ( .A1(G93), .A2(n673), .ZN(n646) );
  NAND2_X1 U736 ( .A1(G80), .A2(n674), .ZN(n645) );
  NAND2_X1 U737 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U738 ( .A1(n648), .A2(n647), .ZN(n687) );
  NAND2_X1 U739 ( .A1(n984), .A2(G559), .ZN(n649) );
  XNOR2_X1 U740 ( .A(n649), .B(KEYINPUT82), .ZN(n685) );
  XOR2_X1 U741 ( .A(n685), .B(n989), .Z(n650) );
  NOR2_X1 U742 ( .A1(G860), .A2(n650), .ZN(n651) );
  XNOR2_X1 U743 ( .A(n687), .B(n651), .ZN(G145) );
  NAND2_X1 U744 ( .A1(G49), .A2(n667), .ZN(n653) );
  NAND2_X1 U745 ( .A1(G74), .A2(G651), .ZN(n652) );
  NAND2_X1 U746 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U747 ( .A1(n669), .A2(n654), .ZN(n655) );
  XOR2_X1 U748 ( .A(KEYINPUT83), .B(n655), .Z(n658) );
  NAND2_X1 U749 ( .A1(n656), .A2(G87), .ZN(n657) );
  NAND2_X1 U750 ( .A1(n658), .A2(n657), .ZN(G288) );
  NAND2_X1 U751 ( .A1(n669), .A2(G61), .ZN(n665) );
  NAND2_X1 U752 ( .A1(G86), .A2(n673), .ZN(n660) );
  NAND2_X1 U753 ( .A1(G48), .A2(n667), .ZN(n659) );
  NAND2_X1 U754 ( .A1(n660), .A2(n659), .ZN(n663) );
  NAND2_X1 U755 ( .A1(n674), .A2(G73), .ZN(n661) );
  XOR2_X1 U756 ( .A(KEYINPUT2), .B(n661), .Z(n662) );
  NOR2_X1 U757 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U758 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U759 ( .A(n666), .B(KEYINPUT84), .ZN(G305) );
  NAND2_X1 U760 ( .A1(n667), .A2(G50), .ZN(n668) );
  XOR2_X1 U761 ( .A(KEYINPUT85), .B(n668), .Z(n671) );
  NAND2_X1 U762 ( .A1(G62), .A2(n669), .ZN(n670) );
  NAND2_X1 U763 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U764 ( .A(KEYINPUT86), .B(n672), .ZN(n678) );
  NAND2_X1 U765 ( .A1(G88), .A2(n673), .ZN(n676) );
  NAND2_X1 U766 ( .A1(G75), .A2(n674), .ZN(n675) );
  NAND2_X1 U767 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U768 ( .A1(n678), .A2(n677), .ZN(G166) );
  INV_X1 U769 ( .A(G166), .ZN(G303) );
  XOR2_X1 U770 ( .A(G299), .B(n989), .Z(n679) );
  XNOR2_X1 U771 ( .A(n679), .B(G288), .ZN(n682) );
  XOR2_X1 U772 ( .A(KEYINPUT19), .B(n687), .Z(n680) );
  XNOR2_X1 U773 ( .A(G290), .B(n680), .ZN(n681) );
  XOR2_X1 U774 ( .A(n682), .B(n681), .Z(n684) );
  XOR2_X1 U775 ( .A(G305), .B(G303), .Z(n683) );
  XNOR2_X1 U776 ( .A(n684), .B(n683), .ZN(n922) );
  XNOR2_X1 U777 ( .A(n685), .B(n922), .ZN(n686) );
  NAND2_X1 U778 ( .A1(n686), .A2(G868), .ZN(n690) );
  NAND2_X1 U779 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U780 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U781 ( .A(KEYINPUT87), .B(n691), .ZN(G295) );
  NAND2_X1 U782 ( .A1(G2084), .A2(G2078), .ZN(n693) );
  XOR2_X1 U783 ( .A(KEYINPUT88), .B(KEYINPUT20), .Z(n692) );
  XNOR2_X1 U784 ( .A(n693), .B(n692), .ZN(n694) );
  NAND2_X1 U785 ( .A1(G2090), .A2(n694), .ZN(n695) );
  XNOR2_X1 U786 ( .A(KEYINPUT21), .B(n695), .ZN(n696) );
  NAND2_X1 U787 ( .A1(n696), .A2(G2072), .ZN(G158) );
  NOR2_X1 U788 ( .A1(G235), .A2(G236), .ZN(n697) );
  XNOR2_X1 U789 ( .A(n697), .B(KEYINPUT89), .ZN(n698) );
  NOR2_X1 U790 ( .A1(G237), .A2(n698), .ZN(n699) );
  XNOR2_X1 U791 ( .A(KEYINPUT90), .B(n699), .ZN(n700) );
  NAND2_X1 U792 ( .A1(n700), .A2(G108), .ZN(n852) );
  NAND2_X1 U793 ( .A1(G567), .A2(n852), .ZN(n701) );
  XNOR2_X1 U794 ( .A(n701), .B(KEYINPUT91), .ZN(n706) );
  NOR2_X1 U795 ( .A1(G220), .A2(G219), .ZN(n702) );
  XNOR2_X1 U796 ( .A(KEYINPUT22), .B(n702), .ZN(n703) );
  NAND2_X1 U797 ( .A1(n703), .A2(G96), .ZN(n704) );
  OR2_X1 U798 ( .A1(G218), .A2(n704), .ZN(n853) );
  AND2_X1 U799 ( .A1(G2106), .A2(n853), .ZN(n705) );
  NOR2_X1 U800 ( .A1(n706), .A2(n705), .ZN(G319) );
  INV_X1 U801 ( .A(G319), .ZN(n708) );
  NAND2_X1 U802 ( .A1(G661), .A2(G483), .ZN(n707) );
  NOR2_X1 U803 ( .A1(n708), .A2(n707), .ZN(n851) );
  NAND2_X1 U804 ( .A1(n851), .A2(G36), .ZN(G176) );
  NOR2_X1 U805 ( .A1(G164), .A2(G1384), .ZN(n810) );
  NOR2_X1 U806 ( .A1(G1981), .A2(G305), .ZN(n710) );
  XOR2_X1 U807 ( .A(n710), .B(KEYINPUT24), .Z(n711) );
  NOR2_X1 U808 ( .A1(n791), .A2(n711), .ZN(n797) );
  NAND2_X1 U809 ( .A1(G1348), .A2(n750), .ZN(n713) );
  NAND2_X1 U810 ( .A1(G2067), .A2(n736), .ZN(n712) );
  NAND2_X1 U811 ( .A1(n713), .A2(n712), .ZN(n716) );
  NOR2_X1 U812 ( .A1(n717), .A2(n716), .ZN(n723) );
  NAND2_X1 U813 ( .A1(G1996), .A2(n736), .ZN(n714) );
  XNOR2_X1 U814 ( .A(n714), .B(KEYINPUT26), .ZN(n715) );
  NAND2_X1 U815 ( .A1(n715), .A2(n989), .ZN(n721) );
  NAND2_X1 U816 ( .A1(n717), .A2(n716), .ZN(n719) );
  NAND2_X1 U817 ( .A1(G1341), .A2(n750), .ZN(n718) );
  NAND2_X1 U818 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U819 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U820 ( .A1(n723), .A2(n722), .ZN(n728) );
  NAND2_X1 U821 ( .A1(n736), .A2(G2072), .ZN(n724) );
  XNOR2_X1 U822 ( .A(n724), .B(KEYINPUT27), .ZN(n726) );
  INV_X1 U823 ( .A(G1956), .ZN(n991) );
  NOR2_X1 U824 ( .A1(n991), .A2(n736), .ZN(n725) );
  INV_X1 U825 ( .A(G299), .ZN(n990) );
  NAND2_X1 U826 ( .A1(n729), .A2(n990), .ZN(n727) );
  NAND2_X1 U827 ( .A1(n728), .A2(n727), .ZN(n733) );
  NOR2_X1 U828 ( .A1(n729), .A2(n990), .ZN(n731) );
  NAND2_X1 U829 ( .A1(n733), .A2(n732), .ZN(n735) );
  INV_X1 U830 ( .A(G1961), .ZN(n867) );
  NAND2_X1 U831 ( .A1(n750), .A2(n867), .ZN(n738) );
  XNOR2_X1 U832 ( .A(G2078), .B(KEYINPUT25), .ZN(n969) );
  NAND2_X1 U833 ( .A1(n736), .A2(n969), .ZN(n737) );
  NAND2_X1 U834 ( .A1(n738), .A2(n737), .ZN(n746) );
  NAND2_X1 U835 ( .A1(G171), .A2(n746), .ZN(n739) );
  XOR2_X1 U836 ( .A(KEYINPUT99), .B(n739), .Z(n740) );
  NAND2_X1 U837 ( .A1(n741), .A2(n740), .ZN(n759) );
  NOR2_X1 U838 ( .A1(G1966), .A2(n791), .ZN(n762) );
  NOR2_X1 U839 ( .A1(G2084), .A2(n750), .ZN(n761) );
  OR2_X1 U840 ( .A1(n762), .A2(n743), .ZN(n744) );
  XNOR2_X1 U841 ( .A(n744), .B(KEYINPUT30), .ZN(n745) );
  XNOR2_X1 U842 ( .A(KEYINPUT100), .B(n748), .ZN(n760) );
  NAND2_X1 U843 ( .A1(n759), .A2(n760), .ZN(n749) );
  NAND2_X1 U844 ( .A1(n749), .A2(G286), .ZN(n756) );
  NOR2_X1 U845 ( .A1(G1971), .A2(n791), .ZN(n752) );
  NOR2_X1 U846 ( .A1(G2090), .A2(n750), .ZN(n751) );
  NOR2_X1 U847 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U848 ( .A1(n753), .A2(G303), .ZN(n754) );
  OR2_X1 U849 ( .A1(n742), .A2(n754), .ZN(n755) );
  NAND2_X1 U850 ( .A1(n756), .A2(n755), .ZN(n758) );
  INV_X1 U851 ( .A(KEYINPUT32), .ZN(n757) );
  AND2_X1 U852 ( .A1(n760), .A2(n759), .ZN(n765) );
  AND2_X1 U853 ( .A1(G8), .A2(n761), .ZN(n763) );
  OR2_X1 U854 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U855 ( .A1(G1976), .A2(G288), .ZN(n987) );
  INV_X1 U856 ( .A(n987), .ZN(n766) );
  OR2_X1 U857 ( .A1(n766), .A2(n791), .ZN(n772) );
  INV_X1 U858 ( .A(n772), .ZN(n767) );
  AND2_X1 U859 ( .A1(n787), .A2(n767), .ZN(n768) );
  NAND2_X1 U860 ( .A1(n786), .A2(n768), .ZN(n774) );
  NOR2_X1 U861 ( .A1(G288), .A2(G1976), .ZN(n769) );
  XOR2_X1 U862 ( .A(n769), .B(KEYINPUT101), .Z(n994) );
  NOR2_X1 U863 ( .A1(G1971), .A2(G303), .ZN(n770) );
  NOR2_X1 U864 ( .A1(n994), .A2(n770), .ZN(n771) );
  OR2_X1 U865 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U866 ( .A1(n774), .A2(n773), .ZN(n776) );
  XNOR2_X1 U867 ( .A(n776), .B(n775), .ZN(n778) );
  NOR2_X1 U868 ( .A1(n791), .A2(KEYINPUT102), .ZN(n777) );
  INV_X1 U869 ( .A(KEYINPUT33), .ZN(n779) );
  NAND2_X1 U870 ( .A1(n524), .A2(n779), .ZN(n785) );
  INV_X1 U871 ( .A(n994), .ZN(n780) );
  OR2_X1 U872 ( .A1(KEYINPUT102), .A2(n780), .ZN(n783) );
  NAND2_X1 U873 ( .A1(n994), .A2(KEYINPUT33), .ZN(n781) );
  NAND2_X1 U874 ( .A1(n781), .A2(KEYINPUT102), .ZN(n782) );
  NAND2_X1 U875 ( .A1(n783), .A2(n782), .ZN(n784) );
  XOR2_X1 U876 ( .A(G1981), .B(G305), .Z(n1005) );
  NAND2_X1 U877 ( .A1(n785), .A2(n526), .ZN(n794) );
  NAND2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n790) );
  NOR2_X1 U879 ( .A1(G2090), .A2(G303), .ZN(n788) );
  NAND2_X1 U880 ( .A1(G8), .A2(n788), .ZN(n789) );
  NAND2_X1 U881 ( .A1(n790), .A2(n789), .ZN(n792) );
  NAND2_X1 U882 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U883 ( .A1(n794), .A2(n793), .ZN(n795) );
  XOR2_X1 U884 ( .A(KEYINPUT103), .B(n795), .Z(n796) );
  NOR2_X1 U885 ( .A1(n797), .A2(n796), .ZN(n830) );
  XNOR2_X1 U886 ( .A(G2067), .B(KEYINPUT37), .ZN(n842) );
  XNOR2_X1 U887 ( .A(KEYINPUT94), .B(KEYINPUT34), .ZN(n801) );
  NAND2_X1 U888 ( .A1(G140), .A2(n903), .ZN(n799) );
  NAND2_X1 U889 ( .A1(G104), .A2(n904), .ZN(n798) );
  NAND2_X1 U890 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U891 ( .A(n801), .B(n800), .ZN(n807) );
  XNOR2_X1 U892 ( .A(KEYINPUT35), .B(KEYINPUT95), .ZN(n805) );
  NAND2_X1 U893 ( .A1(G128), .A2(n896), .ZN(n803) );
  NAND2_X1 U894 ( .A1(G116), .A2(n898), .ZN(n802) );
  NAND2_X1 U895 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U896 ( .A(n805), .B(n804), .ZN(n806) );
  NOR2_X1 U897 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U898 ( .A(n808), .B(KEYINPUT36), .ZN(n919) );
  NOR2_X1 U899 ( .A1(n842), .A2(n919), .ZN(n956) );
  NAND2_X1 U900 ( .A1(G160), .A2(G40), .ZN(n809) );
  NOR2_X1 U901 ( .A1(n810), .A2(n809), .ZN(n844) );
  NAND2_X1 U902 ( .A1(n956), .A2(n844), .ZN(n811) );
  XNOR2_X1 U903 ( .A(n811), .B(KEYINPUT96), .ZN(n840) );
  NAND2_X1 U904 ( .A1(G119), .A2(n896), .ZN(n813) );
  NAND2_X1 U905 ( .A1(G131), .A2(n903), .ZN(n812) );
  NAND2_X1 U906 ( .A1(n813), .A2(n812), .ZN(n817) );
  NAND2_X1 U907 ( .A1(G107), .A2(n898), .ZN(n815) );
  NAND2_X1 U908 ( .A1(G95), .A2(n904), .ZN(n814) );
  NAND2_X1 U909 ( .A1(n815), .A2(n814), .ZN(n816) );
  OR2_X1 U910 ( .A1(n817), .A2(n816), .ZN(n914) );
  NAND2_X1 U911 ( .A1(G1991), .A2(n914), .ZN(n827) );
  NAND2_X1 U912 ( .A1(G129), .A2(n896), .ZN(n819) );
  NAND2_X1 U913 ( .A1(G141), .A2(n903), .ZN(n818) );
  NAND2_X1 U914 ( .A1(n819), .A2(n818), .ZN(n823) );
  NAND2_X1 U915 ( .A1(G105), .A2(n904), .ZN(n820) );
  XNOR2_X1 U916 ( .A(n820), .B(KEYINPUT97), .ZN(n821) );
  XNOR2_X1 U917 ( .A(n821), .B(KEYINPUT38), .ZN(n822) );
  NOR2_X1 U918 ( .A1(n823), .A2(n822), .ZN(n825) );
  NAND2_X1 U919 ( .A1(n898), .A2(G117), .ZN(n824) );
  NAND2_X1 U920 ( .A1(n825), .A2(n824), .ZN(n893) );
  NAND2_X1 U921 ( .A1(G1996), .A2(n893), .ZN(n826) );
  NAND2_X1 U922 ( .A1(n827), .A2(n826), .ZN(n937) );
  NAND2_X1 U923 ( .A1(n937), .A2(n844), .ZN(n828) );
  XNOR2_X1 U924 ( .A(KEYINPUT98), .B(n828), .ZN(n833) );
  NAND2_X1 U925 ( .A1(n840), .A2(n833), .ZN(n829) );
  NOR2_X1 U926 ( .A1(n830), .A2(n829), .ZN(n832) );
  XNOR2_X1 U927 ( .A(G1986), .B(G290), .ZN(n986) );
  NAND2_X1 U928 ( .A1(n986), .A2(n844), .ZN(n831) );
  NAND2_X1 U929 ( .A1(n832), .A2(n831), .ZN(n847) );
  NOR2_X1 U930 ( .A1(G1996), .A2(n893), .ZN(n947) );
  INV_X1 U931 ( .A(n833), .ZN(n837) );
  NOR2_X1 U932 ( .A1(G1991), .A2(n914), .ZN(n834) );
  XNOR2_X1 U933 ( .A(KEYINPUT104), .B(n834), .ZN(n938) );
  NOR2_X1 U934 ( .A1(G1986), .A2(G290), .ZN(n835) );
  NOR2_X1 U935 ( .A1(n938), .A2(n835), .ZN(n836) );
  NOR2_X1 U936 ( .A1(n837), .A2(n836), .ZN(n838) );
  NOR2_X1 U937 ( .A1(n947), .A2(n838), .ZN(n839) );
  XNOR2_X1 U938 ( .A(n839), .B(KEYINPUT39), .ZN(n841) );
  NAND2_X1 U939 ( .A1(n841), .A2(n840), .ZN(n843) );
  NAND2_X1 U940 ( .A1(n842), .A2(n919), .ZN(n953) );
  NAND2_X1 U941 ( .A1(n843), .A2(n953), .ZN(n845) );
  NAND2_X1 U942 ( .A1(n845), .A2(n844), .ZN(n846) );
  NAND2_X1 U943 ( .A1(n847), .A2(n846), .ZN(n848) );
  XNOR2_X1 U944 ( .A(KEYINPUT40), .B(n848), .ZN(G329) );
  NAND2_X1 U945 ( .A1(G2106), .A2(n934), .ZN(G217) );
  AND2_X1 U946 ( .A1(G15), .A2(G2), .ZN(n849) );
  NAND2_X1 U947 ( .A1(G661), .A2(n849), .ZN(G259) );
  NAND2_X1 U948 ( .A1(G3), .A2(G1), .ZN(n850) );
  NAND2_X1 U949 ( .A1(n851), .A2(n850), .ZN(G188) );
  INV_X1 U951 ( .A(G108), .ZN(G238) );
  INV_X1 U952 ( .A(G96), .ZN(G221) );
  NOR2_X1 U953 ( .A1(n853), .A2(n852), .ZN(G325) );
  INV_X1 U954 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U955 ( .A(n854), .B(KEYINPUT42), .ZN(n856) );
  XNOR2_X1 U956 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n855) );
  XNOR2_X1 U957 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U958 ( .A(KEYINPUT43), .B(G2072), .Z(n858) );
  XNOR2_X1 U959 ( .A(G2067), .B(G2090), .ZN(n857) );
  XNOR2_X1 U960 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U961 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U962 ( .A(G2678), .B(G2096), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n862), .B(n861), .ZN(n864) );
  XOR2_X1 U964 ( .A(G2084), .B(G2078), .Z(n863) );
  XNOR2_X1 U965 ( .A(n864), .B(n863), .ZN(G227) );
  XNOR2_X1 U966 ( .A(n991), .B(G1966), .ZN(n866) );
  XNOR2_X1 U967 ( .A(G1991), .B(G1981), .ZN(n865) );
  XNOR2_X1 U968 ( .A(n866), .B(n865), .ZN(n871) );
  XOR2_X1 U969 ( .A(G1976), .B(G1971), .Z(n869) );
  XOR2_X1 U970 ( .A(G1986), .B(n867), .Z(n868) );
  XNOR2_X1 U971 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U972 ( .A(n871), .B(n870), .Z(n873) );
  XNOR2_X1 U973 ( .A(KEYINPUT107), .B(KEYINPUT41), .ZN(n872) );
  XNOR2_X1 U974 ( .A(n873), .B(n872), .ZN(n875) );
  XOR2_X1 U975 ( .A(G1996), .B(G2474), .Z(n874) );
  XNOR2_X1 U976 ( .A(n875), .B(n874), .ZN(G229) );
  NAND2_X1 U977 ( .A1(G112), .A2(n898), .ZN(n877) );
  NAND2_X1 U978 ( .A1(G100), .A2(n904), .ZN(n876) );
  NAND2_X1 U979 ( .A1(n877), .A2(n876), .ZN(n878) );
  XNOR2_X1 U980 ( .A(KEYINPUT108), .B(n878), .ZN(n883) );
  NAND2_X1 U981 ( .A1(n896), .A2(G124), .ZN(n879) );
  XNOR2_X1 U982 ( .A(n879), .B(KEYINPUT44), .ZN(n881) );
  NAND2_X1 U983 ( .A1(G136), .A2(n903), .ZN(n880) );
  NAND2_X1 U984 ( .A1(n881), .A2(n880), .ZN(n882) );
  NOR2_X1 U985 ( .A1(n883), .A2(n882), .ZN(G162) );
  NAND2_X1 U986 ( .A1(G139), .A2(n903), .ZN(n885) );
  NAND2_X1 U987 ( .A1(G103), .A2(n904), .ZN(n884) );
  NAND2_X1 U988 ( .A1(n885), .A2(n884), .ZN(n891) );
  NAND2_X1 U989 ( .A1(n896), .A2(G127), .ZN(n886) );
  XOR2_X1 U990 ( .A(KEYINPUT113), .B(n886), .Z(n888) );
  NAND2_X1 U991 ( .A1(n898), .A2(G115), .ZN(n887) );
  NAND2_X1 U992 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U993 ( .A(KEYINPUT47), .B(n889), .Z(n890) );
  NOR2_X1 U994 ( .A1(n891), .A2(n890), .ZN(n941) );
  XNOR2_X1 U995 ( .A(G164), .B(n941), .ZN(n918) );
  XOR2_X1 U996 ( .A(G160), .B(n936), .Z(n892) );
  XNOR2_X1 U997 ( .A(n893), .B(n892), .ZN(n913) );
  XOR2_X1 U998 ( .A(KEYINPUT114), .B(KEYINPUT112), .Z(n895) );
  XNOR2_X1 U999 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n894) );
  XNOR2_X1 U1000 ( .A(n895), .B(n894), .ZN(n911) );
  NAND2_X1 U1001 ( .A1(n896), .A2(G130), .ZN(n897) );
  XNOR2_X1 U1002 ( .A(KEYINPUT109), .B(n897), .ZN(n901) );
  NAND2_X1 U1003 ( .A1(n898), .A2(G118), .ZN(n899) );
  XOR2_X1 U1004 ( .A(KEYINPUT110), .B(n899), .Z(n900) );
  NOR2_X1 U1005 ( .A1(n901), .A2(n900), .ZN(n902) );
  XNOR2_X1 U1006 ( .A(KEYINPUT111), .B(n902), .ZN(n909) );
  NAND2_X1 U1007 ( .A1(G142), .A2(n903), .ZN(n906) );
  NAND2_X1 U1008 ( .A1(G106), .A2(n904), .ZN(n905) );
  NAND2_X1 U1009 ( .A1(n906), .A2(n905), .ZN(n907) );
  XOR2_X1 U1010 ( .A(n907), .B(KEYINPUT45), .Z(n908) );
  NOR2_X1 U1011 ( .A1(n909), .A2(n908), .ZN(n910) );
  XOR2_X1 U1012 ( .A(n911), .B(n910), .Z(n912) );
  XNOR2_X1 U1013 ( .A(n913), .B(n912), .ZN(n916) );
  XNOR2_X1 U1014 ( .A(n914), .B(G162), .ZN(n915) );
  XNOR2_X1 U1015 ( .A(n916), .B(n915), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(n918), .B(n917), .ZN(n920) );
  XOR2_X1 U1017 ( .A(n920), .B(n919), .Z(n921) );
  NOR2_X1 U1018 ( .A1(G37), .A2(n921), .ZN(G395) );
  XOR2_X1 U1019 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n924) );
  XNOR2_X1 U1020 ( .A(G171), .B(n922), .ZN(n923) );
  XNOR2_X1 U1021 ( .A(n924), .B(n923), .ZN(n926) );
  XNOR2_X1 U1022 ( .A(G286), .B(n984), .ZN(n925) );
  XNOR2_X1 U1023 ( .A(n926), .B(n925), .ZN(n927) );
  NOR2_X1 U1024 ( .A1(G37), .A2(n927), .ZN(G397) );
  NOR2_X1 U1025 ( .A1(G227), .A2(G229), .ZN(n928) );
  XNOR2_X1 U1026 ( .A(n928), .B(KEYINPUT49), .ZN(n929) );
  NOR2_X1 U1027 ( .A1(G401), .A2(n929), .ZN(n930) );
  NAND2_X1 U1028 ( .A1(G319), .A2(n930), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(KEYINPUT117), .B(n931), .ZN(n933) );
  NOR2_X1 U1030 ( .A1(G395), .A2(G397), .ZN(n932) );
  NAND2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(G225) );
  INV_X1 U1032 ( .A(G225), .ZN(G308) );
  INV_X1 U1033 ( .A(n934), .ZN(G223) );
  XNOR2_X1 U1034 ( .A(KEYINPUT52), .B(KEYINPUT119), .ZN(n958) );
  XOR2_X1 U1035 ( .A(G2084), .B(G160), .Z(n935) );
  NOR2_X1 U1036 ( .A1(n936), .A2(n935), .ZN(n940) );
  NOR2_X1 U1037 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n952) );
  XOR2_X1 U1039 ( .A(G2072), .B(n941), .Z(n943) );
  XOR2_X1 U1040 ( .A(G164), .B(G2078), .Z(n942) );
  NOR2_X1 U1041 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1042 ( .A(n944), .B(KEYINPUT118), .ZN(n945) );
  XNOR2_X1 U1043 ( .A(n945), .B(KEYINPUT50), .ZN(n950) );
  XOR2_X1 U1044 ( .A(G2090), .B(G162), .Z(n946) );
  NOR2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1046 ( .A(KEYINPUT51), .B(n948), .Z(n949) );
  NAND2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n954) );
  NAND2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(n958), .B(n957), .ZN(n959) );
  NOR2_X1 U1052 ( .A1(KEYINPUT55), .A2(n959), .ZN(n960) );
  XOR2_X1 U1053 ( .A(KEYINPUT120), .B(n960), .Z(n961) );
  NAND2_X1 U1054 ( .A1(G29), .A2(n961), .ZN(n1041) );
  XNOR2_X1 U1055 ( .A(G2067), .B(G26), .ZN(n963) );
  XNOR2_X1 U1056 ( .A(G33), .B(G2072), .ZN(n962) );
  NOR2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n968) );
  XOR2_X1 U1058 ( .A(G1996), .B(G32), .Z(n964) );
  NAND2_X1 U1059 ( .A1(n964), .A2(G28), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(G25), .B(G1991), .ZN(n965) );
  NOR2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n971) );
  XOR2_X1 U1063 ( .A(G27), .B(n969), .Z(n970) );
  NOR2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(KEYINPUT53), .B(n972), .ZN(n973) );
  XNOR2_X1 U1066 ( .A(n973), .B(KEYINPUT121), .ZN(n977) );
  XOR2_X1 U1067 ( .A(G34), .B(KEYINPUT122), .Z(n975) );
  XNOR2_X1 U1068 ( .A(G2084), .B(KEYINPUT54), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(n975), .B(n974), .ZN(n976) );
  NAND2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(G35), .B(G2090), .ZN(n978) );
  NOR2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1073 ( .A(KEYINPUT55), .B(n980), .ZN(n982) );
  INV_X1 U1074 ( .A(G29), .ZN(n981) );
  NAND2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1076 ( .A1(n983), .A2(G11), .ZN(n1039) );
  INV_X1 U1077 ( .A(G16), .ZN(n1035) );
  XOR2_X1 U1078 ( .A(n1035), .B(KEYINPUT56), .Z(n1013) );
  XOR2_X1 U1079 ( .A(G1348), .B(n984), .Z(n985) );
  NOR2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n988) );
  NAND2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n1003) );
  XNOR2_X1 U1082 ( .A(G1341), .B(n989), .ZN(n1001) );
  XOR2_X1 U1083 ( .A(n991), .B(n990), .Z(n992) );
  XNOR2_X1 U1084 ( .A(n992), .B(KEYINPUT124), .ZN(n996) );
  XOR2_X1 U1085 ( .A(G171), .B(G1961), .Z(n993) );
  NOR2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n999) );
  XNOR2_X1 U1088 ( .A(G1971), .B(G166), .ZN(n997) );
  XNOR2_X1 U1089 ( .A(KEYINPUT125), .B(n997), .ZN(n998) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NOR2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1093 ( .A(KEYINPUT126), .B(n1004), .Z(n1010) );
  XNOR2_X1 U1094 ( .A(G1966), .B(G168), .ZN(n1006) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(n1007), .B(KEYINPUT57), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(KEYINPUT123), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(KEYINPUT127), .B(n1011), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1037) );
  XOR2_X1 U1101 ( .A(G5), .B(G1961), .Z(n1025) );
  XOR2_X1 U1102 ( .A(G20), .B(G1956), .Z(n1017) );
  XNOR2_X1 U1103 ( .A(G1981), .B(G6), .ZN(n1015) );
  XNOR2_X1 U1104 ( .A(G19), .B(G1341), .ZN(n1014) );
  NOR2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1020) );
  XOR2_X1 U1107 ( .A(KEYINPUT59), .B(G1348), .Z(n1018) );
  XNOR2_X1 U1108 ( .A(G4), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1109 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1110 ( .A(KEYINPUT60), .B(n1021), .Z(n1023) );
  XNOR2_X1 U1111 ( .A(G1966), .B(G21), .ZN(n1022) );
  NOR2_X1 U1112 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1113 ( .A1(n1025), .A2(n1024), .ZN(n1032) );
  XNOR2_X1 U1114 ( .A(G1971), .B(G22), .ZN(n1027) );
  XNOR2_X1 U1115 ( .A(G23), .B(G1976), .ZN(n1026) );
  NOR2_X1 U1116 ( .A1(n1027), .A2(n1026), .ZN(n1029) );
  XOR2_X1 U1117 ( .A(G1986), .B(G24), .Z(n1028) );
  NAND2_X1 U1118 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XNOR2_X1 U1119 ( .A(KEYINPUT58), .B(n1030), .ZN(n1031) );
  NOR2_X1 U1120 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1121 ( .A(KEYINPUT61), .B(n1033), .ZN(n1034) );
  NAND2_X1 U1122 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NAND2_X1 U1123 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NOR2_X1 U1124 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  NAND2_X1 U1125 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  XNOR2_X1 U1126 ( .A(KEYINPUT62), .B(n1042), .ZN(G150) );
  INV_X1 U1127 ( .A(G150), .ZN(G311) );
endmodule

