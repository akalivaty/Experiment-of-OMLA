//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 1 0 1 1 1 1 0 1 0 0 0 1 0 0 1 0 0 0 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 1 1 0 0 0 0 1 1 1 0 0 1 0 1 0 1 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  OR2_X1    g002(.A1(KEYINPUT65), .A2(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT65), .A2(G146), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(G143), .A3(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(KEYINPUT1), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n191), .A2(new_n194), .A3(new_n196), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n195), .B1(new_n191), .B2(KEYINPUT1), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n192), .A2(G143), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n189), .A2(new_n190), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n200), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n197), .B1(new_n198), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G104), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G107), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n205), .A2(G107), .ZN(new_n208));
  OAI21_X1  g022(.A(G101), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT3), .B1(new_n205), .B2(G107), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT3), .ZN(new_n211));
  INV_X1    g025(.A(G107), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n212), .A3(G104), .ZN(new_n213));
  INV_X1    g027(.A(G101), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n210), .A2(new_n213), .A3(new_n214), .A4(new_n206), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n209), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  OR2_X1    g031(.A1(new_n204), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT1), .B1(new_n202), .B2(G146), .ZN(new_n219));
  AOI22_X1  g033(.A1(new_n191), .A2(new_n194), .B1(G128), .B2(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n197), .B1(new_n220), .B2(KEYINPUT77), .ZN(new_n221));
  AND2_X1   g035(.A1(KEYINPUT65), .A2(G146), .ZN(new_n222));
  NOR2_X1   g036(.A1(KEYINPUT65), .A2(G146), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n193), .B1(new_n224), .B2(G143), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT77), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n195), .B1(new_n199), .B2(KEYINPUT1), .ZN(new_n227));
  NOR3_X1   g041(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  OAI211_X1 g042(.A(KEYINPUT78), .B(new_n217), .C1(new_n221), .C2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n226), .B1(new_n225), .B2(new_n227), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n191), .A2(new_n194), .ZN(new_n232));
  INV_X1    g046(.A(new_n227), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n232), .A2(new_n233), .A3(KEYINPUT77), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n231), .A2(new_n197), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT78), .B1(new_n235), .B2(new_n217), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n218), .B1(new_n230), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G137), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G134), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT11), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G134), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G137), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT11), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT66), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n239), .B1(new_n241), .B2(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(G131), .B1(new_n245), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n241), .A2(new_n247), .ZN(new_n250));
  INV_X1    g064(.A(new_n239), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n238), .A2(G134), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n253), .B1(new_n239), .B2(new_n241), .ZN(new_n254));
  INV_X1    g068(.A(G131), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n252), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  AND3_X1   g070(.A1(new_n249), .A2(new_n256), .A3(KEYINPUT69), .ZN(new_n257));
  AOI21_X1  g071(.A(KEYINPUT69), .B1(new_n249), .B2(new_n256), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n237), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT12), .ZN(new_n262));
  INV_X1    g076(.A(new_n256), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n255), .B1(new_n252), .B2(new_n254), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT12), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  AOI22_X1  g082(.A1(new_n261), .A2(new_n262), .B1(new_n237), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT10), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(new_n230), .B2(new_n236), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n204), .A2(KEYINPUT10), .A3(new_n217), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n210), .A2(new_n213), .A3(new_n206), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT75), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n210), .A2(new_n213), .A3(KEYINPUT75), .A4(new_n206), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(G101), .A3(new_n277), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n215), .A2(KEYINPUT4), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT76), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n278), .A2(KEYINPUT76), .A3(new_n279), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n199), .B1(new_n224), .B2(G143), .ZN(new_n285));
  NAND2_X1  g099(.A1(KEYINPUT0), .A2(G128), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(KEYINPUT0), .A2(G128), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n285), .A2(new_n289), .B1(new_n225), .B2(new_n287), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT4), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n276), .A2(new_n291), .A3(G101), .A4(new_n277), .ZN(new_n292));
  AND2_X1   g106(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n273), .B1(new_n284), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n271), .A2(new_n294), .A3(new_n259), .ZN(new_n295));
  INV_X1    g109(.A(G953), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G227), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n297), .B(KEYINPUT74), .ZN(new_n298));
  XNOR2_X1  g112(.A(G110), .B(G140), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n298), .B(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n295), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n269), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n283), .ZN(new_n303));
  AOI21_X1  g117(.A(KEYINPUT76), .B1(new_n278), .B2(new_n279), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n293), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n272), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n217), .B1(new_n221), .B2(new_n228), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT78), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT10), .B1(new_n309), .B2(new_n229), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n260), .B1(new_n306), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n300), .B1(new_n311), .B2(new_n295), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n187), .B(new_n188), .C1(new_n302), .C2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT12), .B1(new_n237), .B2(new_n260), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n309), .A2(new_n229), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n267), .B1(new_n315), .B2(new_n218), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n295), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n300), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n311), .A2(new_n295), .A3(new_n300), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(G469), .A3(new_n320), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n187), .A2(new_n188), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n313), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G221), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT9), .B(G234), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n325), .B1(new_n327), .B2(new_n188), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n324), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(G214), .B1(G237), .B2(G902), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(G110), .B(G122), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  XOR2_X1   g148(.A(G116), .B(G119), .Z(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT68), .ZN(new_n336));
  XOR2_X1   g150(.A(KEYINPUT2), .B(G113), .Z(new_n337));
  XNOR2_X1  g151(.A(new_n336), .B(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n292), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n339), .B1(new_n282), .B2(new_n283), .ZN(new_n340));
  INV_X1    g154(.A(new_n335), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n337), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT5), .ZN(new_n343));
  INV_X1    g157(.A(G119), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(new_n344), .A3(G116), .ZN(new_n345));
  OAI211_X1 g159(.A(G113), .B(new_n345), .C1(new_n335), .C2(new_n343), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n217), .A2(new_n342), .A3(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n334), .B1(new_n340), .B2(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n303), .A2(new_n304), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n333), .B(new_n347), .C1(new_n350), .C2(new_n339), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n349), .A2(new_n351), .A3(KEYINPUT6), .ZN(new_n352));
  INV_X1    g166(.A(new_n290), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(G125), .ZN(new_n354));
  OR2_X1    g168(.A1(new_n204), .A2(G125), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G224), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n357), .A2(G953), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n356), .B(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT6), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n360), .B(new_n334), .C1(new_n340), .C2(new_n348), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n352), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(KEYINPUT79), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT79), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n352), .A2(new_n364), .A3(new_n359), .A4(new_n361), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n333), .B(KEYINPUT8), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n217), .B1(new_n342), .B2(new_n346), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n366), .B1(new_n348), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT80), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT7), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n356), .B1(new_n370), .B2(new_n358), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT80), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n372), .B(new_n366), .C1(new_n348), .C2(new_n367), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n358), .A2(new_n370), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n354), .A2(new_n355), .A3(new_n374), .ZN(new_n375));
  AND4_X1   g189(.A1(new_n369), .A2(new_n371), .A3(new_n373), .A4(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(G902), .B1(new_n376), .B2(new_n351), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n363), .A2(new_n365), .A3(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(G210), .B1(G237), .B2(G902), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n363), .A2(new_n379), .A3(new_n365), .A4(new_n377), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n332), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT18), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n384), .A2(new_n255), .ZN(new_n385));
  INV_X1    g199(.A(G237), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(new_n296), .A3(G214), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n202), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n386), .A2(new_n296), .A3(G143), .A4(G214), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT82), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n385), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NOR4_X1   g207(.A1(new_n390), .A2(KEYINPUT82), .A3(new_n384), .A4(new_n255), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT81), .ZN(new_n395));
  XNOR2_X1  g209(.A(G125), .B(G140), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n224), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G140), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G125), .ZN(new_n399));
  INV_X1    g213(.A(G125), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G140), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G146), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n395), .B1(new_n397), .B2(new_n403), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n397), .A2(new_n403), .A3(new_n395), .ZN(new_n405));
  OAI22_X1  g219(.A1(new_n393), .A2(new_n394), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(G113), .B(G122), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n407), .B(new_n205), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n396), .A2(KEYINPUT16), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT71), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT16), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n410), .A2(new_n411), .A3(new_n398), .A4(G125), .ZN(new_n412));
  AND2_X1   g226(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(KEYINPUT71), .B1(new_n399), .B2(KEYINPUT16), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n413), .A2(KEYINPUT72), .A3(G146), .A4(new_n414), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n409), .A2(G146), .A3(new_n414), .A4(new_n412), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT72), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n409), .A2(new_n414), .A3(new_n412), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n192), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n415), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n390), .A2(G131), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT17), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n388), .A2(new_n255), .A3(new_n389), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n390), .A2(KEYINPUT17), .A3(G131), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n406), .B(new_n408), .C1(new_n421), .C2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT83), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AND2_X1   g244(.A1(new_n418), .A2(new_n420), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n431), .A2(new_n415), .A3(new_n426), .A4(new_n425), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n432), .A2(KEYINPUT83), .A3(new_n408), .A4(new_n406), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n422), .A2(new_n424), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n402), .B(KEYINPUT19), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n435), .B(new_n416), .C1(new_n201), .C2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n406), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n408), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n434), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n442));
  NOR2_X1   g256(.A1(G475), .A2(G902), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n430), .A2(new_n433), .B1(new_n439), .B2(new_n438), .ZN(new_n445));
  INV_X1    g259(.A(new_n443), .ZN(new_n446));
  OAI21_X1  g260(.A(KEYINPUT20), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(G475), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n432), .A2(new_n406), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n439), .ZN(new_n451));
  AOI21_X1  g265(.A(G902), .B1(new_n434), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n449), .B1(new_n452), .B2(KEYINPUT84), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT84), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n430), .A2(new_n433), .B1(new_n439), .B2(new_n450), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n454), .B1(new_n455), .B2(G902), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(G234), .A2(G237), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n458), .A2(G902), .A3(G953), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n459), .B(KEYINPUT88), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(KEYINPUT21), .B(G898), .ZN(new_n462));
  XNOR2_X1  g276(.A(KEYINPUT87), .B(G952), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n463), .A2(G953), .ZN(new_n464));
  AOI22_X1  g278(.A1(new_n461), .A2(new_n462), .B1(new_n458), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(G116), .ZN(new_n467));
  OR2_X1    g281(.A1(new_n467), .A2(G122), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n212), .B1(new_n468), .B2(KEYINPUT14), .ZN(new_n469));
  XOR2_X1   g283(.A(G116), .B(G122), .Z(new_n470));
  OR2_X1    g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n469), .A2(new_n470), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n195), .A2(G143), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT85), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n473), .B(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n202), .A2(G128), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(new_n243), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n243), .B1(new_n475), .B2(new_n476), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n471), .B(new_n472), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n475), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT13), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n476), .B(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(G134), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n470), .B(G107), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n477), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(G217), .ZN(new_n487));
  NOR3_X1   g301(.A1(new_n326), .A2(new_n487), .A3(G953), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n480), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT86), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT86), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n480), .A2(new_n486), .A3(new_n491), .A4(new_n488), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n480), .A2(new_n486), .ZN(new_n493));
  INV_X1    g307(.A(new_n488), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n490), .A2(new_n492), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n188), .ZN(new_n497));
  INV_X1    g311(.A(G478), .ZN(new_n498));
  OR2_X1    g312(.A1(new_n498), .A2(KEYINPUT15), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n497), .B(new_n499), .ZN(new_n500));
  AND4_X1   g314(.A1(new_n448), .A2(new_n457), .A3(new_n466), .A4(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n330), .A2(new_n383), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT89), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT89), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n330), .A2(new_n504), .A3(new_n383), .A4(new_n501), .ZN(new_n505));
  INV_X1    g319(.A(G472), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n290), .B1(new_n257), .B2(new_n258), .ZN(new_n507));
  INV_X1    g321(.A(new_n338), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n255), .B1(new_n239), .B2(new_n244), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(KEYINPUT67), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n204), .A2(new_n510), .A3(new_n256), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n507), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(KEYINPUT28), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n507), .A2(new_n511), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n338), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n386), .A2(new_n296), .A3(G210), .ZN(new_n517));
  XOR2_X1   g331(.A(new_n517), .B(KEYINPUT27), .Z(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT26), .B(G101), .ZN(new_n519));
  XOR2_X1   g333(.A(new_n518), .B(new_n519), .Z(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT29), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(G902), .B1(new_n516), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n507), .A2(KEYINPUT30), .A3(new_n511), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n511), .B1(new_n353), .B2(new_n265), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n525), .A2(new_n528), .A3(new_n338), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n512), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n521), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n526), .A2(new_n338), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n513), .A2(new_n532), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n531), .B(new_n522), .C1(new_n533), .C2(new_n521), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n506), .B1(new_n524), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n520), .B1(new_n513), .B2(new_n532), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n529), .A2(new_n512), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT70), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(KEYINPUT31), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(KEYINPUT31), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n537), .A2(new_n520), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n529), .A2(new_n512), .A3(new_n520), .A4(new_n541), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n539), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n536), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(G472), .A2(G902), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT32), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n533), .A2(new_n521), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n543), .A2(new_n539), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n543), .A2(new_n539), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT32), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n553), .A3(new_n546), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n535), .B1(new_n548), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n487), .B1(G234), .B2(new_n188), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT23), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n557), .B1(new_n344), .B2(G128), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n195), .A2(KEYINPUT23), .A3(G119), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n558), .B(new_n559), .C1(G119), .C2(new_n195), .ZN(new_n560));
  OR2_X1    g374(.A1(new_n560), .A2(G110), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT73), .ZN(new_n562));
  OR2_X1    g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n562), .ZN(new_n564));
  XNOR2_X1  g378(.A(G119), .B(G128), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(KEYINPUT24), .B(G110), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n563), .A2(new_n564), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n569), .A2(new_n397), .A3(new_n416), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n560), .A2(G110), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n421), .B(new_n571), .C1(new_n566), .C2(new_n567), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT22), .B(G137), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n296), .A2(G221), .A3(G234), .ZN(new_n575));
  XOR2_X1   g389(.A(new_n574), .B(new_n575), .Z(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n570), .A2(new_n572), .A3(new_n576), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT25), .B1(new_n580), .B2(new_n188), .ZN(new_n581));
  AND4_X1   g395(.A1(KEYINPUT25), .A2(new_n578), .A3(new_n188), .A4(new_n579), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n556), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n556), .A2(G902), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n555), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n503), .A2(new_n505), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(G101), .ZN(G3));
  OAI21_X1  g403(.A(G472), .B1(new_n545), .B2(G902), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n552), .A2(new_n546), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n324), .A2(new_n329), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n592), .A2(new_n593), .A3(new_n586), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n381), .A2(new_n382), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n331), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(new_n465), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n457), .A2(new_n448), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT33), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n496), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n495), .A2(KEYINPUT33), .A3(new_n489), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n498), .A2(G902), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(KEYINPUT90), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n497), .A2(new_n498), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT90), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n601), .A2(new_n607), .A3(new_n602), .A4(new_n603), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n605), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n599), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n598), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT34), .B(G104), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G6));
  XOR2_X1   g427(.A(new_n497), .B(new_n499), .Z(new_n614));
  NAND2_X1  g428(.A1(new_n457), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n444), .A2(new_n447), .A3(KEYINPUT91), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n616), .B1(KEYINPUT91), .B2(new_n444), .ZN(new_n617));
  OR2_X1    g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n598), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(new_n212), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT92), .B(KEYINPUT35), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G9));
  NOR2_X1   g436(.A1(new_n577), .A2(KEYINPUT36), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n573), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n584), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n583), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n592), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n503), .A2(new_n505), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT37), .B(G110), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT93), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n629), .B(new_n631), .ZN(G12));
  NAND4_X1  g446(.A1(new_n595), .A2(new_n331), .A3(new_n329), .A4(new_n324), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n555), .A2(new_n627), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n464), .A2(new_n458), .ZN(new_n636));
  XOR2_X1   g450(.A(new_n636), .B(KEYINPUT94), .Z(new_n637));
  OAI21_X1  g451(.A(new_n637), .B1(G900), .B2(new_n460), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n618), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n634), .A2(new_n635), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G128), .ZN(G30));
  XOR2_X1   g456(.A(KEYINPUT97), .B(KEYINPUT39), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n638), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n330), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(KEYINPUT40), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n595), .B(new_n647), .ZN(new_n648));
  AOI22_X1  g462(.A1(new_n453), .A2(new_n456), .B1(new_n447), .B2(new_n444), .ZN(new_n649));
  NOR4_X1   g463(.A1(new_n626), .A2(new_n332), .A3(new_n649), .A4(new_n500), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT40), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n330), .A2(new_n651), .A3(new_n644), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n646), .A2(new_n648), .A3(new_n650), .A4(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n548), .A2(new_n554), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n537), .A2(new_n521), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n512), .A2(new_n521), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n515), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n188), .ZN(new_n659));
  OAI21_X1  g473(.A(G472), .B1(new_n655), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n654), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT96), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n653), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(new_n202), .ZN(G45));
  AND3_X1   g479(.A1(new_n605), .A2(new_n606), .A3(new_n608), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(new_n649), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n638), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n634), .A2(new_n635), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G146), .ZN(G48));
  INV_X1    g485(.A(new_n312), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n672), .B1(new_n269), .B2(new_n301), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n188), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(G469), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n675), .A2(new_n329), .A3(new_n313), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n597), .A2(new_n587), .A3(new_n667), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT41), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G113), .ZN(G15));
  INV_X1    g494(.A(new_n618), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n597), .A2(new_n587), .A3(new_n681), .A4(new_n677), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G116), .ZN(G18));
  NAND2_X1  g497(.A1(new_n635), .A2(new_n501), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n677), .A2(new_n383), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT98), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n686), .B1(new_n684), .B2(new_n685), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G119), .ZN(G21));
  INV_X1    g505(.A(KEYINPUT100), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n692), .B1(new_n649), .B2(new_n500), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n599), .A2(KEYINPUT100), .A3(new_n614), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n383), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n586), .ZN(new_n696));
  OAI22_X1  g510(.A1(new_n550), .A2(new_n551), .B1(new_n516), .B2(new_n520), .ZN(new_n697));
  XOR2_X1   g511(.A(new_n546), .B(KEYINPUT99), .Z(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AND3_X1   g513(.A1(new_n696), .A2(new_n590), .A3(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n695), .A2(new_n700), .A3(new_n466), .A4(new_n677), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G122), .ZN(G24));
  NOR2_X1   g516(.A1(new_n596), .A2(new_n676), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n626), .A2(new_n590), .A3(new_n699), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n668), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G125), .ZN(G27));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n381), .A2(new_n331), .A3(new_n382), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n319), .A2(KEYINPUT101), .A3(G469), .A4(new_n320), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n313), .A2(new_n710), .A3(new_n323), .ZN(new_n711));
  AND2_X1   g525(.A1(new_n295), .A2(new_n300), .ZN(new_n712));
  AOI22_X1  g526(.A1(new_n317), .A2(new_n318), .B1(new_n712), .B2(new_n311), .ZN(new_n713));
  AOI21_X1  g527(.A(KEYINPUT101), .B1(new_n713), .B2(G469), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n329), .B1(new_n711), .B2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT102), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n709), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  OAI211_X1 g531(.A(KEYINPUT102), .B(new_n329), .C1(new_n711), .C2(new_n714), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n717), .A2(new_n587), .A3(new_n669), .A4(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT103), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT42), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n723), .B1(new_n719), .B2(new_n720), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n708), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n715), .A2(new_n716), .ZN(new_n726));
  INV_X1    g540(.A(new_n709), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n726), .A2(new_n718), .A3(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n728), .A2(KEYINPUT103), .A3(new_n587), .A4(new_n669), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n729), .A2(KEYINPUT104), .A3(new_n721), .A4(new_n723), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n545), .A2(KEYINPUT32), .A3(new_n547), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n553), .B1(new_n552), .B2(new_n546), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n524), .A2(new_n534), .ZN(new_n733));
  OAI22_X1  g547(.A1(new_n731), .A2(new_n732), .B1(new_n733), .B2(new_n506), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT105), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n734), .A2(new_n735), .A3(new_n696), .ZN(new_n736));
  OAI21_X1  g550(.A(KEYINPUT105), .B1(new_n555), .B2(new_n586), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n736), .A2(new_n737), .A3(KEYINPUT42), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n717), .A2(new_n669), .A3(new_n718), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n738), .A2(new_n739), .A3(KEYINPUT106), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT106), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n736), .A2(new_n737), .A3(KEYINPUT42), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n717), .A2(new_n669), .A3(new_n718), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n725), .A2(new_n730), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G131), .ZN(G33));
  NAND4_X1  g561(.A1(new_n728), .A2(KEYINPUT107), .A3(new_n587), .A4(new_n640), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT107), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n717), .A2(new_n718), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n587), .A2(new_n640), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G134), .ZN(G36));
  OAI21_X1  g568(.A(G469), .B1(new_n713), .B2(KEYINPUT45), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n713), .A2(KEYINPUT45), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT108), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n713), .A2(KEYINPUT108), .A3(KEYINPUT45), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n755), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n322), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(KEYINPUT46), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT46), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n763), .B1(new_n760), .B2(new_n322), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n762), .A2(new_n313), .A3(new_n764), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n765), .A2(new_n329), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n592), .A2(new_n626), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n649), .B(new_n609), .C1(KEYINPUT109), .C2(KEYINPUT43), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n599), .A2(new_n666), .ZN(new_n769));
  XOR2_X1   g583(.A(KEYINPUT109), .B(KEYINPUT43), .Z(new_n770));
  OAI21_X1  g584(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n767), .A2(KEYINPUT44), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT44), .B1(new_n767), .B2(new_n771), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n772), .A2(new_n773), .A3(new_n709), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n766), .A2(new_n644), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(KEYINPUT110), .B(G137), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n775), .B(new_n776), .ZN(G39));
  NOR4_X1   g591(.A1(new_n734), .A2(new_n668), .A3(new_n696), .A4(new_n709), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n765), .A2(KEYINPUT47), .A3(new_n329), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT47), .B1(new_n765), .B2(new_n329), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n778), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT111), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT111), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n784), .B(new_n778), .C1(new_n780), .C2(new_n781), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G140), .ZN(G42));
  XOR2_X1   g601(.A(new_n595), .B(new_n647), .Z(new_n788));
  NAND3_X1  g602(.A1(new_n788), .A2(new_n332), .A3(new_n677), .ZN(new_n789));
  INV_X1    g603(.A(new_n637), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n771), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n700), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT50), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n791), .A2(new_n677), .A3(new_n727), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT116), .ZN(new_n796));
  INV_X1    g610(.A(new_n704), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR4_X1   g612(.A1(new_n676), .A2(new_n709), .A3(new_n636), .A4(new_n586), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n663), .A2(new_n649), .A3(new_n666), .A4(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n794), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n780), .A2(new_n781), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n187), .B1(new_n673), .B2(new_n188), .ZN(new_n803));
  INV_X1    g617(.A(new_n313), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n802), .B1(new_n329), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n792), .A2(new_n709), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n801), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(KEYINPUT51), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(KEYINPUT117), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n809), .A2(KEYINPUT51), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n663), .A2(new_n667), .A3(new_n799), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n813), .B(new_n464), .C1(new_n685), .C2(new_n792), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n796), .A2(new_n737), .A3(new_n736), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n815), .A2(KEYINPUT48), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(KEYINPUT48), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n814), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n811), .A2(new_n812), .A3(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n717), .A2(new_n669), .A3(new_n797), .A4(new_n718), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n457), .A2(new_n500), .A3(new_n638), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n593), .A2(new_n617), .A3(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n635), .A2(new_n822), .A3(new_n727), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n824), .B1(new_n748), .B2(new_n752), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n610), .A2(KEYINPUT113), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT113), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n667), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n826), .B(new_n828), .C1(new_n599), .C2(new_n500), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n829), .A2(new_n597), .A3(new_n594), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n588), .A2(new_n629), .A3(new_n830), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n825), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n678), .A2(new_n682), .A3(new_n701), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n833), .B1(new_n688), .B2(new_n689), .ZN(new_n834));
  INV_X1    g648(.A(new_n715), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n583), .A2(new_n625), .A3(new_n638), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n836), .B1(new_n654), .B2(new_n660), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n695), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n641), .A2(new_n670), .A3(new_n838), .A4(new_n706), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT52), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n633), .A2(new_n555), .A3(new_n627), .ZN(new_n842));
  AOI22_X1  g656(.A1(new_n842), .A2(new_n640), .B1(new_n703), .B2(new_n705), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n843), .A2(KEYINPUT52), .A3(new_n670), .A4(new_n838), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n746), .A2(new_n832), .A3(new_n834), .A4(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n843), .ZN(new_n849));
  AOI21_X1  g663(.A(KEYINPUT53), .B1(new_n849), .B2(KEYINPUT52), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n848), .B1(new_n846), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT54), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n745), .A2(new_n730), .ZN(new_n853));
  AND4_X1   g667(.A1(new_n587), .A2(new_n717), .A3(new_n669), .A4(new_n718), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT42), .B1(new_n854), .B2(KEYINPUT103), .ZN(new_n855));
  AOI21_X1  g669(.A(KEYINPUT104), .B1(new_n855), .B2(new_n721), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n834), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT114), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n746), .A2(KEYINPUT114), .A3(new_n834), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n847), .B1(new_n849), .B2(KEYINPUT52), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n845), .A2(new_n831), .A3(new_n825), .A4(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n859), .A2(new_n860), .A3(new_n863), .ZN(new_n864));
  XOR2_X1   g678(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n865));
  NAND3_X1  g679(.A1(new_n864), .A2(new_n848), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n852), .A2(new_n866), .ZN(new_n867));
  OAI22_X1  g681(.A1(new_n819), .A2(new_n867), .B1(G952), .B2(G953), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n586), .A2(new_n332), .A3(new_n328), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(KEYINPUT112), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n806), .A2(KEYINPUT49), .ZN(new_n871));
  OR2_X1    g685(.A1(new_n806), .A2(KEYINPUT49), .ZN(new_n872));
  AND4_X1   g686(.A1(new_n769), .A2(new_n870), .A3(new_n871), .A4(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n873), .A2(new_n663), .A3(new_n788), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n868), .A2(new_n874), .ZN(G75));
  NOR2_X1   g689(.A1(new_n296), .A2(G952), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n864), .A2(new_n848), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n878), .A2(new_n188), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT56), .B1(new_n879), .B2(G210), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n352), .A2(new_n361), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(new_n359), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(KEYINPUT55), .Z(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n877), .B1(new_n880), .B2(new_n884), .ZN(new_n885));
  AOI211_X1 g699(.A(KEYINPUT56), .B(new_n883), .C1(new_n879), .C2(G210), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n885), .A2(new_n886), .ZN(G51));
  XOR2_X1   g701(.A(new_n760), .B(KEYINPUT119), .Z(new_n888));
  NOR3_X1   g702(.A1(new_n878), .A2(new_n188), .A3(new_n888), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n322), .B(KEYINPUT57), .ZN(new_n890));
  INV_X1    g704(.A(new_n865), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n862), .B1(new_n857), .B2(new_n858), .ZN(new_n892));
  AOI221_X4 g706(.A(new_n891), .B1(new_n846), .B2(new_n847), .C1(new_n892), .C2(new_n860), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n865), .B1(new_n864), .B2(new_n848), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n890), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n673), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n889), .B1(new_n896), .B2(KEYINPUT118), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT118), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n895), .A2(new_n898), .A3(new_n673), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n876), .B1(new_n897), .B2(new_n899), .ZN(G54));
  AND2_X1   g714(.A1(KEYINPUT58), .A2(G475), .ZN(new_n901));
  AOI211_X1 g715(.A(KEYINPUT120), .B(new_n441), .C1(new_n879), .C2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n878), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n903), .A2(G902), .A3(new_n901), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n877), .B1(new_n904), .B2(new_n445), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT120), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n906), .B1(new_n904), .B2(new_n445), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n902), .A2(new_n905), .A3(new_n907), .ZN(G60));
  NAND2_X1  g722(.A1(G478), .A2(G902), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(KEYINPUT59), .Z(new_n910));
  AOI21_X1  g724(.A(new_n910), .B1(new_n852), .B2(new_n866), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n601), .A2(new_n602), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  OR3_X1    g727(.A1(new_n911), .A2(KEYINPUT121), .A3(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(KEYINPUT121), .B1(new_n911), .B2(new_n913), .ZN(new_n915));
  OR2_X1    g729(.A1(new_n893), .A2(new_n894), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n912), .A2(new_n910), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n876), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n914), .A2(new_n915), .A3(new_n918), .ZN(G63));
  INV_X1    g733(.A(KEYINPUT61), .ZN(new_n920));
  NAND2_X1  g734(.A1(G217), .A2(G902), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT60), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n878), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n624), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n877), .B1(new_n923), .B2(new_n580), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n920), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OR2_X1    g741(.A1(new_n923), .A2(new_n580), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n928), .A2(KEYINPUT61), .A3(new_n877), .A4(new_n924), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n927), .A2(new_n929), .ZN(G66));
  OAI21_X1  g744(.A(G953), .B1(new_n462), .B2(new_n357), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n678), .A2(new_n701), .ZN(new_n932));
  INV_X1    g746(.A(new_n689), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n932), .B(new_n682), .C1(new_n933), .C2(new_n687), .ZN(new_n934));
  INV_X1    g748(.A(new_n831), .ZN(new_n935));
  OAI21_X1  g749(.A(KEYINPUT122), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT122), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n834), .A2(new_n937), .A3(new_n831), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n931), .B1(new_n939), .B2(G953), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n881), .B1(G898), .B2(new_n296), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(G69));
  AND2_X1   g756(.A1(new_n525), .A2(new_n528), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(new_n436), .Z(new_n944));
  AND3_X1   g758(.A1(new_n641), .A2(new_n670), .A3(new_n706), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT62), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n945), .B(new_n946), .C1(new_n663), .C2(new_n653), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n641), .A2(new_n670), .A3(new_n706), .ZN(new_n948));
  OAI21_X1  g762(.A(KEYINPUT62), .B1(new_n664), .B2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n645), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n829), .A2(new_n950), .A3(new_n587), .A4(new_n727), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n775), .A2(new_n947), .A3(new_n949), .A4(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n786), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n944), .B1(new_n954), .B2(new_n296), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n736), .A2(new_n737), .A3(new_n695), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n766), .A2(new_n956), .A3(new_n644), .ZN(new_n957));
  AND4_X1   g771(.A1(new_n753), .A2(new_n957), .A3(new_n775), .A4(new_n945), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n786), .A2(new_n746), .A3(new_n958), .ZN(new_n959));
  OR2_X1    g773(.A1(new_n959), .A2(G953), .ZN(new_n960));
  INV_X1    g774(.A(new_n944), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n961), .B1(G900), .B2(G953), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n955), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n296), .B1(G227), .B2(G900), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n963), .B(new_n964), .Z(G72));
  NAND2_X1  g779(.A1(G472), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT63), .Z(new_n967));
  NAND2_X1  g781(.A1(new_n936), .A2(new_n938), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n967), .B1(new_n954), .B2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT123), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n969), .A2(new_n970), .A3(new_n655), .ZN(new_n971));
  INV_X1    g785(.A(new_n967), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n952), .B1(new_n783), .B2(new_n785), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n972), .B1(new_n973), .B2(new_n939), .ZN(new_n974));
  INV_X1    g788(.A(new_n655), .ZN(new_n975));
  OAI21_X1  g789(.A(KEYINPUT123), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n967), .B1(new_n531), .B2(KEYINPUT126), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT126), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n978), .B1(new_n537), .B2(new_n520), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n977), .B1(new_n531), .B2(new_n979), .ZN(new_n980));
  AOI22_X1  g794(.A1(new_n971), .A2(new_n976), .B1(new_n851), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n967), .B1(new_n959), .B2(new_n968), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n657), .A2(new_n529), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT124), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(KEYINPUT125), .B1(new_n985), .B2(new_n877), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT125), .ZN(new_n987));
  AOI211_X1 g801(.A(new_n987), .B(new_n876), .C1(new_n982), .C2(new_n984), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n981), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(KEYINPUT127), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT127), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n981), .B(new_n991), .C1(new_n986), .C2(new_n988), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n990), .A2(new_n992), .ZN(G57));
endmodule


