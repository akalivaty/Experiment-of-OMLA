//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 1 0 0 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 0 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n563,
    new_n564, new_n565, new_n566, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n576, new_n578, new_n579, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n593, new_n594, new_n596, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n624, new_n627, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1171, new_n1172,
    new_n1173;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XOR2_X1   g011(.A(new_n436), .B(KEYINPUT65), .Z(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n437), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT67), .Z(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(KEYINPUT68), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n470), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT69), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n464), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n480), .B1(KEYINPUT3), .B2(new_n466), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n479), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n475), .A2(G137), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n466), .A2(G2105), .ZN(new_n486));
  AOI22_X1  g061(.A1(new_n484), .A2(new_n485), .B1(G101), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n478), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G160));
  NAND2_X1  g064(.A1(new_n484), .A2(new_n471), .ZN(new_n490));
  INV_X1    g065(.A(G136), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g067(.A(new_n492), .B(KEYINPUT71), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n483), .A2(new_n475), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n493), .B1(G124), .B2(new_n494), .ZN(new_n495));
  OAI221_X1 g070(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n475), .C2(G112), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n495), .A2(new_n496), .ZN(G162));
  INV_X1    g072(.A(KEYINPUT73), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n473), .A2(G2105), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n471), .A2(KEYINPUT68), .ZN(new_n500));
  OAI21_X1  g075(.A(G138), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n498), .B1(new_n483), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n467), .A2(KEYINPUT70), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(new_n465), .ZN(new_n504));
  INV_X1    g079(.A(G138), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n505), .B1(new_n472), .B2(new_n474), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n504), .A2(new_n506), .A3(KEYINPUT73), .A4(new_n479), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n502), .A2(KEYINPUT4), .A3(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT74), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT74), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT4), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT3), .B(G2104), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n475), .A2(new_n513), .A3(new_n514), .A4(G138), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT75), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g092(.A1(new_n506), .A2(KEYINPUT75), .A3(new_n514), .A4(new_n513), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n508), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT72), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n486), .A2(G102), .ZN(new_n522));
  OAI211_X1 g097(.A(G126), .B(new_n479), .C1(new_n481), .C2(new_n482), .ZN(new_n523));
  NAND2_X1  g098(.A1(G114), .A2(G2104), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI211_X1 g100(.A(new_n521), .B(new_n522), .C1(new_n525), .C2(new_n471), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n471), .B1(new_n523), .B2(new_n524), .ZN(new_n527));
  INV_X1    g102(.A(new_n522), .ZN(new_n528));
  OAI21_X1  g103(.A(KEYINPUT72), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n520), .A2(new_n526), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT76), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT76), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n520), .A2(new_n526), .A3(new_n532), .A4(new_n529), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(G164));
  AND3_X1   g109(.A1(KEYINPUT77), .A2(KEYINPUT6), .A3(G651), .ZN(new_n535));
  AOI21_X1  g110(.A(KEYINPUT6), .B1(KEYINPUT77), .B2(G651), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G50), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT78), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n538), .A2(KEYINPUT5), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT5), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n546), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G651), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n537), .A2(new_n545), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G88), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n541), .A2(new_n549), .A3(new_n551), .ZN(G303));
  INV_X1    g127(.A(G303), .ZN(G166));
  NAND3_X1  g128(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT79), .ZN(new_n555));
  XOR2_X1   g130(.A(new_n555), .B(KEYINPUT7), .Z(new_n556));
  NAND2_X1  g131(.A1(new_n539), .A2(G51), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n535), .A2(new_n536), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n558), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n557), .B1(new_n559), .B2(new_n545), .ZN(new_n560));
  OR2_X1    g135(.A1(new_n556), .A2(new_n560), .ZN(G286));
  INV_X1    g136(.A(G286), .ZN(G168));
  AOI22_X1  g137(.A1(new_n546), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n563), .A2(new_n548), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n564), .B1(G52), .B2(new_n539), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n550), .A2(G90), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(G301));
  INV_X1    g142(.A(G301), .ZN(G171));
  NAND2_X1  g143(.A1(new_n539), .A2(G43), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n558), .A2(new_n546), .ZN(new_n570));
  XNOR2_X1  g145(.A(KEYINPUT80), .B(G81), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n546), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n572));
  OAI221_X1 g147(.A(new_n569), .B1(new_n570), .B2(new_n571), .C1(new_n572), .C2(new_n548), .ZN(new_n573));
  INV_X1    g148(.A(G860), .ZN(new_n574));
  OR2_X1    g149(.A1(new_n573), .A2(new_n574), .ZN(G153));
  AND3_X1   g150(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G36), .ZN(G176));
  NAND2_X1  g152(.A1(G1), .A2(G3), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT8), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n576), .A2(new_n579), .ZN(G188));
  NAND2_X1  g155(.A1(G78), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G65), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n545), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(G651), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT82), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT81), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n570), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n550), .A2(KEYINPUT81), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(G91), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n539), .A2(G53), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n593), .B(KEYINPUT9), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n592), .A2(new_n594), .ZN(G299));
  OR2_X1    g170(.A1(new_n546), .A2(G74), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G651), .B1(G49), .B2(new_n539), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n550), .B(new_n586), .ZN(new_n598));
  INV_X1    g173(.A(G87), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(G288));
  NAND2_X1  g175(.A1(G73), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G61), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n545), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(G48), .A2(new_n539), .B1(new_n603), .B2(G651), .ZN(new_n604));
  INV_X1    g179(.A(G86), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n598), .B2(new_n605), .ZN(G305));
  NAND2_X1  g181(.A1(new_n550), .A2(G85), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n539), .A2(G47), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n546), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n609));
  OAI211_X1 g184(.A(new_n607), .B(new_n608), .C1(new_n609), .C2(new_n548), .ZN(G290));
  NAND2_X1  g185(.A1(G301), .A2(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n539), .A2(G54), .ZN(new_n612));
  NAND2_X1  g187(.A1(G79), .A2(G543), .ZN(new_n613));
  INV_X1    g188(.A(G66), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n545), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G651), .ZN(new_n616));
  AND3_X1   g191(.A1(new_n589), .A2(KEYINPUT10), .A3(G92), .ZN(new_n617));
  AOI21_X1  g192(.A(KEYINPUT10), .B1(new_n589), .B2(G92), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n612), .B(new_n616), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n611), .B1(new_n620), .B2(G868), .ZN(G284));
  OAI21_X1  g196(.A(new_n611), .B1(new_n620), .B2(G868), .ZN(G321));
  INV_X1    g197(.A(G868), .ZN(new_n623));
  NAND2_X1  g198(.A1(G299), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(new_n623), .B2(G168), .ZN(G297));
  OAI21_X1  g200(.A(new_n624), .B1(new_n623), .B2(G168), .ZN(G280));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n620), .B1(new_n627), .B2(G860), .ZN(G148));
  NAND2_X1  g203(.A1(new_n573), .A2(new_n623), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n619), .A2(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(new_n623), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g207(.A1(new_n514), .A2(new_n486), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT12), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT13), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(G2100), .Z(new_n636));
  NAND2_X1  g211(.A1(new_n494), .A2(G123), .ZN(new_n637));
  OAI21_X1  g212(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n638));
  INV_X1    g213(.A(KEYINPUT83), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n640), .B(new_n641), .C1(G111), .C2(new_n475), .ZN(new_n642));
  INV_X1    g217(.A(G135), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n637), .B(new_n642), .C1(new_n490), .C2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(G2096), .Z(new_n645));
  NAND2_X1  g220(.A1(new_n636), .A2(new_n645), .ZN(G156));
  XNOR2_X1  g221(.A(G2451), .B(G2454), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  XOR2_X1   g223(.A(G2443), .B(G2446), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(KEYINPUT15), .B(G2435), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2438), .ZN(new_n654));
  XOR2_X1   g229(.A(G2427), .B(G2430), .Z(new_n655));
  INV_X1    g230(.A(KEYINPUT14), .ZN(new_n656));
  AOI22_X1  g231(.A1(new_n654), .A2(new_n655), .B1(KEYINPUT84), .B2(new_n656), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(KEYINPUT84), .ZN(new_n658));
  OAI211_X1 g233(.A(new_n657), .B(new_n658), .C1(new_n654), .C2(new_n655), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n652), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(G14), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(G401));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2067), .B(G2678), .Z(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n665), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n667), .A2(new_n668), .A3(KEYINPUT17), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT18), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2072), .B(G2078), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n671), .B(new_n672), .C1(new_n670), .C2(new_n666), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n673), .B1(new_n672), .B2(new_n671), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2096), .B(G2100), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G227));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XOR2_X1   g252(.A(G1961), .B(G1966), .Z(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n677), .A2(new_n678), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT85), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n683), .B1(new_n686), .B2(KEYINPUT20), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n680), .A2(new_n682), .A3(new_n684), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n687), .B(new_n688), .C1(KEYINPUT20), .C2(new_n686), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT86), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G1991), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(G1981), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1986), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n691), .A2(new_n695), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(G229));
  MUX2_X1   g273(.A(G23), .B(G288), .S(G16), .Z(new_n699));
  NOR2_X1   g274(.A1(new_n699), .A2(KEYINPUT33), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n699), .A2(KEYINPUT33), .ZN(new_n702));
  AOI21_X1  g277(.A(G1976), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n702), .ZN(new_n704));
  INV_X1    g279(.A(G1976), .ZN(new_n705));
  NOR3_X1   g280(.A1(new_n704), .A2(new_n700), .A3(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT90), .ZN(new_n708));
  INV_X1    g283(.A(G22), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(G16), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n709), .A2(G16), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G303), .B2(G16), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n710), .B1(new_n712), .B2(new_n708), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT91), .B(G1971), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n714), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G16), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G6), .ZN(new_n719));
  INV_X1    g294(.A(G305), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(new_n718), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT32), .B(G1981), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n707), .A2(new_n717), .A3(new_n723), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n724), .A2(KEYINPUT34), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(KEYINPUT34), .ZN(new_n726));
  INV_X1    g301(.A(G25), .ZN(new_n727));
  OAI21_X1  g302(.A(KEYINPUT87), .B1(new_n727), .B2(G29), .ZN(new_n728));
  OR3_X1    g303(.A1(new_n727), .A2(KEYINPUT87), .A3(G29), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n494), .A2(G119), .ZN(new_n730));
  OAI221_X1 g305(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n475), .C2(G107), .ZN(new_n731));
  INV_X1    g306(.A(G131), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n730), .B(new_n731), .C1(new_n490), .C2(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT88), .ZN(new_n734));
  INV_X1    g309(.A(G29), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n728), .B(new_n729), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT35), .B(G1991), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT89), .Z(new_n738));
  XNOR2_X1  g313(.A(new_n736), .B(new_n738), .ZN(new_n739));
  MUX2_X1   g314(.A(G24), .B(G290), .S(G16), .Z(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(G1986), .Z(new_n741));
  NAND4_X1  g316(.A1(new_n725), .A2(new_n726), .A3(new_n739), .A4(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT92), .B(KEYINPUT36), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n726), .A2(new_n741), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n746), .A2(new_n739), .A3(new_n725), .A4(new_n743), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n718), .A2(G4), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n620), .B2(new_n718), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(G1348), .Z(new_n751));
  AND2_X1   g326(.A1(new_n735), .A2(G26), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n494), .A2(G128), .ZN(new_n753));
  OAI221_X1 g328(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n475), .C2(G116), .ZN(new_n754));
  INV_X1    g329(.A(G140), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n753), .B(new_n754), .C1(new_n490), .C2(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n752), .B1(new_n756), .B2(G29), .ZN(new_n757));
  MUX2_X1   g332(.A(new_n752), .B(new_n757), .S(KEYINPUT28), .Z(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G2067), .ZN(new_n759));
  MUX2_X1   g334(.A(G19), .B(new_n573), .S(G16), .Z(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT93), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G1341), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n751), .A2(new_n759), .A3(new_n762), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT94), .Z(new_n764));
  NOR2_X1   g339(.A1(G27), .A2(G29), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G164), .B2(G29), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G2078), .ZN(new_n767));
  NOR2_X1   g342(.A1(G29), .A2(G32), .ZN(new_n768));
  INV_X1    g343(.A(new_n490), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(G141), .ZN(new_n770));
  NAND3_X1  g345(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT26), .Z(new_n772));
  NAND2_X1  g347(.A1(new_n494), .A2(G129), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n486), .A2(G105), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n770), .A2(new_n772), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n768), .B1(new_n776), .B2(G29), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT27), .B(G1996), .Z(new_n778));
  OR2_X1    g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(G34), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n780), .A2(KEYINPUT24), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(KEYINPUT24), .ZN(new_n782));
  AOI21_X1  g357(.A(G29), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n488), .B2(G29), .ZN(new_n784));
  INV_X1    g359(.A(G2084), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OR2_X1    g361(.A1(G29), .A2(G33), .ZN(new_n787));
  INV_X1    g362(.A(G139), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n514), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n789));
  OAI22_X1  g364(.A1(new_n490), .A2(new_n788), .B1(new_n475), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT25), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT95), .Z(new_n794));
  OAI21_X1  g369(.A(new_n787), .B1(new_n794), .B2(new_n735), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n795), .A2(G2072), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n795), .A2(G2072), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n779), .B(new_n786), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT96), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n767), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(G299), .A2(G16), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n803), .A2(KEYINPUT23), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n718), .A2(G20), .ZN(new_n805));
  MUX2_X1   g380(.A(KEYINPUT23), .B(new_n804), .S(new_n805), .Z(new_n806));
  OR2_X1    g381(.A1(new_n806), .A2(G1956), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(G1956), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n735), .A2(G35), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G162), .B2(new_n735), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT29), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(G2090), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n807), .B(new_n808), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT98), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G5), .B2(G16), .ZN(new_n816));
  OR3_X1    g391(.A1(new_n815), .A2(G5), .A3(G16), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n816), .B(new_n817), .C1(G301), .C2(new_n718), .ZN(new_n818));
  INV_X1    g393(.A(G1961), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n818), .A2(new_n819), .ZN(new_n821));
  INV_X1    g396(.A(G28), .ZN(new_n822));
  AOI21_X1  g397(.A(G29), .B1(new_n822), .B2(KEYINPUT30), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(KEYINPUT30), .B2(new_n822), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n644), .B2(new_n735), .ZN(new_n825));
  NOR3_X1   g400(.A1(new_n820), .A2(new_n821), .A3(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT31), .B(G11), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n718), .A2(G21), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(G168), .B2(new_n718), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT97), .B(G1966), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n777), .A2(new_n778), .B1(new_n785), .B2(new_n784), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n826), .A2(new_n827), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n814), .A2(new_n833), .ZN(new_n834));
  AND3_X1   g409(.A1(new_n764), .A2(new_n802), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n812), .A2(new_n813), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n748), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(KEYINPUT99), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT99), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n748), .A2(new_n835), .A3(new_n839), .A4(new_n836), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n838), .A2(new_n840), .ZN(G311));
  INV_X1    g416(.A(KEYINPUT100), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n837), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n748), .A2(new_n835), .A3(KEYINPUT100), .A4(new_n836), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(G150));
  NAND2_X1  g420(.A1(new_n539), .A2(G55), .ZN(new_n846));
  INV_X1    g421(.A(G93), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n846), .B1(new_n847), .B2(new_n570), .ZN(new_n848));
  NAND2_X1  g423(.A1(G80), .A2(G543), .ZN(new_n849));
  INV_X1    g424(.A(G67), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n849), .B1(new_n545), .B2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT101), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n848), .B1(new_n852), .B2(G651), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n853), .A2(new_n574), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT37), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n620), .A2(G559), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT38), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n853), .A2(new_n573), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n853), .A2(new_n573), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT39), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n857), .B(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n855), .B1(new_n862), .B2(G860), .ZN(G145));
  INV_X1    g438(.A(new_n634), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n644), .B(KEYINPUT102), .Z(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n866), .A2(G160), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n865), .A2(new_n488), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n868), .A2(new_n870), .A3(G162), .ZN(new_n871));
  INV_X1    g446(.A(G162), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n872), .B1(new_n867), .B2(new_n869), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT105), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n871), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n874), .B1(new_n871), .B2(new_n873), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n864), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n871), .A2(new_n873), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(KEYINPUT105), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n871), .A2(new_n873), .A3(new_n874), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(new_n880), .A3(new_n634), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n475), .A2(G118), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n466), .B1(new_n883), .B2(KEYINPUT104), .ZN(new_n884));
  OAI221_X1 g459(.A(new_n884), .B1(KEYINPUT104), .B2(new_n883), .C1(G106), .C2(G2105), .ZN(new_n885));
  AOI22_X1  g460(.A1(new_n769), .A2(G142), .B1(G130), .B2(new_n494), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n733), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n756), .B(KEYINPUT103), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n527), .A2(new_n528), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n890), .A2(new_n520), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n890), .B1(new_n520), .B2(new_n891), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(new_n776), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n775), .B1(new_n892), .B2(new_n893), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n794), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n895), .B(new_n896), .C1(new_n790), .C2(new_n792), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n889), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(new_n889), .A3(new_n900), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n882), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n903), .ZN(new_n905));
  OAI211_X1 g480(.A(new_n881), .B(new_n877), .C1(new_n905), .C2(new_n901), .ZN(new_n906));
  XOR2_X1   g481(.A(KEYINPUT106), .B(G37), .Z(new_n907));
  NAND3_X1  g482(.A1(new_n904), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g484(.A(G303), .B(G290), .Z(new_n910));
  XOR2_X1   g485(.A(G288), .B(G305), .Z(new_n911));
  OR2_X1    g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n911), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n912), .A2(KEYINPUT109), .A3(new_n913), .ZN(new_n915));
  AOI21_X1  g490(.A(KEYINPUT109), .B1(new_n912), .B2(new_n913), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  MUX2_X1   g493(.A(new_n914), .B(new_n918), .S(KEYINPUT42), .Z(new_n919));
  NAND2_X1  g494(.A1(G299), .A2(KEYINPUT107), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n592), .A2(new_n921), .A3(new_n594), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n620), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(G299), .A2(KEYINPUT107), .A3(new_n619), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  XOR2_X1   g501(.A(new_n630), .B(new_n860), .Z(new_n927));
  OR2_X1    g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT108), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT41), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n930), .B1(new_n923), .B2(new_n924), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n923), .A2(new_n930), .A3(new_n924), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n929), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n929), .B1(new_n925), .B2(KEYINPUT41), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(new_n927), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n919), .A2(new_n928), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n919), .B1(new_n928), .B2(new_n938), .ZN(new_n940));
  OAI21_X1  g515(.A(G868), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(G868), .B2(new_n853), .ZN(G295));
  OAI21_X1  g517(.A(new_n941), .B1(G868), .B2(new_n853), .ZN(G331));
  NOR2_X1   g518(.A1(new_n860), .A2(G171), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n860), .A2(G171), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n945), .A2(G168), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(G168), .B1(new_n945), .B2(new_n946), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n926), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n917), .B(new_n950), .C1(new_n937), .C2(new_n949), .ZN(new_n951));
  INV_X1    g526(.A(new_n933), .ZN(new_n952));
  OAI21_X1  g527(.A(KEYINPUT108), .B1(new_n952), .B2(new_n931), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n949), .B1(new_n953), .B2(new_n935), .ZN(new_n954));
  INV_X1    g529(.A(new_n950), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n918), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(G37), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n951), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT43), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n949), .B1(new_n933), .B2(new_n932), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n918), .B1(new_n961), .B2(new_n955), .ZN(new_n962));
  AND4_X1   g537(.A1(KEYINPUT43), .A2(new_n951), .A3(new_n962), .A4(new_n907), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT44), .B1(new_n960), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n951), .A2(new_n962), .A3(new_n959), .A4(new_n907), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n964), .A2(new_n969), .ZN(G397));
  NAND2_X1  g545(.A1(G303), .A2(G8), .ZN(new_n971));
  XOR2_X1   g546(.A(new_n971), .B(KEYINPUT55), .Z(new_n972));
  NAND2_X1  g547(.A1(new_n520), .A2(new_n891), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT50), .ZN(new_n974));
  INV_X1    g549(.A(G1384), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n973), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n478), .A2(G40), .A3(new_n487), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n531), .A2(new_n975), .A3(new_n533), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n978), .B1(new_n979), .B2(KEYINPUT50), .ZN(new_n980));
  XNOR2_X1  g555(.A(KEYINPUT111), .B(G2090), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n973), .A2(KEYINPUT45), .A3(new_n975), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n977), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT45), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n984), .B1(new_n979), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n986), .A2(G1971), .ZN(new_n987));
  OAI211_X1 g562(.A(G8), .B(new_n972), .C1(new_n982), .C2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n973), .A2(new_n975), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n478), .A2(G40), .A3(new_n487), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G8), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(G288), .A2(new_n705), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT52), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NOR2_X1   g572(.A1(G305), .A2(G1981), .ZN(new_n998));
  INV_X1    g573(.A(G1981), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n550), .A2(G86), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n999), .B1(new_n604), .B2(new_n1000), .ZN(new_n1001));
  OR3_X1    g576(.A1(new_n998), .A2(KEYINPUT49), .A3(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT49), .B1(new_n998), .B2(new_n1001), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n994), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT52), .B1(G288), .B2(new_n705), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n994), .B(new_n1006), .C1(new_n705), .C2(G288), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n997), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n989), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(G288), .A2(G1976), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n1010), .B(KEYINPUT112), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1011), .A2(new_n1003), .A3(new_n1002), .ZN(new_n1012));
  INV_X1    g587(.A(new_n998), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n995), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1008), .A2(new_n988), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n531), .A2(KEYINPUT45), .A3(new_n975), .A4(new_n533), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n991), .B1(new_n990), .B2(new_n985), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1966), .ZN(new_n1019));
  AOI22_X1  g594(.A1(new_n980), .A2(new_n785), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n1020), .A2(new_n993), .A3(G286), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT63), .ZN(new_n1022));
  OAI21_X1  g597(.A(G8), .B1(new_n982), .B2(new_n987), .ZN(new_n1023));
  INV_X1    g598(.A(new_n972), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1022), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1015), .A2(new_n1021), .A3(new_n1025), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n531), .A2(new_n974), .A3(new_n975), .A4(new_n533), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n991), .B1(new_n990), .B2(KEYINPUT50), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n1027), .A2(new_n981), .A3(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(G8), .B1(new_n987), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(new_n1024), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1031), .A2(new_n1008), .A3(new_n1021), .A4(new_n988), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n1022), .ZN(new_n1033));
  AOI211_X1 g608(.A(new_n1009), .B(new_n1014), .C1(new_n1026), .C2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n980), .A2(new_n785), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n993), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(G286), .A2(G8), .ZN(new_n1038));
  XOR2_X1   g613(.A(new_n1038), .B(KEYINPUT119), .Z(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT120), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT120), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1042), .B(new_n1039), .C1(new_n1020), .C2(new_n993), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1041), .A2(KEYINPUT51), .A3(new_n1043), .ZN(new_n1044));
  OR2_X1    g619(.A1(new_n1020), .A2(new_n1039), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT51), .ZN(new_n1046));
  OAI211_X1 g621(.A(KEYINPUT120), .B(new_n1046), .C1(new_n1037), .C2(new_n1040), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1044), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT62), .ZN(new_n1049));
  AOI211_X1 g624(.A(G2078), .B(new_n984), .C1(new_n985), .C2(new_n979), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT122), .B1(new_n1050), .B2(KEYINPUT53), .ZN(new_n1051));
  OR2_X1    g626(.A1(new_n980), .A2(G1961), .ZN(new_n1052));
  INV_X1    g627(.A(G2078), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n986), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT122), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1016), .A2(new_n1053), .A3(new_n1017), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT121), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT121), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1016), .A2(new_n1017), .A3(new_n1060), .A4(new_n1053), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1059), .A2(KEYINPUT53), .A3(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1051), .A2(new_n1052), .A3(new_n1057), .A4(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(G171), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT123), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT123), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1063), .A2(new_n1066), .A3(G171), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1015), .A2(new_n1031), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT62), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1044), .A2(new_n1070), .A3(new_n1045), .A4(new_n1047), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1049), .A2(new_n1068), .A3(new_n1069), .A4(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT56), .B(G2072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n986), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1075));
  INV_X1    g650(.A(G1956), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1074), .A2(KEYINPUT116), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(KEYINPUT116), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT114), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n591), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n585), .A2(new_n590), .A3(KEYINPUT114), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1082), .A2(new_n594), .A3(new_n1083), .ZN(new_n1084));
  XOR2_X1   g659(.A(KEYINPUT113), .B(KEYINPUT57), .Z(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n594), .A2(new_n585), .A3(KEYINPUT57), .A4(new_n590), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT115), .ZN(new_n1088));
  XNOR2_X1  g663(.A(new_n1087), .B(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1074), .A2(new_n1090), .A3(new_n1077), .ZN(new_n1092));
  INV_X1    g667(.A(G2067), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n992), .A2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1094), .B1(new_n980), .B2(G1348), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1095), .A2(new_n620), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1080), .A2(new_n1091), .B1(new_n1092), .B2(new_n1096), .ZN(new_n1097));
  OAI211_X1 g672(.A(KEYINPUT60), .B(new_n1094), .C1(new_n980), .C2(G1348), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1098), .A2(KEYINPUT118), .A3(new_n619), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT60), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1095), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1098), .A2(KEYINPUT118), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1103), .A2(new_n619), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1098), .A2(KEYINPUT118), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1102), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT61), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1092), .A2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1074), .A2(new_n1077), .A3(KEYINPUT61), .A4(new_n1090), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1090), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n573), .A2(KEYINPUT117), .ZN(new_n1112));
  AOI211_X1 g687(.A(G1996), .B(new_n984), .C1(new_n985), .C2(new_n979), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT58), .B(G1341), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n992), .A2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1112), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1111), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  OAI211_X1 g693(.A(KEYINPUT59), .B(new_n1112), .C1(new_n1113), .C2(new_n1115), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1110), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1097), .B1(new_n1106), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT124), .ZN(new_n1122));
  OAI21_X1  g697(.A(G40), .B1(new_n487), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1123), .B1(new_n1122), .B2(new_n487), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n983), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(G1384), .B1(new_n520), .B2(new_n891), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1126), .A2(KEYINPUT45), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n477), .A2(KEYINPUT53), .ZN(new_n1128));
  OR4_X1    g703(.A1(G2078), .A2(new_n1125), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1051), .A2(new_n1129), .A3(new_n1052), .A4(new_n1057), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(G171), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1131), .B(KEYINPUT54), .C1(G171), .C2(new_n1063), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1121), .A2(new_n1069), .A3(new_n1132), .A4(new_n1048), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1063), .A2(new_n1066), .A3(G171), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1066), .B1(new_n1063), .B2(G171), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n1130), .A2(G171), .ZN(new_n1137));
  AOI21_X1  g712(.A(KEYINPUT54), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1034), .B(new_n1072), .C1(new_n1133), .C2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1127), .A2(new_n977), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n1140), .B(KEYINPUT110), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n756), .B(new_n1093), .ZN(new_n1142));
  INV_X1    g717(.A(G1996), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1142), .B1(new_n776), .B2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1140), .A2(G1996), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1141), .A2(new_n1144), .B1(new_n776), .B2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n733), .B(new_n737), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1141), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1140), .ZN(new_n1150));
  XNOR2_X1  g725(.A(G290), .B(G1986), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1149), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1139), .A2(new_n1152), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1140), .A2(G1986), .A3(G290), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT127), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(KEYINPUT48), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1156), .A2(new_n1149), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1142), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1141), .B1(new_n775), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1145), .B1(KEYINPUT125), .B2(KEYINPUT46), .ZN(new_n1160));
  XOR2_X1   g735(.A(KEYINPUT125), .B(KEYINPUT46), .Z(new_n1161));
  OAI211_X1 g736(.A(new_n1159), .B(new_n1160), .C1(new_n1145), .C2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1162), .B(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(new_n737), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1146), .A2(new_n734), .A3(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1166), .B1(G2067), .B2(new_n756), .ZN(new_n1167));
  AOI211_X1 g742(.A(new_n1157), .B(new_n1164), .C1(new_n1141), .C2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1153), .A2(new_n1168), .ZN(G329));
  assign    G231 = 1'b0;
  AND3_X1   g744(.A1(new_n696), .A2(new_n661), .A3(new_n697), .ZN(new_n1171));
  AND2_X1   g745(.A1(new_n908), .A2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g746(.A1(G227), .A2(new_n461), .ZN(new_n1173));
  AND3_X1   g747(.A1(new_n1172), .A2(new_n967), .A3(new_n1173), .ZN(G308));
  NAND3_X1  g748(.A1(new_n1172), .A2(new_n967), .A3(new_n1173), .ZN(G225));
endmodule


