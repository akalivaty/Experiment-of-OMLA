

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810;

  INV_X2 U379 ( .A(G146), .ZN(n536) );
  AND2_X1 U380 ( .A1(n454), .A2(n466), .ZN(n361) );
  INV_X1 U381 ( .A(G953), .ZN(n532) );
  AND2_X2 U382 ( .A1(n367), .A2(n532), .ZN(n718) );
  NAND2_X2 U383 ( .A1(n409), .A2(n408), .ZN(n741) );
  NOR2_X2 U384 ( .A1(n395), .A2(n392), .ZN(n386) );
  AND2_X2 U385 ( .A1(n723), .A2(n722), .ZN(n469) );
  NAND2_X2 U386 ( .A1(n361), .A2(n452), .ZN(n632) );
  XNOR2_X2 U387 ( .A(n421), .B(n588), .ZN(n607) );
  XNOR2_X2 U388 ( .A(n609), .B(n608), .ZN(n657) );
  NAND2_X1 U389 ( .A1(n445), .A2(n444), .ZN(n443) );
  NAND2_X1 U390 ( .A1(n470), .A2(n672), .ZN(n468) );
  AND2_X1 U391 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U392 ( .A1(n677), .A2(n774), .ZN(n798) );
  AND2_X1 U393 ( .A1(n485), .A2(n484), .ZN(n483) );
  AND2_X1 U394 ( .A1(n665), .A2(n664), .ZN(n496) );
  NAND2_X1 U395 ( .A1(n741), .A2(n720), .ZN(n662) );
  XNOR2_X1 U396 ( .A(n636), .B(n635), .ZN(n807) );
  XNOR2_X1 U397 ( .A(n462), .B(KEYINPUT32), .ZN(n720) );
  XNOR2_X1 U398 ( .A(n648), .B(n647), .ZN(n769) );
  NAND2_X1 U399 ( .A1(n434), .A2(n431), .ZN(n641) );
  XNOR2_X1 U400 ( .A(n734), .B(n733), .ZN(n735) );
  XNOR2_X1 U401 ( .A(n547), .B(n482), .ZN(n797) );
  INV_X1 U402 ( .A(n785), .ZN(n444) );
  INV_X1 U403 ( .A(KEYINPUT69), .ZN(n499) );
  BUF_X1 U404 ( .A(n742), .Z(n781) );
  XNOR2_X2 U405 ( .A(n384), .B(n479), .ZN(n739) );
  XNOR2_X2 U406 ( .A(n686), .B(n510), .ZN(n654) );
  NOR2_X1 U407 ( .A1(n656), .A2(KEYINPUT101), .ZN(n417) );
  XNOR2_X2 U408 ( .A(n509), .B(n508), .ZN(n686) );
  OR2_X1 U409 ( .A1(n775), .A2(n427), .ZN(n426) );
  NAND2_X1 U410 ( .A1(n428), .A2(n512), .ZN(n427) );
  INV_X1 U411 ( .A(n478), .ZN(n428) );
  AND2_X1 U412 ( .A1(n398), .A2(n430), .ZN(n429) );
  NAND2_X1 U413 ( .A1(n775), .A2(n478), .ZN(n398) );
  NAND2_X1 U414 ( .A1(n359), .A2(n378), .ZN(n611) );
  NOR2_X1 U415 ( .A1(n646), .A2(n439), .ZN(n472) );
  NAND2_X1 U416 ( .A1(n423), .A2(n437), .ZN(n596) );
  AND2_X1 U417 ( .A1(n703), .A2(n632), .ZN(n437) );
  XNOR2_X1 U418 ( .A(n498), .B(KEYINPUT71), .ZN(n482) );
  INV_X1 U419 ( .A(n497), .ZN(n498) );
  XNOR2_X1 U420 ( .A(G131), .B(G134), .ZN(n497) );
  XNOR2_X1 U421 ( .A(G137), .B(G140), .ZN(n537) );
  XNOR2_X1 U422 ( .A(n502), .B(n501), .ZN(n572) );
  INV_X1 U423 ( .A(KEYINPUT75), .ZN(n501) );
  NOR2_X1 U424 ( .A1(G953), .A2(G237), .ZN(n502) );
  INV_X1 U425 ( .A(G107), .ZN(n522) );
  OR2_X1 U426 ( .A1(n657), .A2(KEYINPUT33), .ZN(n475) );
  INV_X1 U427 ( .A(KEYINPUT84), .ZN(n455) );
  AND2_X1 U428 ( .A1(n625), .A2(KEYINPUT33), .ZN(n446) );
  INV_X1 U429 ( .A(KEYINPUT30), .ZN(n449) );
  NOR2_X1 U430 ( .A1(n630), .A2(n373), .ZN(n518) );
  AND2_X1 U431 ( .A1(n375), .A2(n374), .ZN(n373) );
  INV_X1 U432 ( .A(G900), .ZN(n374) );
  NAND2_X1 U433 ( .A1(n589), .A2(n360), .ZN(n466) );
  AND2_X1 U434 ( .A1(n436), .A2(n435), .ZN(n434) );
  NAND2_X1 U435 ( .A1(n433), .A2(n512), .ZN(n432) );
  INV_X1 U436 ( .A(KEYINPUT0), .ZN(n633) );
  XNOR2_X1 U437 ( .A(n481), .B(n480), .ZN(n479) );
  NAND2_X1 U438 ( .A1(n572), .A2(G210), .ZN(n480) );
  XNOR2_X1 U439 ( .A(n505), .B(n507), .ZN(n481) );
  XNOR2_X1 U440 ( .A(G119), .B(G110), .ZN(n548) );
  XNOR2_X1 U441 ( .A(n548), .B(n460), .ZN(n459) );
  XNOR2_X1 U442 ( .A(G128), .B(KEYINPUT24), .ZN(n460) );
  XNOR2_X1 U443 ( .A(n531), .B(KEYINPUT23), .ZN(n458) );
  INV_X1 U444 ( .A(KEYINPUT91), .ZN(n531) );
  XNOR2_X1 U445 ( .A(n586), .B(n585), .ZN(n695) );
  XNOR2_X1 U446 ( .A(n584), .B(KEYINPUT107), .ZN(n585) );
  INV_X1 U447 ( .A(KEYINPUT105), .ZN(n456) );
  INV_X1 U448 ( .A(KEYINPUT102), .ZN(n411) );
  NAND2_X1 U449 ( .A1(n401), .A2(n399), .ZN(n400) );
  NAND2_X1 U450 ( .A1(n425), .A2(KEYINPUT93), .ZN(n402) );
  BUF_X1 U451 ( .A(n686), .Z(n420) );
  XNOR2_X1 U452 ( .A(n539), .B(n362), .ZN(n461) );
  XNOR2_X1 U453 ( .A(G469), .B(n529), .ZN(n478) );
  AND2_X1 U454 ( .A1(n494), .A2(n492), .ZN(n491) );
  NAND2_X1 U455 ( .A1(n490), .A2(n357), .ZN(n484) );
  INV_X1 U456 ( .A(G237), .ZN(n511) );
  XNOR2_X1 U457 ( .A(n377), .B(n376), .ZN(n375) );
  INV_X1 U458 ( .A(KEYINPUT103), .ZN(n376) );
  NOR2_X1 U459 ( .A1(n627), .A2(n532), .ZN(n377) );
  NAND2_X1 U460 ( .A1(n358), .A2(n641), .ZN(n404) );
  INV_X1 U461 ( .A(n461), .ZN(n433) );
  NAND2_X1 U462 ( .A1(n461), .A2(G902), .ZN(n435) );
  XNOR2_X1 U463 ( .A(G137), .B(G119), .ZN(n503) );
  NAND2_X1 U464 ( .A1(G234), .A2(G237), .ZN(n514) );
  XNOR2_X1 U465 ( .A(n379), .B(KEYINPUT87), .ZN(n515) );
  INV_X1 U466 ( .A(KEYINPUT14), .ZN(n379) );
  NOR2_X1 U467 ( .A1(n442), .A2(n441), .ZN(n665) );
  NOR2_X1 U468 ( .A1(n807), .A2(n666), .ZN(n442) );
  INV_X1 U469 ( .A(n747), .ZN(n418) );
  NAND2_X1 U470 ( .A1(n700), .A2(n699), .ZN(n704) );
  XNOR2_X1 U471 ( .A(n620), .B(KEYINPUT38), .ZN(n700) );
  INV_X1 U472 ( .A(KEYINPUT28), .ZN(n382) );
  NOR2_X1 U473 ( .A1(n611), .A2(n637), .ZN(n438) );
  NAND2_X1 U474 ( .A1(n365), .A2(n655), .ZN(n416) );
  INV_X1 U475 ( .A(n429), .ZN(n425) );
  NAND2_X1 U476 ( .A1(n404), .A2(KEYINPUT93), .ZN(n403) );
  XNOR2_X1 U477 ( .A(G122), .B(G134), .ZN(n563) );
  XNOR2_X1 U478 ( .A(G143), .B(G140), .ZN(n573) );
  XNOR2_X1 U479 ( .A(n384), .B(n528), .ZN(n775) );
  XOR2_X1 U480 ( .A(G104), .B(G110), .Z(n526) );
  XNOR2_X1 U481 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n542) );
  NAND2_X1 U482 ( .A1(n393), .A2(n392), .ZN(n387) );
  NAND2_X1 U483 ( .A1(n476), .A2(n473), .ZN(n393) );
  XNOR2_X1 U484 ( .A(n540), .B(KEYINPUT76), .ZN(n597) );
  AND2_X1 U485 ( .A1(n649), .A2(n359), .ZN(n451) );
  NAND2_X1 U486 ( .A1(n453), .A2(n364), .ZN(n452) );
  XNOR2_X1 U487 ( .A(n740), .B(n371), .ZN(n445) );
  XNOR2_X1 U488 ( .A(n464), .B(n463), .ZN(n791) );
  XNOR2_X1 U489 ( .A(n548), .B(KEYINPUT16), .ZN(n463) );
  XNOR2_X1 U490 ( .A(n459), .B(n458), .ZN(n535) );
  INV_X1 U491 ( .A(n698), .ZN(n397) );
  XNOR2_X1 U492 ( .A(n422), .B(n587), .ZN(n810) );
  NAND2_X1 U493 ( .A1(n695), .A2(n423), .ZN(n422) );
  XNOR2_X1 U494 ( .A(n424), .B(n582), .ZN(n808) );
  OR2_X1 U495 ( .A1(n691), .A2(n646), .ZN(n648) );
  NAND2_X1 U496 ( .A1(n412), .A2(n410), .ZN(n409) );
  NAND2_X1 U497 ( .A1(n414), .A2(KEYINPUT102), .ZN(n408) );
  NAND2_X1 U498 ( .A1(n417), .A2(n411), .ZN(n410) );
  NAND2_X1 U499 ( .A1(n440), .A2(n651), .ZN(n752) );
  AND2_X1 U500 ( .A1(n493), .A2(n617), .ZN(n357) );
  AND2_X1 U501 ( .A1(n426), .A2(n684), .ZN(n358) );
  XOR2_X1 U502 ( .A(n518), .B(KEYINPUT78), .Z(n359) );
  XNOR2_X1 U503 ( .A(KEYINPUT68), .B(KEYINPUT19), .ZN(n360) );
  NAND2_X1 U504 ( .A1(n471), .A2(n476), .ZN(n698) );
  NAND2_X1 U505 ( .A1(n474), .A2(n477), .ZN(n473) );
  XOR2_X1 U506 ( .A(KEYINPUT92), .B(KEYINPUT25), .Z(n362) );
  XNOR2_X1 U507 ( .A(n380), .B(n456), .ZN(n592) );
  INV_X1 U508 ( .A(n592), .ZN(n423) );
  AND2_X1 U509 ( .A1(n446), .A2(n659), .ZN(n363) );
  BUF_X1 U510 ( .A(n590), .Z(n620) );
  NOR2_X1 U511 ( .A1(n589), .A2(n360), .ZN(n364) );
  OR2_X1 U512 ( .A1(n682), .A2(KEYINPUT101), .ZN(n365) );
  AND2_X1 U513 ( .A1(n682), .A2(KEYINPUT101), .ZN(n366) );
  AND2_X1 U514 ( .A1(n717), .A2(n495), .ZN(n367) );
  INV_X1 U515 ( .A(n641), .ZN(n378) );
  AND2_X1 U516 ( .A1(n661), .A2(n660), .ZN(n368) );
  AND2_X1 U517 ( .A1(n403), .A2(n402), .ZN(n369) );
  INV_X1 U518 ( .A(KEYINPUT33), .ZN(n477) );
  AND2_X1 U519 ( .A1(n397), .A2(n695), .ZN(n370) );
  INV_X1 U520 ( .A(KEYINPUT34), .ZN(n392) );
  XNOR2_X1 U521 ( .A(KEYINPUT62), .B(n739), .ZN(n371) );
  XNOR2_X1 U522 ( .A(KEYINPUT86), .B(KEYINPUT63), .ZN(n372) );
  XNOR2_X1 U523 ( .A(n557), .B(n556), .ZN(n622) );
  NAND2_X2 U524 ( .A1(n469), .A2(n468), .ZN(n467) );
  NAND2_X1 U525 ( .A1(n483), .A2(n486), .ZN(n677) );
  NAND2_X1 U526 ( .A1(n369), .A2(n400), .ZN(n649) );
  NAND2_X1 U527 ( .A1(n656), .A2(n366), .ZN(n396) );
  XNOR2_X2 U528 ( .A(n640), .B(n639), .ZN(n656) );
  NAND2_X1 U529 ( .A1(n381), .A2(n457), .ZN(n380) );
  XNOR2_X1 U530 ( .A(n383), .B(n382), .ZN(n381) );
  NAND2_X1 U531 ( .A1(n654), .A2(n699), .ZN(n513) );
  NAND2_X1 U532 ( .A1(n438), .A2(n654), .ZN(n383) );
  XNOR2_X2 U533 ( .A(n797), .B(n500), .ZN(n384) );
  INV_X1 U534 ( .A(n472), .ZN(n391) );
  NAND2_X1 U535 ( .A1(n385), .A2(n472), .ZN(n390) );
  NAND2_X1 U536 ( .A1(n476), .A2(n386), .ZN(n385) );
  NAND2_X1 U537 ( .A1(n388), .A2(n387), .ZN(n394) );
  NAND2_X1 U538 ( .A1(n390), .A2(n389), .ZN(n388) );
  NAND2_X1 U539 ( .A1(n391), .A2(KEYINPUT34), .ZN(n389) );
  NAND2_X1 U540 ( .A1(n394), .A2(n634), .ZN(n636) );
  INV_X1 U541 ( .A(n473), .ZN(n395) );
  NAND2_X1 U542 ( .A1(n415), .A2(n396), .ZN(n414) );
  NAND2_X1 U543 ( .A1(n413), .A2(n396), .ZN(n407) );
  OR2_X1 U544 ( .A1(n786), .A2(KEYINPUT2), .ZN(n673) );
  NAND2_X1 U545 ( .A1(n678), .A2(n786), .ZN(n723) );
  NAND2_X1 U546 ( .A1(n405), .A2(n786), .ZN(n470) );
  XNOR2_X2 U547 ( .A(n671), .B(KEYINPUT45), .ZN(n786) );
  INV_X1 U548 ( .A(n700), .ZN(n583) );
  NOR2_X1 U549 ( .A1(n702), .A2(n704), .ZN(n586) );
  INV_X1 U550 ( .A(n404), .ZN(n399) );
  NOR2_X1 U551 ( .A1(n425), .A2(KEYINPUT93), .ZN(n401) );
  INV_X1 U552 ( .A(n798), .ZN(n405) );
  NAND2_X1 U553 ( .A1(n407), .A2(n406), .ZN(n412) );
  INV_X1 U554 ( .A(n417), .ZN(n406) );
  NOR2_X1 U555 ( .A1(n416), .A2(KEYINPUT102), .ZN(n413) );
  INV_X1 U556 ( .A(n416), .ZN(n415) );
  NAND2_X1 U557 ( .A1(n650), .A2(n638), .ZN(n640) );
  NAND2_X1 U558 ( .A1(n419), .A2(n418), .ZN(n441) );
  XNOR2_X1 U559 ( .A(n653), .B(KEYINPUT98), .ZN(n419) );
  XNOR2_X1 U560 ( .A(n513), .B(n449), .ZN(n448) );
  NAND2_X1 U561 ( .A1(n808), .A2(n810), .ZN(n421) );
  NAND2_X1 U562 ( .A1(n622), .A2(n762), .ZN(n424) );
  NAND2_X1 U563 ( .A1(n429), .A2(n426), .ZN(n609) );
  NAND2_X1 U564 ( .A1(n478), .A2(G902), .ZN(n430) );
  OR2_X1 U565 ( .A1(n782), .A2(n432), .ZN(n431) );
  NAND2_X1 U566 ( .A1(n782), .A2(n461), .ZN(n436) );
  XNOR2_X1 U567 ( .A(n538), .B(n796), .ZN(n782) );
  NOR2_X1 U568 ( .A1(n592), .A2(n591), .ZN(n763) );
  INV_X1 U569 ( .A(n475), .ZN(n439) );
  INV_X1 U570 ( .A(n646), .ZN(n440) );
  XNOR2_X1 U571 ( .A(n443), .B(n372), .ZN(G57) );
  XNOR2_X1 U572 ( .A(n447), .B(n546), .ZN(n551) );
  XNOR2_X1 U573 ( .A(n545), .B(n547), .ZN(n447) );
  NAND2_X1 U574 ( .A1(n451), .A2(n448), .ZN(n540) );
  NAND2_X1 U575 ( .A1(n670), .A2(n496), .ZN(n671) );
  XNOR2_X1 U576 ( .A(n662), .B(n455), .ZN(n668) );
  XNOR2_X2 U577 ( .A(n450), .B(n633), .ZN(n650) );
  NAND2_X1 U578 ( .A1(n632), .A2(n631), .ZN(n450) );
  XNOR2_X1 U579 ( .A(n559), .B(n549), .ZN(n550) );
  XNOR2_X2 U580 ( .A(KEYINPUT73), .B(KEYINPUT3), .ZN(n549) );
  XNOR2_X2 U581 ( .A(G116), .B(G107), .ZN(n559) );
  INV_X1 U582 ( .A(n590), .ZN(n453) );
  NAND2_X1 U583 ( .A1(n590), .A2(n360), .ZN(n454) );
  XNOR2_X2 U584 ( .A(n555), .B(n554), .ZN(n590) );
  NAND2_X1 U585 ( .A1(n607), .A2(n494), .ZN(n488) );
  INV_X1 U586 ( .A(n609), .ZN(n457) );
  NAND2_X1 U587 ( .A1(n656), .A2(n368), .ZN(n462) );
  XNOR2_X1 U588 ( .A(n550), .B(n569), .ZN(n464) );
  XNOR2_X2 U589 ( .A(n465), .B(G104), .ZN(n569) );
  XNOR2_X2 U590 ( .A(G122), .B(G113), .ZN(n465) );
  XNOR2_X2 U591 ( .A(n499), .B(G101), .ZN(n543) );
  XNOR2_X2 U592 ( .A(n536), .B(G125), .ZN(n544) );
  XNOR2_X2 U593 ( .A(n467), .B(KEYINPUT65), .ZN(n742) );
  AND2_X1 U594 ( .A1(n473), .A2(n475), .ZN(n471) );
  AND2_X1 U595 ( .A1(n657), .A2(n625), .ZN(n645) );
  NAND2_X1 U596 ( .A1(n625), .A2(n659), .ZN(n474) );
  NAND2_X1 U597 ( .A1(n363), .A2(n657), .ZN(n476) );
  XNOR2_X2 U598 ( .A(n561), .B(KEYINPUT4), .ZN(n547) );
  NAND2_X1 U599 ( .A1(n488), .A2(n357), .ZN(n485) );
  NAND2_X1 U600 ( .A1(n607), .A2(n487), .ZN(n486) );
  AND2_X1 U601 ( .A1(n606), .A2(n489), .ZN(n487) );
  AND2_X1 U602 ( .A1(n491), .A2(n493), .ZN(n489) );
  INV_X1 U603 ( .A(n606), .ZN(n490) );
  INV_X1 U604 ( .A(n617), .ZN(n492) );
  INV_X1 U605 ( .A(n721), .ZN(n493) );
  INV_X1 U606 ( .A(n772), .ZN(n494) );
  XOR2_X1 U607 ( .A(KEYINPUT121), .B(n716), .Z(n495) );
  AND2_X1 U608 ( .A1(n807), .A2(n666), .ZN(n667) );
  XNOR2_X1 U609 ( .A(n669), .B(KEYINPUT74), .ZN(n670) );
  XNOR2_X1 U610 ( .A(n523), .B(n522), .ZN(n525) );
  XNOR2_X1 U611 ( .A(n525), .B(n524), .ZN(n527) );
  INV_X1 U612 ( .A(n681), .ZN(n625) );
  XNOR2_X1 U613 ( .A(n535), .B(n534), .ZN(n538) );
  INV_X1 U614 ( .A(KEYINPUT2), .ZN(n672) );
  XNOR2_X2 U615 ( .A(G143), .B(G128), .ZN(n561) );
  XNOR2_X1 U616 ( .A(n543), .B(G146), .ZN(n500) );
  XOR2_X1 U617 ( .A(G116), .B(G113), .Z(n504) );
  XNOR2_X1 U618 ( .A(n504), .B(n503), .ZN(n505) );
  INV_X1 U619 ( .A(KEYINPUT5), .ZN(n506) );
  XNOR2_X1 U620 ( .A(n549), .B(n506), .ZN(n507) );
  INV_X1 U621 ( .A(G902), .ZN(n512) );
  NAND2_X1 U622 ( .A1(n739), .A2(n512), .ZN(n509) );
  INV_X1 U623 ( .A(G472), .ZN(n508) );
  INV_X1 U624 ( .A(KEYINPUT100), .ZN(n510) );
  NAND2_X1 U625 ( .A1(n512), .A2(n511), .ZN(n553) );
  NAND2_X1 U626 ( .A1(n553), .A2(G214), .ZN(n699) );
  XNOR2_X1 U627 ( .A(n515), .B(n514), .ZN(n517) );
  NAND2_X1 U628 ( .A1(n517), .A2(G952), .ZN(n516) );
  XNOR2_X1 U629 ( .A(n516), .B(KEYINPUT88), .ZN(n714) );
  NOR2_X1 U630 ( .A1(n714), .A2(G953), .ZN(n630) );
  NAND2_X1 U631 ( .A1(G902), .A2(n517), .ZN(n627) );
  XNOR2_X1 U632 ( .A(G902), .B(KEYINPUT15), .ZN(n552) );
  NAND2_X1 U633 ( .A1(G234), .A2(n552), .ZN(n519) );
  XNOR2_X1 U634 ( .A(KEYINPUT20), .B(n519), .ZN(n530) );
  NAND2_X1 U635 ( .A1(n530), .A2(G221), .ZN(n521) );
  INV_X1 U636 ( .A(KEYINPUT21), .ZN(n520) );
  XNOR2_X1 U637 ( .A(n521), .B(n520), .ZN(n684) );
  INV_X1 U638 ( .A(n684), .ZN(n637) );
  NAND2_X1 U639 ( .A1(G227), .A2(n532), .ZN(n523) );
  INV_X1 U640 ( .A(n537), .ZN(n524) );
  XNOR2_X1 U641 ( .A(n527), .B(n526), .ZN(n528) );
  INV_X1 U642 ( .A(KEYINPUT72), .ZN(n529) );
  NAND2_X1 U643 ( .A1(n530), .A2(G217), .ZN(n539) );
  NAND2_X1 U644 ( .A1(G234), .A2(n532), .ZN(n533) );
  XOR2_X1 U645 ( .A(KEYINPUT8), .B(n533), .Z(n558) );
  NAND2_X1 U646 ( .A1(G221), .A2(n558), .ZN(n534) );
  XOR2_X1 U647 ( .A(KEYINPUT10), .B(n544), .Z(n571) );
  XNOR2_X1 U648 ( .A(n537), .B(n571), .ZN(n796) );
  NAND2_X1 U649 ( .A1(n532), .A2(G224), .ZN(n541) );
  XNOR2_X1 U650 ( .A(n542), .B(n541), .ZN(n546) );
  XNOR2_X1 U651 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U652 ( .A(n551), .B(n791), .ZN(n726) );
  INV_X1 U653 ( .A(n552), .ZN(n722) );
  OR2_X2 U654 ( .A1(n726), .A2(n722), .ZN(n555) );
  NAND2_X1 U655 ( .A1(n553), .A2(G210), .ZN(n554) );
  NOR2_X2 U656 ( .A1(n597), .A2(n583), .ZN(n557) );
  INV_X1 U657 ( .A(KEYINPUT39), .ZN(n556) );
  NAND2_X1 U658 ( .A1(G217), .A2(n558), .ZN(n560) );
  XNOR2_X1 U659 ( .A(n559), .B(n560), .ZN(n567) );
  XNOR2_X1 U660 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n562) );
  XNOR2_X1 U661 ( .A(n561), .B(n562), .ZN(n565) );
  XNOR2_X1 U662 ( .A(n563), .B(KEYINPUT96), .ZN(n564) );
  XNOR2_X1 U663 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U664 ( .A(n567), .B(n566), .ZN(n743) );
  NOR2_X1 U665 ( .A1(G902), .A2(n743), .ZN(n568) );
  XNOR2_X1 U666 ( .A(G478), .B(n568), .ZN(n599) );
  XNOR2_X1 U667 ( .A(n569), .B(G131), .ZN(n570) );
  XNOR2_X1 U668 ( .A(n571), .B(n570), .ZN(n579) );
  NAND2_X1 U669 ( .A1(G214), .A2(n572), .ZN(n576) );
  XOR2_X1 U670 ( .A(KEYINPUT12), .B(KEYINPUT95), .Z(n574) );
  XNOR2_X1 U671 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U672 ( .A(n576), .B(n575), .ZN(n577) );
  XOR2_X1 U673 ( .A(n577), .B(KEYINPUT11), .Z(n578) );
  XNOR2_X1 U674 ( .A(n579), .B(n578), .ZN(n734) );
  NOR2_X1 U675 ( .A1(G902), .A2(n734), .ZN(n581) );
  XNOR2_X1 U676 ( .A(KEYINPUT13), .B(G475), .ZN(n580) );
  XNOR2_X1 U677 ( .A(n581), .B(n580), .ZN(n593) );
  NAND2_X1 U678 ( .A1(n599), .A2(n593), .ZN(n766) );
  INV_X1 U679 ( .A(n766), .ZN(n762) );
  XNOR2_X1 U680 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n582) );
  XOR2_X1 U681 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n587) );
  INV_X1 U682 ( .A(n593), .ZN(n600) );
  NAND2_X1 U683 ( .A1(n600), .A2(n599), .ZN(n702) );
  XNOR2_X1 U684 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n584) );
  XOR2_X1 U685 ( .A(KEYINPUT46), .B(KEYINPUT64), .Z(n588) );
  INV_X1 U686 ( .A(n699), .ZN(n589) );
  INV_X1 U687 ( .A(n632), .ZN(n591) );
  NOR2_X1 U688 ( .A1(n593), .A2(n599), .ZN(n757) );
  NOR2_X1 U689 ( .A1(n757), .A2(n762), .ZN(n594) );
  XNOR2_X1 U690 ( .A(n594), .B(KEYINPUT97), .ZN(n703) );
  XNOR2_X1 U691 ( .A(KEYINPUT70), .B(KEYINPUT47), .ZN(n595) );
  NOR2_X1 U692 ( .A1(n596), .A2(n595), .ZN(n605) );
  NAND2_X1 U693 ( .A1(KEYINPUT47), .A2(n596), .ZN(n602) );
  NOR2_X1 U694 ( .A1(n597), .A2(n620), .ZN(n598) );
  XNOR2_X1 U695 ( .A(n598), .B(KEYINPUT104), .ZN(n601) );
  NOR2_X1 U696 ( .A1(n600), .A2(n599), .ZN(n634) );
  NAND2_X1 U697 ( .A1(n601), .A2(n634), .ZN(n761) );
  NAND2_X1 U698 ( .A1(n602), .A2(n761), .ZN(n603) );
  XNOR2_X1 U699 ( .A(KEYINPUT80), .B(n603), .ZN(n604) );
  NOR2_X1 U700 ( .A1(n605), .A2(n604), .ZN(n606) );
  INV_X1 U701 ( .A(KEYINPUT1), .ZN(n608) );
  INV_X1 U702 ( .A(n657), .ZN(n682) );
  NAND2_X1 U703 ( .A1(n699), .A2(n684), .ZN(n610) );
  NOR2_X1 U704 ( .A1(n611), .A2(n610), .ZN(n614) );
  XNOR2_X1 U705 ( .A(n686), .B(KEYINPUT6), .ZN(n659) );
  INV_X1 U706 ( .A(n659), .ZN(n612) );
  NOR2_X1 U707 ( .A1(n612), .A2(n766), .ZN(n613) );
  NAND2_X1 U708 ( .A1(n614), .A2(n613), .ZN(n618) );
  NOR2_X1 U709 ( .A1(n618), .A2(n620), .ZN(n615) );
  XOR2_X1 U710 ( .A(KEYINPUT36), .B(n615), .Z(n616) );
  NOR2_X1 U711 ( .A1(n682), .A2(n616), .ZN(n772) );
  XNOR2_X1 U712 ( .A(KEYINPUT83), .B(KEYINPUT48), .ZN(n617) );
  NOR2_X1 U713 ( .A1(n657), .A2(n618), .ZN(n619) );
  XNOR2_X1 U714 ( .A(n619), .B(KEYINPUT43), .ZN(n621) );
  NOR2_X1 U715 ( .A1(n621), .A2(n453), .ZN(n721) );
  BUF_X1 U716 ( .A(n622), .Z(n623) );
  NAND2_X1 U717 ( .A1(n623), .A2(n757), .ZN(n774) );
  AND2_X1 U718 ( .A1(n672), .A2(n798), .ZN(n624) );
  XNOR2_X1 U719 ( .A(n624), .B(KEYINPUT81), .ZN(n674) );
  NAND2_X1 U720 ( .A1(n641), .A2(n684), .ZN(n681) );
  NOR2_X1 U721 ( .A1(G898), .A2(n532), .ZN(n626) );
  XNOR2_X1 U722 ( .A(KEYINPUT89), .B(n626), .ZN(n792) );
  NOR2_X1 U723 ( .A1(n627), .A2(n792), .ZN(n628) );
  XNOR2_X1 U724 ( .A(n628), .B(KEYINPUT90), .ZN(n629) );
  OR2_X1 U725 ( .A1(n630), .A2(n629), .ZN(n631) );
  INV_X1 U726 ( .A(n650), .ZN(n646) );
  INV_X1 U727 ( .A(KEYINPUT35), .ZN(n635) );
  INV_X1 U728 ( .A(KEYINPUT44), .ZN(n666) );
  NOR2_X1 U729 ( .A1(n702), .A2(n637), .ZN(n638) );
  INV_X1 U730 ( .A(KEYINPUT22), .ZN(n639) );
  OR2_X1 U731 ( .A1(n657), .A2(n378), .ZN(n642) );
  NOR2_X1 U732 ( .A1(n659), .A2(n642), .ZN(n643) );
  AND2_X1 U733 ( .A1(n656), .A2(n643), .ZN(n747) );
  INV_X1 U734 ( .A(n420), .ZN(n644) );
  NAND2_X1 U735 ( .A1(n645), .A2(n644), .ZN(n691) );
  XOR2_X1 U736 ( .A(KEYINPUT31), .B(KEYINPUT94), .Z(n647) );
  AND2_X1 U737 ( .A1(n420), .A2(n649), .ZN(n651) );
  NAND2_X1 U738 ( .A1(n769), .A2(n752), .ZN(n652) );
  NAND2_X1 U739 ( .A1(n652), .A2(n703), .ZN(n653) );
  NOR2_X1 U740 ( .A1(n654), .A2(n641), .ZN(n655) );
  NAND2_X1 U741 ( .A1(n657), .A2(n378), .ZN(n658) );
  XNOR2_X1 U742 ( .A(n658), .B(KEYINPUT99), .ZN(n661) );
  XNOR2_X1 U743 ( .A(n659), .B(KEYINPUT77), .ZN(n660) );
  NAND2_X1 U744 ( .A1(n662), .A2(KEYINPUT44), .ZN(n663) );
  XNOR2_X1 U745 ( .A(n663), .B(KEYINPUT66), .ZN(n664) );
  NAND2_X1 U746 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U747 ( .A1(n674), .A2(n673), .ZN(n679) );
  NAND2_X1 U748 ( .A1(n774), .A2(KEYINPUT2), .ZN(n675) );
  XNOR2_X1 U749 ( .A(n675), .B(KEYINPUT79), .ZN(n676) );
  NAND2_X1 U750 ( .A1(n679), .A2(n723), .ZN(n680) );
  XNOR2_X1 U751 ( .A(n680), .B(KEYINPUT82), .ZN(n717) );
  NAND2_X1 U752 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U753 ( .A(n683), .B(KEYINPUT50), .ZN(n690) );
  NOR2_X1 U754 ( .A1(n641), .A2(n684), .ZN(n685) );
  XNOR2_X1 U755 ( .A(n685), .B(KEYINPUT49), .ZN(n687) );
  NAND2_X1 U756 ( .A1(n687), .A2(n420), .ZN(n688) );
  XNOR2_X1 U757 ( .A(KEYINPUT117), .B(n688), .ZN(n689) );
  NAND2_X1 U758 ( .A1(n690), .A2(n689), .ZN(n692) );
  NAND2_X1 U759 ( .A1(n692), .A2(n691), .ZN(n694) );
  XOR2_X1 U760 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n693) );
  XNOR2_X1 U761 ( .A(n694), .B(n693), .ZN(n696) );
  NAND2_X1 U762 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U763 ( .A(n697), .B(KEYINPUT119), .ZN(n711) );
  NOR2_X1 U764 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U765 ( .A1(n702), .A2(n701), .ZN(n707) );
  INV_X1 U766 ( .A(n703), .ZN(n705) );
  NOR2_X1 U767 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U768 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U769 ( .A(KEYINPUT120), .B(n708), .ZN(n709) );
  NOR2_X1 U770 ( .A1(n698), .A2(n709), .ZN(n710) );
  NOR2_X1 U771 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U772 ( .A(n712), .B(KEYINPUT52), .ZN(n713) );
  NOR2_X1 U773 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U774 ( .A1(n715), .A2(n370), .ZN(n716) );
  XNOR2_X1 U775 ( .A(n718), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U776 ( .A(G119), .B(KEYINPUT127), .Z(n719) );
  XNOR2_X1 U777 ( .A(n720), .B(n719), .ZN(G21) );
  XOR2_X1 U778 ( .A(G140), .B(n721), .Z(G42) );
  NAND2_X1 U779 ( .A1(n742), .A2(G210), .ZN(n728) );
  XNOR2_X1 U780 ( .A(KEYINPUT85), .B(KEYINPUT54), .ZN(n724) );
  XNOR2_X1 U781 ( .A(n724), .B(KEYINPUT55), .ZN(n725) );
  XNOR2_X1 U782 ( .A(n726), .B(n725), .ZN(n727) );
  XNOR2_X1 U783 ( .A(n728), .B(n727), .ZN(n730) );
  INV_X1 U784 ( .A(G952), .ZN(n729) );
  AND2_X1 U785 ( .A1(n729), .A2(G953), .ZN(n785) );
  NOR2_X2 U786 ( .A1(n730), .A2(n785), .ZN(n731) );
  XNOR2_X1 U787 ( .A(n731), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U788 ( .A1(n742), .A2(G475), .ZN(n736) );
  XNOR2_X1 U789 ( .A(KEYINPUT67), .B(KEYINPUT123), .ZN(n732) );
  XOR2_X1 U790 ( .A(n732), .B(KEYINPUT59), .Z(n733) );
  XNOR2_X1 U791 ( .A(n736), .B(n735), .ZN(n737) );
  NOR2_X2 U792 ( .A1(n737), .A2(n785), .ZN(n738) );
  XNOR2_X1 U793 ( .A(n738), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U794 ( .A1(n742), .A2(G472), .ZN(n740) );
  XNOR2_X1 U795 ( .A(n741), .B(G110), .ZN(G12) );
  NAND2_X1 U796 ( .A1(n781), .A2(G478), .ZN(n745) );
  XNOR2_X1 U797 ( .A(n743), .B(KEYINPUT124), .ZN(n744) );
  XNOR2_X1 U798 ( .A(n745), .B(n744), .ZN(n746) );
  NOR2_X1 U799 ( .A1(n746), .A2(n785), .ZN(G63) );
  XOR2_X1 U800 ( .A(G101), .B(n747), .Z(G3) );
  NOR2_X1 U801 ( .A1(n752), .A2(n766), .ZN(n748) );
  XOR2_X1 U802 ( .A(KEYINPUT110), .B(n748), .Z(n749) );
  XNOR2_X1 U803 ( .A(G104), .B(n749), .ZN(G6) );
  XOR2_X1 U804 ( .A(KEYINPUT113), .B(KEYINPUT112), .Z(n751) );
  XNOR2_X1 U805 ( .A(KEYINPUT111), .B(KEYINPUT27), .ZN(n750) );
  XNOR2_X1 U806 ( .A(n751), .B(n750), .ZN(n756) );
  INV_X1 U807 ( .A(n757), .ZN(n768) );
  NOR2_X1 U808 ( .A1(n752), .A2(n768), .ZN(n754) );
  XNOR2_X1 U809 ( .A(G107), .B(KEYINPUT26), .ZN(n753) );
  XNOR2_X1 U810 ( .A(n754), .B(n753), .ZN(n755) );
  XOR2_X1 U811 ( .A(n756), .B(n755), .Z(G9) );
  XOR2_X1 U812 ( .A(KEYINPUT114), .B(KEYINPUT29), .Z(n759) );
  NAND2_X1 U813 ( .A1(n763), .A2(n757), .ZN(n758) );
  XNOR2_X1 U814 ( .A(n759), .B(n758), .ZN(n760) );
  XNOR2_X1 U815 ( .A(G128), .B(n760), .ZN(G30) );
  XNOR2_X1 U816 ( .A(G143), .B(n761), .ZN(G45) );
  XOR2_X1 U817 ( .A(G146), .B(KEYINPUT115), .Z(n765) );
  NAND2_X1 U818 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U819 ( .A(n765), .B(n764), .ZN(G48) );
  NOR2_X1 U820 ( .A1(n769), .A2(n766), .ZN(n767) );
  XOR2_X1 U821 ( .A(G113), .B(n767), .Z(G15) );
  NOR2_X1 U822 ( .A1(n769), .A2(n768), .ZN(n770) );
  XOR2_X1 U823 ( .A(KEYINPUT116), .B(n770), .Z(n771) );
  XNOR2_X1 U824 ( .A(G116), .B(n771), .ZN(G18) );
  XNOR2_X1 U825 ( .A(G125), .B(n772), .ZN(n773) );
  XNOR2_X1 U826 ( .A(n773), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U827 ( .A(G134), .B(n774), .ZN(G36) );
  NAND2_X1 U828 ( .A1(n781), .A2(G469), .ZN(n779) );
  XOR2_X1 U829 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n777) );
  XNOR2_X1 U830 ( .A(n775), .B(KEYINPUT122), .ZN(n776) );
  XNOR2_X1 U831 ( .A(n777), .B(n776), .ZN(n778) );
  XNOR2_X1 U832 ( .A(n779), .B(n778), .ZN(n780) );
  NOR2_X1 U833 ( .A1(n785), .A2(n780), .ZN(G54) );
  NAND2_X1 U834 ( .A1(n781), .A2(G217), .ZN(n783) );
  XNOR2_X1 U835 ( .A(n783), .B(n782), .ZN(n784) );
  NOR2_X1 U836 ( .A1(n785), .A2(n784), .ZN(G66) );
  NAND2_X1 U837 ( .A1(n786), .A2(n532), .ZN(n790) );
  NAND2_X1 U838 ( .A1(G953), .A2(G224), .ZN(n787) );
  XNOR2_X1 U839 ( .A(KEYINPUT61), .B(n787), .ZN(n788) );
  NAND2_X1 U840 ( .A1(n788), .A2(G898), .ZN(n789) );
  NAND2_X1 U841 ( .A1(n790), .A2(n789), .ZN(n795) );
  XNOR2_X1 U842 ( .A(n791), .B(G101), .ZN(n793) );
  NAND2_X1 U843 ( .A1(n793), .A2(n792), .ZN(n794) );
  XOR2_X1 U844 ( .A(n795), .B(n794), .Z(G69) );
  XOR2_X1 U845 ( .A(n797), .B(n796), .Z(n801) );
  XOR2_X1 U846 ( .A(n801), .B(n798), .Z(n799) );
  NOR2_X1 U847 ( .A1(G953), .A2(n799), .ZN(n800) );
  XNOR2_X1 U848 ( .A(KEYINPUT125), .B(n800), .ZN(n805) );
  XNOR2_X1 U849 ( .A(G227), .B(n801), .ZN(n802) );
  NAND2_X1 U850 ( .A1(n802), .A2(G900), .ZN(n803) );
  NAND2_X1 U851 ( .A1(n803), .A2(G953), .ZN(n804) );
  NAND2_X1 U852 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U853 ( .A(n806), .B(KEYINPUT126), .ZN(G72) );
  XNOR2_X1 U854 ( .A(G122), .B(n807), .ZN(G24) );
  BUF_X1 U855 ( .A(n808), .Z(n809) );
  XNOR2_X1 U856 ( .A(G131), .B(n809), .ZN(G33) );
  XNOR2_X1 U857 ( .A(G137), .B(n810), .ZN(G39) );
endmodule

