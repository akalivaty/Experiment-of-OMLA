//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 0 0 0 0 1 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 1 0 0 0 0 1 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:52 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G13), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n209), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(KEYINPUT1), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G87), .A2(G250), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n225));
  AND4_X1   g0025(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  XOR2_X1   g0026(.A(KEYINPUT65), .B(G244), .Z(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G77), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n210), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n215), .B(new_n220), .C1(new_n221), .C2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n229), .A2(new_n221), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT66), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n230), .A2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT69), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G250), .ZN(new_n236));
  INV_X1    g0036(.A(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n239));
  XNOR2_X1  g0039(.A(G226), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n241), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n238), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT70), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  NAND2_X1  g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT71), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n218), .ZN(new_n257));
  NAND3_X1  g0057(.A1(KEYINPUT71), .A2(G33), .A3(G41), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G41), .ZN(new_n260));
  INV_X1    g0060(.A(G45), .ZN(new_n261));
  AOI21_X1  g0061(.A(G1), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n259), .A2(G274), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  INV_X1    g0064(.A(G97), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G226), .A2(G1698), .ZN(new_n267));
  INV_X1    g0067(.A(G232), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n267), .B1(new_n268), .B2(G1698), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT3), .B(G33), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n266), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n257), .A2(new_n254), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n263), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n262), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n259), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT76), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT76), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n259), .A2(new_n275), .A3(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n277), .A2(G238), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n274), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(KEYINPUT13), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT77), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT13), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n274), .A2(new_n284), .A3(new_n280), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n282), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n281), .A2(KEYINPUT77), .A3(KEYINPUT13), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n286), .A2(G169), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(KEYINPUT14), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT14), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n286), .A2(new_n290), .A3(G169), .A4(new_n287), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n282), .A2(G179), .A3(new_n285), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n289), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n218), .ZN(new_n295));
  NOR2_X1   g0095(.A1(G20), .A2(G33), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  OAI22_X1  g0097(.A1(new_n297), .A2(new_n201), .B1(new_n209), .B2(G68), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n209), .A2(G33), .ZN(new_n299));
  INV_X1    g0099(.A(G77), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n295), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n302), .B(KEYINPUT11), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT78), .B1(new_n304), .B2(G68), .ZN(new_n305));
  XOR2_X1   g0105(.A(new_n305), .B(KEYINPUT12), .Z(new_n306));
  INV_X1    g0106(.A(new_n304), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n307), .A2(new_n295), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n208), .A2(G20), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n308), .A2(G68), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n303), .A2(new_n306), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n293), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n286), .A2(G200), .A3(new_n287), .ZN(new_n314));
  INV_X1    g0114(.A(G190), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n315), .B1(new_n281), .B2(KEYINPUT13), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n311), .B1(new_n316), .B2(new_n285), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n313), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n201), .B1(new_n208), .B2(G20), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n308), .A2(new_n321), .B1(new_n201), .B2(new_n307), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT8), .B(G58), .ZN(new_n323));
  INV_X1    g0123(.A(G150), .ZN(new_n324));
  OAI22_X1  g0124(.A1(new_n323), .A2(new_n299), .B1(new_n324), .B2(new_n297), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n325), .B1(G20), .B2(new_n204), .ZN(new_n326));
  INV_X1    g0126(.A(new_n295), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n322), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  XNOR2_X1  g0128(.A(new_n328), .B(KEYINPUT9), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT10), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n276), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(G226), .ZN(new_n333));
  INV_X1    g0133(.A(G1698), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G222), .ZN(new_n335));
  INV_X1    g0135(.A(G223), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n270), .B(new_n335), .C1(new_n336), .C2(new_n334), .ZN(new_n337));
  INV_X1    g0137(.A(new_n272), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n337), .B(new_n338), .C1(G77), .C2(new_n270), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n333), .A2(new_n339), .A3(G190), .A4(new_n263), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT74), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n340), .B(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n333), .A2(new_n339), .A3(new_n263), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(G200), .ZN(new_n344));
  OR2_X1    g0144(.A1(new_n344), .A2(KEYINPUT73), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(KEYINPUT73), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n331), .A2(new_n342), .A3(new_n345), .A4(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n342), .A2(new_n329), .A3(new_n344), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT10), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(G169), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n343), .A2(new_n351), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n352), .B(new_n328), .C1(G179), .C2(new_n343), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n332), .A2(new_n227), .ZN(new_n354));
  NAND2_X1  g0154(.A1(G238), .A2(G1698), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n270), .B(new_n355), .C1(new_n268), .C2(G1698), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n356), .B(new_n338), .C1(G107), .C2(new_n270), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n354), .A2(new_n357), .A3(new_n263), .ZN(new_n358));
  OR2_X1    g0158(.A1(new_n358), .A2(G179), .ZN(new_n359));
  NAND2_X1  g0159(.A1(G20), .A2(G77), .ZN(new_n360));
  XNOR2_X1  g0160(.A(KEYINPUT15), .B(G87), .ZN(new_n361));
  OAI221_X1 g0161(.A(new_n360), .B1(new_n323), .B2(new_n297), .C1(new_n299), .C2(new_n361), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n362), .A2(new_n295), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n308), .A2(G77), .A3(new_n309), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(G77), .B2(new_n304), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n358), .A2(new_n351), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n359), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n358), .A2(G200), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n370), .B(new_n366), .C1(new_n315), .C2(new_n358), .ZN(new_n371));
  AND3_X1   g0171(.A1(new_n369), .A2(KEYINPUT72), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(KEYINPUT72), .B1(new_n369), .B2(new_n371), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n350), .A2(new_n353), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT75), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n350), .A2(new_n374), .A3(KEYINPUT75), .A4(new_n353), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n259), .A2(new_n275), .A3(G232), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n263), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(KEYINPUT79), .B1(new_n264), .B2(KEYINPUT3), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT79), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT3), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(new_n384), .A3(G33), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n264), .A2(KEYINPUT3), .ZN(new_n386));
  AND2_X1   g0186(.A1(G226), .A2(G1698), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n382), .A2(new_n385), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  AND2_X1   g0188(.A1(new_n388), .A2(KEYINPUT81), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n388), .A2(KEYINPUT81), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n336), .A2(G1698), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n382), .A2(new_n385), .A3(new_n386), .A4(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G33), .A2(G87), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NOR3_X1   g0194(.A1(new_n389), .A2(new_n390), .A3(new_n394), .ZN(new_n395));
  OAI211_X1 g0195(.A(G179), .B(new_n381), .C1(new_n395), .C2(new_n272), .ZN(new_n396));
  NOR3_X1   g0196(.A1(new_n264), .A2(KEYINPUT79), .A3(KEYINPUT3), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n384), .A2(G33), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT81), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n399), .A2(new_n400), .A3(new_n382), .A4(new_n387), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n388), .A2(KEYINPUT81), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n401), .A2(new_n402), .A3(new_n393), .A4(new_n392), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n380), .B1(new_n403), .B2(new_n338), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n396), .B1(new_n351), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT16), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT7), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n270), .B2(G20), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n384), .A2(G33), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n386), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n410), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n203), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  AND2_X1   g0212(.A1(G58), .A2(G68), .ZN(new_n413));
  NOR2_X1   g0213(.A1(G58), .A2(G68), .ZN(new_n414));
  OAI21_X1  g0214(.A(G20), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT80), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OAI211_X1 g0217(.A(KEYINPUT80), .B(G20), .C1(new_n413), .C2(new_n414), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n296), .A2(G159), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n406), .B1(new_n412), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n382), .A2(new_n385), .A3(new_n386), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n422), .A2(new_n407), .A3(new_n209), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n407), .B1(new_n422), .B2(new_n209), .ZN(new_n424));
  NOR3_X1   g0224(.A1(new_n423), .A2(new_n424), .A3(new_n203), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n417), .A2(KEYINPUT16), .A3(new_n418), .A4(new_n419), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n421), .B(new_n295), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n323), .B1(new_n208), .B2(G20), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n428), .A2(new_n308), .B1(new_n307), .B2(new_n323), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n405), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT18), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT18), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n405), .A2(new_n433), .A3(new_n430), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n403), .A2(new_n338), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n435), .A2(new_n315), .A3(new_n381), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(G200), .B2(new_n404), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT17), .ZN(new_n438));
  INV_X1    g0238(.A(new_n429), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n382), .A2(new_n385), .A3(new_n386), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT7), .B1(new_n440), .B2(G20), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n422), .A2(new_n407), .A3(new_n209), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n441), .A2(G68), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n426), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n327), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n439), .B1(new_n445), .B2(new_n421), .ZN(new_n446));
  AND3_X1   g0246(.A1(new_n437), .A2(new_n438), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n438), .B1(new_n437), .B2(new_n446), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n432), .B(new_n434), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  AND4_X1   g0250(.A1(new_n320), .A2(new_n377), .A3(new_n378), .A4(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT23), .ZN(new_n452));
  INV_X1    g0252(.A(G107), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n452), .A2(new_n453), .A3(G20), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT86), .ZN(new_n455));
  AOI21_X1  g0255(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n456));
  OAI22_X1  g0256(.A1(new_n454), .A2(new_n455), .B1(new_n456), .B2(G20), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n209), .A2(G87), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT22), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n461), .A2(new_n386), .A3(new_n382), .A4(new_n385), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n460), .B1(new_n410), .B2(new_n459), .ZN(new_n463));
  AOI22_X1  g0263(.A1(new_n454), .A2(new_n455), .B1(KEYINPUT23), .B2(G107), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n458), .A2(new_n462), .A3(new_n463), .A4(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT24), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n209), .A2(KEYINPUT23), .A3(G107), .ZN(new_n467));
  OAI22_X1  g0267(.A1(new_n467), .A2(KEYINPUT86), .B1(new_n452), .B2(new_n453), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(new_n457), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT24), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n469), .A2(new_n470), .A3(new_n462), .A4(new_n463), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n295), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT25), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n474), .B1(new_n304), .B2(G107), .ZN(new_n475));
  NOR3_X1   g0275(.A1(new_n304), .A2(new_n474), .A3(G107), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n208), .A2(G33), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n304), .A2(new_n478), .A3(new_n218), .A4(new_n294), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n475), .A2(new_n477), .B1(new_n480), .B2(G107), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n473), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n237), .A2(G1698), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(G250), .B2(G1698), .ZN(new_n484));
  INV_X1    g0284(.A(G294), .ZN(new_n485));
  OAI22_X1  g0285(.A1(new_n422), .A2(new_n484), .B1(new_n264), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n261), .A2(G1), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT5), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G41), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n260), .A2(KEYINPUT5), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n487), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n259), .A2(new_n491), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n338), .A2(new_n486), .B1(new_n492), .B2(G264), .ZN(new_n493));
  INV_X1    g0293(.A(G179), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n487), .A2(new_n490), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n495), .A2(new_n259), .A3(G274), .A4(new_n489), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n493), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n486), .A2(new_n338), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n492), .A2(G264), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n498), .A2(new_n499), .A3(new_n496), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n351), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n482), .A2(KEYINPUT87), .A3(new_n497), .A4(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT87), .ZN(new_n503));
  INV_X1    g0303(.A(new_n481), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n504), .B1(new_n472), .B2(new_n295), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n501), .A2(new_n497), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n503), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n500), .A2(G200), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n315), .B2(new_n500), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n482), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G283), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT4), .ZN(new_n514));
  INV_X1    g0314(.A(G244), .ZN(new_n515));
  NOR3_X1   g0315(.A1(new_n514), .A2(new_n515), .A3(G1698), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n270), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n514), .B1(new_n270), .B2(G250), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n513), .B(new_n517), .C1(new_n518), .C2(new_n334), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT4), .B1(new_n440), .B2(G244), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n338), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n259), .A2(new_n491), .A3(G257), .ZN(new_n522));
  XNOR2_X1  g0322(.A(new_n522), .B(KEYINPUT83), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n521), .A2(new_n523), .A3(new_n496), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(G200), .ZN(new_n525));
  XNOR2_X1  g0325(.A(KEYINPUT82), .B(KEYINPUT6), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n265), .B2(G107), .ZN(new_n527));
  XNOR2_X1  g0327(.A(G97), .B(G107), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n527), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  OAI22_X1  g0329(.A1(new_n529), .A2(new_n209), .B1(new_n300), .B2(new_n297), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n453), .B1(new_n408), .B2(new_n411), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n295), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n304), .A2(G97), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n533), .B1(new_n480), .B2(G97), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n521), .A2(new_n523), .A3(G190), .A4(new_n496), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n525), .A2(new_n532), .A3(new_n534), .A4(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n524), .A2(new_n351), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n532), .A2(new_n534), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n521), .A2(new_n523), .A3(new_n494), .A4(new_n496), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(G116), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n307), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n479), .B2(new_n542), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n294), .A2(new_n218), .B1(G20), .B2(new_n542), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n513), .B(new_n209), .C1(G33), .C2(new_n265), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(KEYINPUT20), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n545), .A2(new_n546), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT20), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n544), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n410), .A2(G303), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n237), .A2(new_n334), .ZN(new_n554));
  INV_X1    g0354(.A(G264), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G1698), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n553), .B1(new_n422), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n338), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n259), .A2(new_n491), .A3(G270), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n559), .A2(new_n496), .A3(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n552), .A2(new_n561), .A3(KEYINPUT21), .A4(G169), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n399), .A2(new_n382), .A3(new_n556), .A4(new_n554), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n272), .B1(new_n563), .B2(new_n553), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n496), .A2(new_n560), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n566), .A2(new_n552), .A3(G179), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT21), .ZN(new_n569));
  OAI21_X1  g0369(.A(G169), .B1(new_n564), .B2(new_n565), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n569), .B1(new_n570), .B2(new_n551), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n561), .A2(G200), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n572), .B(new_n551), .C1(new_n315), .C2(new_n561), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n568), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n515), .A2(G1698), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(G238), .B2(G1698), .ZN(new_n576));
  OAI22_X1  g0376(.A1(new_n422), .A2(new_n576), .B1(new_n264), .B2(new_n542), .ZN(new_n577));
  OR3_X1    g0377(.A1(new_n261), .A2(G1), .A3(G274), .ZN(new_n578));
  INV_X1    g0378(.A(G250), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(new_n261), .B2(G1), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n577), .A2(new_n338), .B1(new_n259), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(G190), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT85), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n582), .A2(KEYINPUT85), .A3(G190), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n577), .A2(new_n338), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n581), .A2(new_n259), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(G200), .ZN(new_n590));
  INV_X1    g0390(.A(new_n361), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n591), .A2(new_n304), .ZN(new_n592));
  INV_X1    g0392(.A(G87), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n479), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n593), .A2(new_n265), .A3(new_n453), .ZN(new_n595));
  OAI211_X1 g0395(.A(KEYINPUT19), .B(new_n595), .C1(new_n266), .C2(G20), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT19), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(new_n299), .B2(new_n265), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n209), .A2(G68), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n596), .B(new_n598), .C1(new_n422), .C2(new_n599), .ZN(new_n600));
  AOI211_X1 g0400(.A(new_n592), .B(new_n594), .C1(new_n600), .C2(new_n295), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n585), .A2(new_n586), .A3(new_n590), .A4(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n589), .A2(new_n351), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n592), .B1(new_n600), .B2(new_n295), .ZN(new_n604));
  OR2_X1    g0404(.A1(new_n361), .A2(KEYINPUT84), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n361), .A2(KEYINPUT84), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(new_n480), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n582), .A2(new_n494), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n603), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n602), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n574), .A2(new_n611), .ZN(new_n612));
  AND4_X1   g0412(.A1(new_n451), .A2(new_n512), .A3(new_n541), .A4(new_n612), .ZN(G372));
  AND3_X1   g0413(.A1(new_n537), .A2(new_n539), .A3(new_n538), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT26), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n590), .A2(new_n583), .A3(new_n601), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n614), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(KEYINPUT26), .B1(new_n611), .B2(new_n540), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n618), .A2(new_n619), .A3(new_n610), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n505), .A2(new_n506), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n571), .A2(new_n567), .A3(new_n562), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT88), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n610), .A2(new_n616), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n511), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n571), .A2(new_n567), .A3(new_n562), .ZN(new_n628));
  OAI21_X1  g0428(.A(KEYINPUT88), .B1(new_n628), .B2(new_n621), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n625), .A2(new_n541), .A3(new_n627), .A4(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n620), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n451), .A2(new_n631), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n319), .A2(new_n369), .ZN(new_n633));
  AOI21_X1  g0433(.A(G200), .B1(new_n435), .B2(new_n381), .ZN(new_n634));
  AOI211_X1 g0434(.A(G190), .B(new_n380), .C1(new_n403), .C2(new_n338), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n427), .B(new_n429), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT17), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n437), .A2(new_n438), .A3(new_n446), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n633), .A2(new_n312), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n405), .A2(new_n433), .A3(new_n430), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n433), .B1(new_n405), .B2(new_n430), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n350), .B1(new_n639), .B2(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n644), .A2(new_n353), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n632), .A2(new_n645), .ZN(G369));
  INV_X1    g0446(.A(KEYINPUT89), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n648), .A2(KEYINPUT27), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(KEYINPUT27), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n649), .A2(G213), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(G343), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n551), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n568), .A2(new_n571), .A3(new_n573), .A4(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n628), .A2(new_n653), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n647), .B1(new_n657), .B2(G330), .ZN(new_n658));
  INV_X1    g0458(.A(G330), .ZN(new_n659));
  AOI211_X1 g0459(.A(KEYINPUT89), .B(new_n659), .C1(new_n655), .C2(new_n656), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n505), .B(new_n509), .C1(new_n315), .C2(new_n500), .ZN(new_n662));
  INV_X1    g0462(.A(new_n652), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n482), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n502), .A2(new_n662), .A3(new_n507), .A4(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n621), .A2(new_n663), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT90), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n665), .A2(KEYINPUT90), .A3(new_n666), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n661), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n622), .A2(new_n663), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n669), .A2(new_n670), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n628), .A2(new_n652), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n673), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n672), .A2(new_n677), .ZN(G399));
  OR3_X1    g0478(.A1(new_n212), .A2(KEYINPUT91), .A3(G41), .ZN(new_n679));
  OAI21_X1  g0479(.A(KEYINPUT91), .B1(new_n212), .B2(G41), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n595), .A2(G116), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G1), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n216), .B2(new_n681), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT28), .ZN(new_n685));
  INV_X1    g0485(.A(new_n524), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n561), .A2(new_n494), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n493), .A2(new_n582), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n686), .A2(KEYINPUT30), .A3(new_n687), .A4(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT30), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n566), .A2(G179), .A3(new_n493), .A4(new_n582), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n690), .B1(new_n691), .B2(new_n524), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n566), .A2(G179), .A3(new_n582), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n693), .A2(new_n500), .A3(new_n524), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n689), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(KEYINPUT31), .B1(new_n695), .B2(new_n663), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT92), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n695), .A2(KEYINPUT31), .A3(new_n663), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n512), .A2(new_n541), .A3(new_n612), .A4(new_n652), .ZN(new_n700));
  INV_X1    g0500(.A(new_n698), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT92), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n699), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G330), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n502), .A2(new_n623), .A3(new_n507), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n662), .A2(new_n536), .A3(new_n540), .A4(new_n617), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n614), .A2(new_n615), .A3(new_n610), .A4(new_n602), .ZN(new_n709));
  OAI21_X1  g0509(.A(KEYINPUT26), .B1(new_n540), .B2(new_n626), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(new_n610), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n652), .B1(new_n708), .B2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT93), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n610), .ZN(new_n715));
  AOI22_X1  g0515(.A1(new_n524), .A2(new_n351), .B1(new_n532), .B2(new_n534), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n617), .A2(new_n539), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n715), .B1(new_n717), .B2(KEYINPUT26), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n718), .B(new_n709), .C1(new_n706), .C2(new_n707), .ZN(new_n719));
  AOI21_X1  g0519(.A(KEYINPUT93), .B1(new_n719), .B2(new_n652), .ZN(new_n720));
  OAI21_X1  g0520(.A(KEYINPUT29), .B1(new_n714), .B2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n663), .B1(new_n620), .B2(new_n630), .ZN(new_n722));
  OR2_X1    g0522(.A1(new_n722), .A2(KEYINPUT29), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n705), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n685), .B1(new_n724), .B2(G1), .ZN(G364));
  INV_X1    g0525(.A(new_n681), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n209), .A2(G13), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT94), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n208), .B1(new_n728), .B2(G45), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OAI221_X1 g0530(.A(new_n661), .B1(G330), .B2(new_n657), .C1(new_n726), .C2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n726), .A2(new_n730), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n212), .A2(new_n410), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n733), .B(KEYINPUT95), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G355), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n735), .B1(G116), .B2(new_n213), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n249), .A2(G45), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n440), .A2(new_n212), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n739), .B1(new_n261), .B2(new_n217), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n736), .B1(new_n737), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G13), .A2(G33), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G20), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n218), .B1(G20), .B2(new_n351), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n732), .B1(new_n741), .B2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n745), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n209), .A2(new_n494), .ZN(new_n750));
  INV_X1    g0550(.A(G200), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n750), .A2(G190), .A3(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n209), .A2(G179), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G190), .A2(G200), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(G159), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT32), .ZN(new_n758));
  OAI221_X1 g0558(.A(new_n270), .B1(new_n752), .B2(new_n202), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n750), .A2(G200), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n315), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n760), .B1(new_n763), .B2(new_n201), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n750), .A2(new_n754), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(KEYINPUT96), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n765), .A2(KEYINPUT96), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI211_X1 g0570(.A(new_n759), .B(new_n764), .C1(G77), .C2(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n753), .A2(G190), .A3(G200), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT97), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n772), .A2(new_n773), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n593), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n753), .A2(new_n315), .A3(G200), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n778), .B(KEYINPUT98), .Z(new_n779));
  AOI21_X1  g0579(.A(new_n777), .B1(G107), .B2(new_n779), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n315), .A2(G179), .A3(G200), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n209), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n761), .A2(G190), .ZN(new_n784));
  AOI22_X1  g0584(.A1(G97), .A2(new_n783), .B1(new_n784), .B2(G68), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT99), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n771), .A2(new_n780), .A3(new_n786), .ZN(new_n787));
  XNOR2_X1  g0587(.A(KEYINPUT33), .B(G317), .ZN(new_n788));
  INV_X1    g0588(.A(new_n752), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n784), .A2(new_n788), .B1(new_n789), .B2(G322), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(KEYINPUT100), .Z(new_n791));
  NAND2_X1  g0591(.A1(new_n762), .A2(G326), .ZN(new_n792));
  INV_X1    g0592(.A(new_n755), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n270), .B1(new_n793), .B2(G329), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n792), .B(new_n794), .C1(new_n485), .C2(new_n782), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n795), .B1(G311), .B2(new_n770), .ZN(new_n796));
  INV_X1    g0596(.A(new_n776), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n797), .A2(G303), .B1(new_n779), .B2(G283), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n791), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n749), .B1(new_n787), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n748), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n744), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n801), .B1(new_n657), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n731), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(G396));
  NAND2_X1  g0605(.A1(new_n369), .A2(KEYINPUT105), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT105), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n359), .A2(new_n367), .A3(new_n807), .A4(new_n368), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n809), .A2(new_n371), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n722), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n367), .A2(new_n663), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n806), .A2(new_n371), .A3(new_n812), .A4(new_n808), .ZN(new_n813));
  OR2_X1    g0613(.A1(new_n369), .A2(new_n652), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n811), .B1(new_n722), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n732), .B1(new_n816), .B2(new_n704), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n704), .B2(new_n816), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n745), .A2(new_n742), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT101), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n732), .B1(G77), .B2(new_n820), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT102), .ZN(new_n822));
  INV_X1    g0622(.A(new_n779), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n823), .A2(new_n593), .B1(new_n453), .B2(new_n776), .ZN(new_n824));
  AOI22_X1  g0624(.A1(G97), .A2(new_n783), .B1(new_n762), .B2(G303), .ZN(new_n825));
  INV_X1    g0625(.A(G283), .ZN(new_n826));
  INV_X1    g0626(.A(new_n784), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n769), .A2(new_n542), .ZN(new_n829));
  INV_X1    g0629(.A(G311), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n410), .B1(new_n755), .B2(new_n830), .C1(new_n752), .C2(new_n485), .ZN(new_n831));
  NOR4_X1   g0631(.A1(new_n824), .A2(new_n828), .A3(new_n829), .A4(new_n831), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(KEYINPUT103), .ZN(new_n833));
  INV_X1    g0633(.A(G132), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n440), .B1(new_n834), .B2(new_n755), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n823), .A2(new_n203), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n835), .B(new_n836), .C1(G58), .C2(new_n783), .ZN(new_n837));
  AOI22_X1  g0637(.A1(G150), .A2(new_n784), .B1(new_n789), .B2(G143), .ZN(new_n838));
  INV_X1    g0638(.A(G137), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n838), .B1(new_n839), .B2(new_n763), .C1(new_n769), .C2(new_n756), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT34), .ZN(new_n841));
  OR2_X1    g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n840), .A2(new_n841), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n797), .A2(G50), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n837), .A2(new_n842), .A3(new_n843), .A4(new_n844), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n833), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n822), .B1(new_n846), .B2(new_n749), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n847), .B(KEYINPUT104), .Z(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n743), .B2(new_n815), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n818), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(G384));
  INV_X1    g0651(.A(KEYINPUT35), .ZN(new_n852));
  OAI211_X1 g0652(.A(G116), .B(new_n219), .C1(new_n529), .C2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(new_n852), .B2(new_n529), .ZN(new_n854));
  XOR2_X1   g0654(.A(KEYINPUT106), .B(KEYINPUT36), .Z(new_n855));
  XNOR2_X1  g0655(.A(new_n854), .B(new_n855), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n217), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n201), .A2(G68), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n208), .B(G13), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT38), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n430), .A2(new_n651), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n431), .A2(new_n636), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(KEYINPUT37), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT37), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n431), .A2(new_n636), .A3(new_n862), .A4(new_n865), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n637), .A2(new_n638), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n862), .B1(new_n642), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n861), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n295), .B1(new_n425), .B2(new_n426), .ZN(new_n871));
  INV_X1    g0671(.A(new_n420), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT16), .B1(new_n443), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n429), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n651), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n405), .A2(new_n874), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n877), .A2(new_n875), .A3(new_n636), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT37), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n449), .A2(new_n876), .B1(new_n879), .B2(new_n866), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n870), .A2(KEYINPUT109), .B1(KEYINPUT38), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT39), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT109), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n883), .B(new_n861), .C1(new_n867), .C2(new_n869), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n881), .A2(KEYINPUT110), .A3(new_n882), .A4(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n862), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n449), .A2(new_n886), .B1(new_n864), .B2(new_n866), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT109), .B1(new_n887), .B2(KEYINPUT38), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n880), .A2(KEYINPUT38), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n888), .A2(new_n884), .A3(new_n882), .A4(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT110), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n449), .A2(new_n876), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n879), .A2(new_n866), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n861), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n889), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(KEYINPUT39), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n885), .A2(new_n892), .A3(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT108), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n313), .B2(new_n652), .ZN(new_n901));
  NOR3_X1   g0701(.A1(new_n312), .A2(KEYINPUT108), .A3(new_n663), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n899), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n642), .A2(new_n651), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT107), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n893), .A2(KEYINPUT38), .A3(new_n894), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT38), .B1(new_n893), .B2(new_n894), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n896), .A2(KEYINPUT107), .A3(new_n889), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n311), .A2(new_n663), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n312), .A2(new_n318), .A3(new_n913), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n311), .B(new_n663), .C1(new_n293), .C2(new_n319), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n809), .A2(new_n663), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(new_n722), .B2(new_n810), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n906), .B1(new_n912), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n905), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n721), .A2(new_n451), .A3(new_n723), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n645), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n922), .B(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n815), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n701), .A2(new_n696), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n926), .B1(new_n927), .B2(new_n700), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n928), .A2(new_n916), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n888), .A2(new_n884), .A3(new_n889), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n929), .A2(KEYINPUT40), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n928), .A2(new_n916), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n910), .B2(new_n911), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n931), .B1(new_n933), .B2(KEYINPUT40), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n927), .A2(new_n700), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n451), .A2(new_n935), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n934), .A2(new_n936), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n937), .A2(G330), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n925), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n208), .B2(new_n728), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n925), .A2(new_n939), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n860), .B1(new_n941), .B2(new_n942), .ZN(G367));
  NOR2_X1   g0743(.A1(new_n601), .A2(new_n652), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n610), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n617), .B2(new_n944), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT111), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT43), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n675), .B1(new_n669), .B2(new_n670), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n538), .A2(new_n663), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n541), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n614), .A2(new_n663), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n950), .A2(new_n954), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n955), .A2(KEYINPUT42), .ZN(new_n956));
  INV_X1    g0756(.A(new_n508), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n540), .B1(new_n952), .B2(new_n957), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n955), .A2(KEYINPUT42), .B1(new_n652), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n949), .B1(new_n956), .B2(new_n959), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n947), .A2(new_n948), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n956), .A2(new_n959), .A3(new_n948), .A4(new_n947), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n954), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n672), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n963), .A2(new_n967), .A3(new_n964), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n681), .B(KEYINPUT112), .Z(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT41), .Z(new_n974));
  INV_X1    g0774(.A(new_n661), .ZN(new_n975));
  AND3_X1   g0775(.A1(new_n665), .A2(KEYINPUT90), .A3(new_n666), .ZN(new_n976));
  AOI21_X1  g0776(.A(KEYINPUT90), .B1(new_n665), .B2(new_n666), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n676), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n669), .A2(new_n670), .A3(new_n675), .ZN(new_n979));
  AND3_X1   g0779(.A1(new_n975), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n975), .B1(new_n978), .B2(new_n979), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n724), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT114), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n672), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n966), .B1(new_n950), .B2(new_n673), .ZN(new_n987));
  XNOR2_X1  g0787(.A(KEYINPUT113), .B(KEYINPUT44), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n966), .B(new_n988), .C1(new_n950), .C2(new_n673), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n671), .A2(KEYINPUT114), .ZN(new_n992));
  AND3_X1   g0792(.A1(new_n990), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n677), .A2(KEYINPUT45), .A3(new_n954), .ZN(new_n994));
  INV_X1    g0794(.A(new_n673), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n978), .A2(new_n995), .A3(new_n954), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT45), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n994), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n986), .B1(new_n993), .B2(new_n999), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n987), .A2(new_n989), .B1(new_n671), .B2(KEYINPUT114), .ZN(new_n1001));
  AND4_X1   g0801(.A1(new_n986), .A2(new_n999), .A3(new_n1001), .A4(new_n991), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n984), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n974), .B1(new_n1003), .B2(new_n724), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n972), .B1(new_n1004), .B2(new_n730), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n238), .A2(new_n738), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1006), .B(new_n746), .C1(new_n213), .C2(new_n361), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n410), .B1(new_n793), .B2(G137), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1008), .B1(new_n300), .B2(new_n778), .C1(new_n827), .C2(new_n756), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(G50), .B2(new_n770), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n202), .B2(new_n776), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(G143), .A2(new_n762), .B1(new_n789), .B2(G150), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n203), .B2(new_n782), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT115), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n776), .A2(new_n542), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT46), .ZN(new_n1016));
  INV_X1    g0816(.A(G317), .ZN(new_n1017));
  INV_X1    g0817(.A(G303), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n422), .B1(new_n755), .B2(new_n1017), .C1(new_n752), .C2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(new_n770), .B2(G283), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n778), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n783), .A2(G107), .B1(new_n1021), .B2(G97), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(G294), .A2(new_n784), .B1(new_n762), .B2(G311), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1020), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n1011), .A2(new_n1014), .B1(new_n1016), .B2(new_n1024), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT47), .Z(new_n1026));
  OAI211_X1 g0826(.A(new_n732), .B(new_n1007), .C1(new_n1026), .C2(new_n749), .ZN(new_n1027));
  AND2_X1   g0827(.A1(new_n947), .A2(new_n744), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1005), .A2(new_n1030), .ZN(G387));
  OR2_X1    g0831(.A1(new_n724), .A2(new_n982), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1032), .A2(new_n726), .A3(new_n983), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n982), .A2(new_n730), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n776), .A2(new_n300), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(G97), .B2(new_n779), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n756), .A2(new_n763), .B1(new_n827), .B2(new_n323), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(KEYINPUT116), .B(G150), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n752), .A2(new_n201), .B1(new_n755), .B2(new_n1038), .ZN(new_n1039));
  NOR3_X1   g0839(.A1(new_n1037), .A2(new_n422), .A3(new_n1039), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n605), .A2(new_n783), .A3(new_n606), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n770), .A2(G68), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1036), .A2(new_n1040), .A3(new_n1041), .A4(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n440), .B1(G326), .B2(new_n793), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n776), .A2(new_n485), .B1(new_n826), .B2(new_n782), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G311), .A2(new_n784), .B1(new_n789), .B2(G317), .ZN(new_n1046));
  INV_X1    g0846(.A(G322), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1046), .B1(new_n1047), .B2(new_n763), .C1(new_n769), .C2(new_n1018), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT48), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1045), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n1049), .B2(new_n1048), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT49), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1044), .B1(new_n542), .B2(new_n778), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  AND2_X1   g0853(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1043), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n745), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n739), .B1(new_n244), .B2(G45), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n682), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1057), .B1(new_n1058), .B2(new_n734), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n323), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n201), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT50), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n261), .B1(new_n203), .B2(new_n300), .ZN(new_n1063));
  NOR3_X1   g0863(.A1(new_n1062), .A2(new_n1058), .A3(new_n1063), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n1059), .A2(new_n1064), .B1(G107), .B2(new_n213), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n726), .B(new_n730), .C1(new_n1065), .C2(new_n746), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1056), .B(new_n1066), .C1(new_n674), .C2(new_n802), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n1034), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1033), .A2(new_n1068), .ZN(G393));
  INV_X1    g0869(.A(new_n986), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n999), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n990), .A2(new_n992), .A3(new_n991), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n999), .A2(new_n1001), .A3(new_n986), .A4(new_n991), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1073), .A2(new_n983), .A3(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1003), .A2(new_n726), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n966), .A2(new_n744), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n746), .B1(new_n265), .B2(new_n213), .C1(new_n739), .C2(new_n252), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n732), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n763), .A2(new_n1017), .B1(new_n830), .B2(new_n752), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT52), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n797), .A2(G283), .B1(new_n779), .B2(G107), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n770), .A2(G294), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n410), .B1(new_n755), .B2(new_n1047), .C1(new_n782), .C2(new_n542), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(G303), .B2(new_n784), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .A4(new_n1086), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n827), .A2(new_n201), .B1(new_n300), .B2(new_n782), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n422), .B(new_n1088), .C1(G143), .C2(new_n793), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n797), .A2(G68), .B1(new_n779), .B2(G87), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1089), .B(new_n1090), .C1(new_n323), .C2(new_n769), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(G150), .A2(new_n762), .B1(new_n789), .B2(G159), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT51), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1087), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1080), .B1(new_n1094), .B2(new_n745), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n1077), .A2(new_n730), .B1(new_n1078), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1076), .A2(new_n1096), .ZN(G390));
  AOI22_X1  g0897(.A1(new_n890), .A2(new_n891), .B1(KEYINPUT39), .B2(new_n897), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n903), .B1(new_n919), .B2(new_n917), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1098), .A2(new_n885), .A3(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n712), .A2(new_n713), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n719), .A2(KEYINPUT93), .A3(new_n652), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n926), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n916), .B1(new_n1103), .B2(new_n918), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n930), .A2(new_n903), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n705), .A2(new_n815), .A3(new_n916), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1100), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n932), .A2(new_n659), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n1100), .B2(new_n1106), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n1109), .A2(new_n729), .A3(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1098), .A2(new_n742), .A3(new_n885), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n732), .B1(new_n1060), .B2(new_n820), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n782), .A2(new_n300), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n410), .B1(new_n755), .B2(new_n485), .C1(new_n752), .C2(new_n542), .ZN(new_n1117));
  NOR4_X1   g0917(.A1(new_n836), .A2(new_n777), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(G107), .A2(new_n784), .B1(new_n762), .B2(G283), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n769), .B2(new_n265), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT118), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT119), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n776), .A2(new_n1038), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT53), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n762), .A2(G128), .B1(new_n1021), .B2(G50), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(G159), .A2(new_n783), .B1(new_n784), .B2(G137), .ZN(new_n1127));
  INV_X1    g0927(.A(G125), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n270), .B1(new_n755), .B2(new_n1128), .C1(new_n752), .C2(new_n834), .ZN(new_n1129));
  XOR2_X1   g0929(.A(KEYINPUT54), .B(G143), .Z(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT117), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1129), .B1(new_n770), .B2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .A4(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(KEYINPUT120), .B1(new_n1123), .B2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1134), .A2(new_n749), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1123), .A2(KEYINPUT120), .A3(new_n1133), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1115), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1113), .B1(new_n1114), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n659), .B1(new_n927), .B2(new_n700), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n451), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n923), .A2(new_n1140), .A3(new_n645), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n919), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n916), .B1(new_n705), .B2(new_n815), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1142), .B1(new_n1143), .B2(new_n1110), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1103), .A2(new_n918), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1139), .A2(new_n815), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n917), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1145), .A2(new_n1107), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1141), .B1(new_n1144), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1100), .A2(new_n1106), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n1110), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1153), .A2(new_n1149), .A3(new_n1108), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1151), .A2(new_n726), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1138), .A2(new_n1155), .ZN(G378));
  NAND2_X1  g0956(.A1(new_n350), .A2(new_n353), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1157), .B(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n328), .A2(new_n651), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1159), .B(new_n1160), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1161), .A2(KEYINPUT121), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  OAI211_X1 g0963(.A(G330), .B(new_n931), .C1(new_n933), .C2(KEYINPUT40), .ZN(new_n1164));
  AND3_X1   g0964(.A1(new_n905), .A2(new_n921), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1164), .B1(new_n905), .B2(new_n921), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1163), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1164), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n903), .B1(new_n1098), .B2(new_n885), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n921), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1168), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n905), .A2(new_n921), .A3(new_n1164), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1171), .A2(new_n1162), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1167), .A2(new_n1173), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1161), .A2(new_n743), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n732), .B1(G50), .B2(new_n820), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n422), .A2(new_n260), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n752), .A2(new_n453), .B1(new_n755), .B2(new_n826), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1177), .B(new_n1178), .C1(G68), .C2(new_n783), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n605), .A2(new_n606), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1179), .B1(new_n1180), .B2(new_n769), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n778), .A2(new_n202), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(G97), .B2(new_n784), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n542), .B2(new_n763), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n1181), .A2(new_n1035), .A3(new_n1184), .ZN(new_n1185));
  OR2_X1    g0985(.A1(new_n1185), .A2(KEYINPUT58), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n770), .A2(G137), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n797), .A2(new_n1131), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(G125), .A2(new_n762), .B1(new_n789), .B2(G128), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(G150), .A2(new_n783), .B1(new_n784), .B2(G132), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n1191), .A2(KEYINPUT59), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(KEYINPUT59), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1021), .A2(G159), .ZN(new_n1194));
  AOI211_X1 g0994(.A(G33), .B(G41), .C1(new_n793), .C2(G124), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1185), .A2(KEYINPUT58), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1177), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1186), .A2(new_n1196), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1176), .B1(new_n1199), .B2(new_n745), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n1174), .A2(new_n730), .B1(new_n1175), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1141), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1167), .A2(new_n1173), .B1(new_n1202), .B2(new_n1154), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n726), .B1(new_n1203), .B2(KEYINPUT57), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1154), .A2(new_n1202), .ZN(new_n1205));
  AND3_X1   g1005(.A1(new_n1174), .A2(KEYINPUT57), .A3(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1201), .B1(new_n1204), .B2(new_n1206), .ZN(G375));
  INV_X1    g1007(.A(KEYINPUT123), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n1144), .A2(new_n1148), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1208), .B1(new_n1209), .B2(new_n729), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1144), .A2(new_n1148), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1211), .A2(KEYINPUT123), .A3(new_n730), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n732), .B1(G68), .B2(new_n820), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1041), .B1(new_n826), .B2(new_n752), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT124), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n410), .B1(new_n755), .B2(new_n1018), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(G116), .B2(new_n784), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n485), .B2(new_n763), .C1(new_n769), .C2(new_n453), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n823), .A2(new_n300), .B1(new_n776), .B2(new_n265), .ZN(new_n1219));
  NOR3_X1   g1019(.A1(new_n1215), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1220), .B(KEYINPUT125), .ZN(new_n1221));
  INV_X1    g1021(.A(G128), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n440), .B1(new_n1222), .B2(new_n755), .C1(new_n839), .C2(new_n752), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(new_n770), .B2(G150), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1131), .A2(new_n784), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n797), .A2(G159), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n782), .A2(new_n201), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n1182), .B(new_n1227), .C1(G132), .C2(new_n762), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .A4(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1221), .A2(new_n1229), .ZN(new_n1230));
  OR2_X1    g1030(.A1(new_n1230), .A2(KEYINPUT126), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n749), .B1(new_n1230), .B2(KEYINPUT126), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1213), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(new_n743), .B2(new_n916), .ZN(new_n1234));
  AND3_X1   g1034(.A1(new_n1210), .A2(new_n1212), .A3(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1209), .A2(new_n1141), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n974), .B(KEYINPUT122), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1236), .A2(new_n1150), .A3(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1235), .A2(new_n1238), .ZN(G381));
  AND2_X1   g1039(.A1(new_n1076), .A2(new_n1096), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1005), .A2(new_n1240), .A3(new_n1030), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1033), .A2(new_n804), .A3(new_n1068), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1235), .A2(new_n850), .A3(new_n1238), .A4(new_n1243), .ZN(new_n1244));
  OR4_X1    g1044(.A1(G378), .A2(G375), .A3(new_n1241), .A4(new_n1244), .ZN(G407));
  INV_X1    g1045(.A(G378), .ZN(new_n1246));
  INV_X1    g1046(.A(G213), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1247), .A2(G343), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1246), .A2(new_n1248), .ZN(new_n1249));
  OAI211_X1 g1049(.A(G407), .B(G213), .C1(G375), .C2(new_n1249), .ZN(G409));
  AOI21_X1  g1050(.A(new_n804), .B1(new_n1033), .B2(new_n1068), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1243), .A2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1240), .B1(new_n1005), .B2(new_n1030), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n974), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n983), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n724), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1254), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n971), .B1(new_n1257), .B2(new_n729), .ZN(new_n1258));
  NOR3_X1   g1058(.A1(new_n1258), .A2(G390), .A3(new_n1029), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1252), .B1(new_n1253), .B2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT61), .ZN(new_n1261));
  OAI21_X1  g1061(.A(G390), .B1(new_n1258), .B2(new_n1029), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1252), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1241), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1260), .A2(new_n1261), .A3(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT127), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1265), .B(new_n1266), .ZN(new_n1267));
  OAI211_X1 g1067(.A(G378), .B(new_n1201), .C1(new_n1204), .C2(new_n1206), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1174), .A2(new_n1205), .A3(new_n1237), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1201), .A2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1246), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1248), .B1(new_n1268), .B2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT60), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1236), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1209), .A2(KEYINPUT60), .A3(new_n1141), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1274), .A2(new_n726), .A3(new_n1150), .A4(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(new_n1235), .A3(G384), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(G384), .B1(new_n1276), .B2(new_n1235), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1272), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT63), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  OAI211_X1 g1083(.A(G2897), .B(new_n1248), .C1(new_n1278), .C2(new_n1279), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1279), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1248), .A2(G2897), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1285), .A2(new_n1277), .A3(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1284), .A2(new_n1287), .ZN(new_n1288));
  OR2_X1    g1088(.A1(new_n1272), .A2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1272), .A2(KEYINPUT63), .A3(new_n1280), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1267), .A2(new_n1283), .A3(new_n1289), .A4(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT62), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1272), .A2(new_n1292), .A3(new_n1280), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1261), .B1(new_n1272), .B2(new_n1288), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1292), .B1(new_n1272), .B2(new_n1280), .ZN(new_n1295));
  NOR3_X1   g1095(.A1(new_n1293), .A2(new_n1294), .A3(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1260), .A2(new_n1264), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1291), .B1(new_n1296), .B2(new_n1298), .ZN(G405));
  NAND2_X1  g1099(.A1(G375), .A2(new_n1246), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1268), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1298), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1297), .A2(new_n1300), .A3(new_n1268), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1280), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(new_n1304), .B(new_n1305), .ZN(G402));
endmodule


