

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X2 U322 ( .A(n409), .B(n408), .ZN(n515) );
  XNOR2_X1 U323 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U324 ( .A(n410), .B(n293), .ZN(n411) );
  XOR2_X1 U325 ( .A(n436), .B(KEYINPUT28), .Z(n519) );
  XOR2_X1 U326 ( .A(n398), .B(n397), .Z(n525) );
  XOR2_X1 U327 ( .A(n301), .B(n300), .Z(n290) );
  XOR2_X1 U328 ( .A(n405), .B(n394), .Z(n291) );
  XOR2_X1 U329 ( .A(n416), .B(n415), .Z(n292) );
  AND2_X1 U330 ( .A1(G228GAT), .A2(G233GAT), .ZN(n293) );
  OR2_X1 U331 ( .A1(n454), .A2(n453), .ZN(n455) );
  XNOR2_X1 U332 ( .A(n465), .B(KEYINPUT121), .ZN(n466) );
  XNOR2_X1 U333 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U334 ( .A(KEYINPUT113), .B(KEYINPUT48), .ZN(n462) );
  XNOR2_X1 U335 ( .A(n417), .B(n292), .ZN(n418) );
  XNOR2_X1 U336 ( .A(n302), .B(n290), .ZN(n303) );
  XNOR2_X1 U337 ( .A(n463), .B(n462), .ZN(n524) );
  XNOR2_X1 U338 ( .A(n419), .B(n418), .ZN(n424) );
  XNOR2_X1 U339 ( .A(n304), .B(n303), .ZN(n305) );
  INV_X1 U340 ( .A(G29GAT), .ZN(n447) );
  XNOR2_X1 U341 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U342 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U343 ( .A(n477), .B(n476), .ZN(G1351GAT) );
  XNOR2_X1 U344 ( .A(n450), .B(n449), .ZN(G1328GAT) );
  XNOR2_X1 U345 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n294) );
  XNOR2_X1 U346 ( .A(n294), .B(KEYINPUT7), .ZN(n328) );
  XOR2_X1 U347 ( .A(G36GAT), .B(G8GAT), .Z(n405) );
  XNOR2_X1 U348 ( .A(G43GAT), .B(G15GAT), .ZN(n295) );
  XNOR2_X1 U349 ( .A(n295), .B(G113GAT), .ZN(n394) );
  XNOR2_X1 U350 ( .A(G169GAT), .B(G197GAT), .ZN(n296) );
  XNOR2_X1 U351 ( .A(n291), .B(n296), .ZN(n304) );
  XOR2_X1 U352 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n298) );
  XNOR2_X1 U353 ( .A(KEYINPUT71), .B(KEYINPUT70), .ZN(n297) );
  XNOR2_X1 U354 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U355 ( .A(n299), .B(KEYINPUT72), .ZN(n302) );
  XOR2_X1 U356 ( .A(KEYINPUT69), .B(G1GAT), .Z(n301) );
  NAND2_X1 U357 ( .A1(G229GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U358 ( .A(n328), .B(n305), .ZN(n307) );
  XOR2_X1 U359 ( .A(G50GAT), .B(G22GAT), .Z(n306) );
  XOR2_X1 U360 ( .A(G141GAT), .B(n306), .Z(n420) );
  XOR2_X1 U361 ( .A(n307), .B(n420), .Z(n568) );
  XNOR2_X1 U362 ( .A(KEYINPUT73), .B(n568), .ZN(n555) );
  XNOR2_X1 U363 ( .A(G99GAT), .B(G71GAT), .ZN(n308) );
  XNOR2_X1 U364 ( .A(n308), .B(G120GAT), .ZN(n389) );
  XNOR2_X1 U365 ( .A(G204GAT), .B(G92GAT), .ZN(n309) );
  XNOR2_X1 U366 ( .A(n309), .B(G64GAT), .ZN(n401) );
  XOR2_X1 U367 ( .A(n389), .B(n401), .Z(n321) );
  XOR2_X1 U368 ( .A(G85GAT), .B(G57GAT), .Z(n371) );
  XOR2_X1 U369 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n311) );
  XNOR2_X1 U370 ( .A(G176GAT), .B(KEYINPUT75), .ZN(n310) );
  XNOR2_X1 U371 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U372 ( .A(n371), .B(n312), .Z(n314) );
  NAND2_X1 U373 ( .A1(G230GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U374 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U375 ( .A(n315), .B(KEYINPUT13), .Z(n319) );
  XOR2_X1 U376 ( .A(G78GAT), .B(G148GAT), .Z(n317) );
  XNOR2_X1 U377 ( .A(G106GAT), .B(KEYINPUT74), .ZN(n316) );
  XNOR2_X1 U378 ( .A(n317), .B(n316), .ZN(n414) );
  XNOR2_X1 U379 ( .A(n414), .B(KEYINPUT31), .ZN(n318) );
  XNOR2_X1 U380 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U381 ( .A(n321), .B(n320), .ZN(n572) );
  NAND2_X1 U382 ( .A1(n555), .A2(n572), .ZN(n482) );
  XOR2_X1 U383 ( .A(KEYINPUT76), .B(G162GAT), .Z(n410) );
  XOR2_X1 U384 ( .A(KEYINPUT78), .B(KEYINPUT10), .Z(n323) );
  XNOR2_X1 U385 ( .A(G218GAT), .B(G85GAT), .ZN(n322) );
  XNOR2_X1 U386 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U387 ( .A(n410), .B(n324), .Z(n326) );
  NAND2_X1 U388 ( .A1(G232GAT), .A2(G233GAT), .ZN(n325) );
  XNOR2_X1 U389 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U390 ( .A(n327), .B(G43GAT), .ZN(n330) );
  XOR2_X1 U391 ( .A(n328), .B(G50GAT), .Z(n329) );
  XNOR2_X1 U392 ( .A(n330), .B(n329), .ZN(n334) );
  XOR2_X1 U393 ( .A(KEYINPUT66), .B(KEYINPUT11), .Z(n332) );
  XNOR2_X1 U394 ( .A(G190GAT), .B(KEYINPUT77), .ZN(n331) );
  XNOR2_X1 U395 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U396 ( .A(n334), .B(n333), .ZN(n342) );
  XOR2_X1 U397 ( .A(KEYINPUT64), .B(G92GAT), .Z(n336) );
  XNOR2_X1 U398 ( .A(G99GAT), .B(G106GAT), .ZN(n335) );
  XNOR2_X1 U399 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U400 ( .A(KEYINPUT67), .B(KEYINPUT9), .Z(n338) );
  XNOR2_X1 U401 ( .A(G36GAT), .B(G134GAT), .ZN(n337) );
  XNOR2_X1 U402 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U403 ( .A(n340), .B(n339), .Z(n341) );
  XNOR2_X1 U404 ( .A(n342), .B(n341), .ZN(n536) );
  INV_X1 U405 ( .A(n536), .ZN(n553) );
  XOR2_X1 U406 ( .A(KEYINPUT36), .B(n553), .Z(n581) );
  XOR2_X1 U407 ( .A(KEYINPUT13), .B(G64GAT), .Z(n344) );
  XNOR2_X1 U408 ( .A(G1GAT), .B(G57GAT), .ZN(n343) );
  XNOR2_X1 U409 ( .A(n344), .B(n343), .ZN(n348) );
  XOR2_X1 U410 ( .A(KEYINPUT80), .B(KEYINPUT12), .Z(n346) );
  XNOR2_X1 U411 ( .A(G8GAT), .B(KEYINPUT81), .ZN(n345) );
  XNOR2_X1 U412 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U413 ( .A(n348), .B(n347), .ZN(n361) );
  XOR2_X1 U414 ( .A(G155GAT), .B(G78GAT), .Z(n350) );
  XNOR2_X1 U415 ( .A(G22GAT), .B(G211GAT), .ZN(n349) );
  XNOR2_X1 U416 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U417 ( .A(G127GAT), .B(G71GAT), .Z(n352) );
  XNOR2_X1 U418 ( .A(G15GAT), .B(G183GAT), .ZN(n351) );
  XNOR2_X1 U419 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U420 ( .A(n354), .B(n353), .Z(n359) );
  XOR2_X1 U421 ( .A(KEYINPUT79), .B(KEYINPUT15), .Z(n356) );
  NAND2_X1 U422 ( .A1(G231GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U423 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U424 ( .A(KEYINPUT14), .B(n357), .ZN(n358) );
  XNOR2_X1 U425 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U426 ( .A(n361), .B(n360), .Z(n563) );
  XOR2_X1 U427 ( .A(KEYINPUT6), .B(KEYINPUT90), .Z(n363) );
  XNOR2_X1 U428 ( .A(KEYINPUT91), .B(KEYINPUT1), .ZN(n362) );
  XNOR2_X1 U429 ( .A(n363), .B(n362), .ZN(n382) );
  XOR2_X1 U430 ( .A(KEYINPUT89), .B(G120GAT), .Z(n365) );
  XNOR2_X1 U431 ( .A(G1GAT), .B(G113GAT), .ZN(n364) );
  XNOR2_X1 U432 ( .A(n365), .B(n364), .ZN(n369) );
  XOR2_X1 U433 ( .A(G162GAT), .B(G148GAT), .Z(n367) );
  XNOR2_X1 U434 ( .A(G29GAT), .B(G141GAT), .ZN(n366) );
  XNOR2_X1 U435 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U436 ( .A(n369), .B(n368), .ZN(n380) );
  XNOR2_X1 U437 ( .A(G134GAT), .B(G127GAT), .ZN(n370) );
  XNOR2_X1 U438 ( .A(n370), .B(KEYINPUT0), .ZN(n393) );
  XOR2_X1 U439 ( .A(n371), .B(n393), .Z(n373) );
  NAND2_X1 U440 ( .A1(G225GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U441 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U442 ( .A(n374), .B(KEYINPUT4), .Z(n378) );
  XOR2_X1 U443 ( .A(G155GAT), .B(KEYINPUT3), .Z(n376) );
  XNOR2_X1 U444 ( .A(KEYINPUT87), .B(KEYINPUT2), .ZN(n375) );
  XNOR2_X1 U445 ( .A(n376), .B(n375), .ZN(n412) );
  XNOR2_X1 U446 ( .A(n412), .B(KEYINPUT5), .ZN(n377) );
  XNOR2_X1 U447 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U448 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U449 ( .A(n382), .B(n381), .ZN(n511) );
  XOR2_X1 U450 ( .A(G176GAT), .B(G183GAT), .Z(n384) );
  XNOR2_X1 U451 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n383) );
  XNOR2_X1 U452 ( .A(n384), .B(n383), .ZN(n388) );
  XOR2_X1 U453 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n386) );
  XNOR2_X1 U454 ( .A(G190GAT), .B(KEYINPUT83), .ZN(n385) );
  XNOR2_X1 U455 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U456 ( .A(n388), .B(n387), .Z(n409) );
  XNOR2_X1 U457 ( .A(n409), .B(n389), .ZN(n398) );
  XOR2_X1 U458 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n391) );
  NAND2_X1 U459 ( .A1(G227GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U460 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U461 ( .A(n392), .B(KEYINPUT84), .Z(n396) );
  XNOR2_X1 U462 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U463 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U464 ( .A(KEYINPUT92), .B(KEYINPUT78), .Z(n403) );
  XOR2_X1 U465 ( .A(G211GAT), .B(KEYINPUT21), .Z(n400) );
  XNOR2_X1 U466 ( .A(G197GAT), .B(G218GAT), .ZN(n399) );
  XNOR2_X1 U467 ( .A(n400), .B(n399), .ZN(n421) );
  XNOR2_X1 U468 ( .A(n421), .B(n401), .ZN(n402) );
  XNOR2_X1 U469 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U470 ( .A(n405), .B(n404), .Z(n407) );
  NAND2_X1 U471 ( .A1(G226GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U472 ( .A(n407), .B(n406), .ZN(n408) );
  NAND2_X1 U473 ( .A1(n525), .A2(n515), .ZN(n425) );
  XOR2_X1 U474 ( .A(n413), .B(G204GAT), .Z(n419) );
  XNOR2_X1 U475 ( .A(n414), .B(KEYINPUT22), .ZN(n417) );
  XOR2_X1 U476 ( .A(KEYINPUT88), .B(KEYINPUT23), .Z(n416) );
  XNOR2_X1 U477 ( .A(KEYINPUT24), .B(KEYINPUT86), .ZN(n415) );
  INV_X1 U478 ( .A(n420), .ZN(n422) );
  XOR2_X1 U479 ( .A(n422), .B(n421), .Z(n423) );
  XNOR2_X1 U480 ( .A(n424), .B(n423), .ZN(n469) );
  NAND2_X1 U481 ( .A1(n425), .A2(n469), .ZN(n426) );
  XNOR2_X1 U482 ( .A(n426), .B(KEYINPUT96), .ZN(n427) );
  XNOR2_X1 U483 ( .A(n427), .B(KEYINPUT25), .ZN(n431) );
  XNOR2_X1 U484 ( .A(KEYINPUT27), .B(n515), .ZN(n434) );
  NOR2_X1 U485 ( .A1(n469), .A2(n525), .ZN(n429) );
  XNOR2_X1 U486 ( .A(KEYINPUT95), .B(KEYINPUT26), .ZN(n428) );
  XOR2_X1 U487 ( .A(n429), .B(n428), .Z(n566) );
  AND2_X1 U488 ( .A1(n434), .A2(n566), .ZN(n430) );
  NOR2_X1 U489 ( .A1(n431), .A2(n430), .ZN(n432) );
  XOR2_X1 U490 ( .A(KEYINPUT97), .B(n432), .Z(n433) );
  NOR2_X1 U491 ( .A1(n511), .A2(n433), .ZN(n441) );
  NAND2_X1 U492 ( .A1(n511), .A2(n434), .ZN(n435) );
  XNOR2_X1 U493 ( .A(n435), .B(KEYINPUT93), .ZN(n540) );
  XNOR2_X1 U494 ( .A(n469), .B(KEYINPUT68), .ZN(n436) );
  INV_X1 U495 ( .A(n519), .ZN(n437) );
  NAND2_X1 U496 ( .A1(n540), .A2(n437), .ZN(n527) );
  XOR2_X1 U497 ( .A(KEYINPUT85), .B(n525), .Z(n438) );
  NOR2_X1 U498 ( .A1(n527), .A2(n438), .ZN(n439) );
  XNOR2_X1 U499 ( .A(n439), .B(KEYINPUT94), .ZN(n440) );
  NOR2_X1 U500 ( .A1(n441), .A2(n440), .ZN(n442) );
  XNOR2_X1 U501 ( .A(KEYINPUT98), .B(n442), .ZN(n480) );
  NOR2_X1 U502 ( .A1(n563), .A2(n480), .ZN(n443) );
  NAND2_X1 U503 ( .A1(n581), .A2(n443), .ZN(n444) );
  XOR2_X1 U504 ( .A(KEYINPUT37), .B(n444), .Z(n510) );
  NOR2_X1 U505 ( .A1(n482), .A2(n510), .ZN(n446) );
  XNOR2_X1 U506 ( .A(KEYINPUT104), .B(KEYINPUT38), .ZN(n445) );
  XNOR2_X1 U507 ( .A(n446), .B(n445), .ZN(n495) );
  NAND2_X1 U508 ( .A1(n495), .A2(n511), .ZN(n450) );
  XOR2_X1 U509 ( .A(KEYINPUT39), .B(KEYINPUT105), .Z(n448) );
  XOR2_X1 U510 ( .A(n572), .B(KEYINPUT41), .Z(n545) );
  OR2_X1 U511 ( .A1(n568), .A2(n545), .ZN(n452) );
  XOR2_X1 U512 ( .A(KEYINPUT46), .B(KEYINPUT112), .Z(n451) );
  XNOR2_X1 U513 ( .A(n452), .B(n451), .ZN(n454) );
  INV_X1 U514 ( .A(n563), .ZN(n578) );
  NAND2_X1 U515 ( .A1(n553), .A2(n578), .ZN(n453) );
  XNOR2_X1 U516 ( .A(n455), .B(KEYINPUT47), .ZN(n461) );
  NAND2_X1 U517 ( .A1(n563), .A2(n581), .ZN(n457) );
  XNOR2_X1 U518 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n456) );
  XNOR2_X1 U519 ( .A(n457), .B(n456), .ZN(n458) );
  NAND2_X1 U520 ( .A1(n458), .A2(n572), .ZN(n459) );
  NOR2_X1 U521 ( .A1(n459), .A2(n555), .ZN(n460) );
  NOR2_X1 U522 ( .A1(n461), .A2(n460), .ZN(n463) );
  XNOR2_X1 U523 ( .A(KEYINPUT120), .B(n515), .ZN(n464) );
  NAND2_X1 U524 ( .A1(n524), .A2(n464), .ZN(n467) );
  INV_X1 U525 ( .A(KEYINPUT54), .ZN(n465) );
  NOR2_X1 U526 ( .A1(n511), .A2(n468), .ZN(n565) );
  NAND2_X1 U527 ( .A1(n469), .A2(n565), .ZN(n470) );
  XNOR2_X1 U528 ( .A(KEYINPUT55), .B(n470), .ZN(n471) );
  NAND2_X1 U529 ( .A1(n471), .A2(n525), .ZN(n473) );
  INV_X1 U530 ( .A(KEYINPUT122), .ZN(n472) );
  XNOR2_X1 U531 ( .A(n473), .B(n472), .ZN(n558) );
  NAND2_X1 U532 ( .A1(n558), .A2(n536), .ZN(n477) );
  XOR2_X1 U533 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n475) );
  INV_X1 U534 ( .A(G190GAT), .ZN(n474) );
  XOR2_X1 U535 ( .A(KEYINPUT34), .B(KEYINPUT101), .Z(n485) );
  NOR2_X1 U536 ( .A1(n536), .A2(n578), .ZN(n478) );
  XOR2_X1 U537 ( .A(KEYINPUT16), .B(n478), .Z(n479) );
  NOR2_X1 U538 ( .A1(n480), .A2(n479), .ZN(n481) );
  XNOR2_X1 U539 ( .A(KEYINPUT99), .B(n481), .ZN(n500) );
  NOR2_X1 U540 ( .A1(n482), .A2(n500), .ZN(n483) );
  XNOR2_X1 U541 ( .A(n483), .B(KEYINPUT100), .ZN(n492) );
  NAND2_X1 U542 ( .A1(n492), .A2(n511), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U544 ( .A(G1GAT), .B(n486), .ZN(G1324GAT) );
  NAND2_X1 U545 ( .A1(n492), .A2(n515), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n487), .B(KEYINPUT102), .ZN(n488) );
  XNOR2_X1 U547 ( .A(G8GAT), .B(n488), .ZN(G1325GAT) );
  XOR2_X1 U548 ( .A(KEYINPUT103), .B(KEYINPUT35), .Z(n490) );
  NAND2_X1 U549 ( .A1(n492), .A2(n525), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(n491) );
  XOR2_X1 U551 ( .A(G15GAT), .B(n491), .Z(G1326GAT) );
  NAND2_X1 U552 ( .A1(n492), .A2(n519), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n493), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U554 ( .A1(n515), .A2(n495), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n494), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT106), .B(KEYINPUT40), .Z(n497) );
  NAND2_X1 U557 ( .A1(n495), .A2(n525), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U559 ( .A(G43GAT), .B(n498), .Z(G1330GAT) );
  NAND2_X1 U560 ( .A1(n519), .A2(n495), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n499), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT42), .B(KEYINPUT107), .Z(n502) );
  INV_X1 U563 ( .A(n545), .ZN(n557) );
  NAND2_X1 U564 ( .A1(n557), .A2(n568), .ZN(n509) );
  NOR2_X1 U565 ( .A1(n500), .A2(n509), .ZN(n506) );
  NAND2_X1 U566 ( .A1(n506), .A2(n511), .ZN(n501) );
  XNOR2_X1 U567 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(n503), .ZN(G1332GAT) );
  NAND2_X1 U569 ( .A1(n515), .A2(n506), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n504), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U571 ( .A1(n525), .A2(n506), .ZN(n505) );
  XNOR2_X1 U572 ( .A(n505), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U573 ( .A(G78GAT), .B(KEYINPUT43), .Z(n508) );
  NAND2_X1 U574 ( .A1(n506), .A2(n519), .ZN(n507) );
  XNOR2_X1 U575 ( .A(n508), .B(n507), .ZN(G1335GAT) );
  XOR2_X1 U576 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n513) );
  NOR2_X1 U577 ( .A1(n510), .A2(n509), .ZN(n520) );
  NAND2_X1 U578 ( .A1(n520), .A2(n511), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U580 ( .A(G85GAT), .B(n514), .ZN(G1336GAT) );
  NAND2_X1 U581 ( .A1(n515), .A2(n520), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n516), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U583 ( .A1(n525), .A2(n520), .ZN(n517) );
  XNOR2_X1 U584 ( .A(n517), .B(KEYINPUT110), .ZN(n518) );
  XNOR2_X1 U585 ( .A(G99GAT), .B(n518), .ZN(G1338GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n522) );
  NAND2_X1 U587 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  NAND2_X1 U590 ( .A1(n524), .A2(n525), .ZN(n526) );
  NOR2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n537) );
  NAND2_X1 U592 ( .A1(n537), .A2(n555), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n528), .B(KEYINPUT114), .ZN(n529) );
  XNOR2_X1 U594 ( .A(G113GAT), .B(n529), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(G120GAT), .B(KEYINPUT49), .Z(n531) );
  NAND2_X1 U596 ( .A1(n537), .A2(n557), .ZN(n530) );
  XNOR2_X1 U597 ( .A(n531), .B(n530), .ZN(G1341GAT) );
  XNOR2_X1 U598 ( .A(G127GAT), .B(KEYINPUT116), .ZN(n535) );
  XOR2_X1 U599 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n533) );
  NAND2_X1 U600 ( .A1(n537), .A2(n563), .ZN(n532) );
  XNOR2_X1 U601 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(G1342GAT) );
  XOR2_X1 U603 ( .A(G134GAT), .B(KEYINPUT51), .Z(n539) );
  NAND2_X1 U604 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(G1343GAT) );
  NAND2_X1 U606 ( .A1(n524), .A2(n540), .ZN(n542) );
  INV_X1 U607 ( .A(n566), .ZN(n541) );
  NOR2_X1 U608 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n543), .B(KEYINPUT117), .ZN(n552) );
  NOR2_X1 U610 ( .A1(n568), .A2(n552), .ZN(n544) );
  XOR2_X1 U611 ( .A(G141GAT), .B(n544), .Z(G1344GAT) );
  NOR2_X1 U612 ( .A1(n545), .A2(n552), .ZN(n550) );
  XOR2_X1 U613 ( .A(KEYINPUT119), .B(KEYINPUT53), .Z(n547) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U616 ( .A(KEYINPUT118), .B(n548), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(G1345GAT) );
  NOR2_X1 U618 ( .A1(n578), .A2(n552), .ZN(n551) );
  XOR2_X1 U619 ( .A(G155GAT), .B(n551), .Z(G1346GAT) );
  NOR2_X1 U620 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U621 ( .A(G162GAT), .B(n554), .Z(G1347GAT) );
  NAND2_X1 U622 ( .A1(n558), .A2(n555), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n560) );
  XOR2_X1 U625 ( .A(G176GAT), .B(KEYINPUT56), .Z(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(n562) );
  XOR2_X1 U627 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1349GAT) );
  NAND2_X1 U629 ( .A1(n558), .A2(n563), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U632 ( .A(KEYINPUT125), .B(n567), .ZN(n580) );
  INV_X1 U633 ( .A(n580), .ZN(n577) );
  NOR2_X1 U634 ( .A1(n568), .A2(n577), .ZN(n570) );
  XNOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(n571), .ZN(G1352GAT) );
  NOR2_X1 U638 ( .A1(n577), .A2(n572), .ZN(n576) );
  XOR2_X1 U639 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n574) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT127), .ZN(n573) );
  XNOR2_X1 U641 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(G1353GAT) );
  NOR2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U644 ( .A(G211GAT), .B(n579), .Z(G1354GAT) );
  NAND2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(n582), .B(KEYINPUT62), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

