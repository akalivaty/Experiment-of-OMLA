//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 0 0 0 1 1 1 0 0 0 1 0 0 1 1 1 1 0 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 0 0 0 0 1 1 1 1 0 1 1 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:03 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n572,
    new_n573, new_n574, new_n575, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n593, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n629, new_n630, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AND2_X1   g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n459), .A2(KEYINPUT68), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n456), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(KEYINPUT68), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n465), .A2(G2105), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n470), .A2(G137), .B1(G101), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n473), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n476), .A2(KEYINPUT69), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n476), .A2(KEYINPUT69), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n472), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n482), .ZN(new_n483));
  XOR2_X1   g058(.A(new_n483), .B(KEYINPUT71), .Z(new_n484));
  AND2_X1   g059(.A1(new_n466), .A2(new_n468), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(new_n482), .ZN(new_n486));
  INV_X1    g061(.A(G136), .ZN(new_n487));
  OR3_X1    g062(.A1(new_n486), .A2(KEYINPUT70), .A3(new_n487), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n469), .A2(new_n482), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  OAI21_X1  g065(.A(KEYINPUT70), .B1(new_n486), .B2(new_n487), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n484), .A2(new_n488), .A3(new_n490), .A4(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT4), .B1(new_n486), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n470), .A2(new_n496), .A3(G138), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n495), .A2(new_n497), .B1(G126), .B2(new_n489), .ZN(new_n498));
  OR2_X1    g073(.A1(G102), .A2(G2105), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n499), .B(G2104), .C1(G114), .C2(new_n482), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT73), .B1(new_n505), .B2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(new_n503), .A3(G543), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n504), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT72), .B(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT6), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G651), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n509), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n511), .A2(G543), .A3(new_n513), .ZN(new_n516));
  INV_X1    g091(.A(G50), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n514), .A2(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n519), .A2(new_n510), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n518), .A2(new_n520), .ZN(G166));
  INV_X1    g096(.A(new_n504), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n507), .B1(new_n503), .B2(G543), .ZN(new_n523));
  NOR3_X1   g098(.A1(new_n505), .A2(KEYINPUT73), .A3(KEYINPUT5), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT74), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n509), .A2(KEYINPUT74), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AND3_X1   g104(.A1(new_n529), .A2(G63), .A3(G651), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  INV_X1    g107(.A(G51), .ZN(new_n533));
  INV_X1    g108(.A(G89), .ZN(new_n534));
  OAI221_X1 g109(.A(new_n532), .B1(new_n516), .B2(new_n533), .C1(new_n534), .C2(new_n514), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n530), .A2(new_n535), .ZN(G168));
  INV_X1    g111(.A(new_n514), .ZN(new_n537));
  XOR2_X1   g112(.A(KEYINPUT76), .B(G90), .Z(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n516), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G52), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT75), .ZN(new_n542));
  AOI211_X1 g117(.A(new_n526), .B(new_n504), .C1(new_n506), .C2(new_n508), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n506), .A2(new_n508), .ZN(new_n544));
  AOI21_X1  g119(.A(KEYINPUT74), .B1(new_n544), .B2(new_n522), .ZN(new_n545));
  OAI21_X1  g120(.A(G64), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(G77), .A2(G543), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n510), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n542), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI211_X1 g125(.A(KEYINPUT75), .B(new_n510), .C1(new_n546), .C2(new_n547), .ZN(new_n551));
  OAI211_X1 g126(.A(new_n539), .B(new_n541), .C1(new_n550), .C2(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  OAI21_X1  g128(.A(G56), .B1(new_n543), .B2(new_n545), .ZN(new_n554));
  NAND2_X1  g129(.A1(G68), .A2(G543), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n510), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND4_X1  g131(.A1(new_n509), .A2(new_n511), .A3(G81), .A4(new_n513), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n511), .A2(G43), .A3(G543), .A4(new_n513), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NOR3_X1   g134(.A1(new_n556), .A2(KEYINPUT77), .A3(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT77), .ZN(new_n561));
  INV_X1    g136(.A(G56), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n562), .B1(new_n527), .B2(new_n528), .ZN(new_n563));
  INV_X1    g138(.A(new_n555), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n549), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n559), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n561), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n560), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(G153));
  NAND4_X1  g145(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g146(.A(KEYINPUT78), .B(KEYINPUT8), .Z(new_n572));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n572), .B(new_n573), .ZN(new_n574));
  NAND4_X1  g149(.A1(G319), .A2(G483), .A3(G661), .A4(new_n574), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT79), .ZN(G188));
  XOR2_X1   g151(.A(KEYINPUT81), .B(G65), .Z(new_n577));
  NAND2_X1  g152(.A1(new_n509), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(G78), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n579), .B2(new_n505), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT82), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI211_X1 g157(.A(new_n578), .B(KEYINPUT82), .C1(new_n579), .C2(new_n505), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n582), .A2(G651), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n537), .A2(G91), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n511), .A2(G53), .A3(G543), .A4(new_n513), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT9), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n587), .A2(KEYINPUT80), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n586), .B(new_n588), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n584), .A2(new_n585), .A3(new_n589), .ZN(G299));
  INV_X1    g165(.A(G168), .ZN(G286));
  XOR2_X1   g166(.A(G166), .B(KEYINPUT83), .Z(G303));
  AOI22_X1  g167(.A1(G87), .A2(new_n537), .B1(new_n540), .B2(G49), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n529), .B2(G74), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g170(.A(new_n595), .B(KEYINPUT84), .Z(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G288));
  AOI22_X1  g172(.A1(new_n509), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n598), .A2(new_n510), .ZN(new_n599));
  INV_X1    g174(.A(G48), .ZN(new_n600));
  INV_X1    g175(.A(G86), .ZN(new_n601));
  OAI221_X1 g176(.A(new_n599), .B1(new_n600), .B2(new_n516), .C1(new_n601), .C2(new_n514), .ZN(G305));
  AOI22_X1  g177(.A1(new_n529), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n603), .A2(new_n510), .ZN(new_n604));
  INV_X1    g179(.A(G85), .ZN(new_n605));
  INV_X1    g180(.A(G47), .ZN(new_n606));
  OAI22_X1  g181(.A1(new_n514), .A2(new_n605), .B1(new_n516), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(new_n511), .A2(new_n513), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  NAND4_X1  g187(.A1(new_n611), .A2(new_n612), .A3(G92), .A4(new_n509), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n540), .A2(G54), .ZN(new_n614));
  INV_X1    g189(.A(G92), .ZN(new_n615));
  OAI21_X1  g190(.A(KEYINPUT10), .B1(new_n514), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(G79), .A2(G543), .ZN(new_n617));
  XOR2_X1   g192(.A(KEYINPUT85), .B(G66), .Z(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n525), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G651), .ZN(new_n620));
  NAND4_X1  g195(.A1(new_n613), .A2(new_n614), .A3(new_n616), .A4(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(G868), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G171), .B2(new_n622), .ZN(G284));
  OAI21_X1  g199(.A(new_n623), .B1(G171), .B2(new_n622), .ZN(G321));
  NAND2_X1  g200(.A1(G299), .A2(new_n622), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(new_n622), .B2(G168), .ZN(G297));
  OAI21_X1  g202(.A(new_n626), .B1(new_n622), .B2(G168), .ZN(G280));
  INV_X1    g203(.A(new_n621), .ZN(new_n629));
  INV_X1    g204(.A(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(G860), .ZN(G148));
  NAND2_X1  g206(.A1(new_n568), .A2(new_n622), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n621), .A2(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(new_n622), .B2(new_n633), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g210(.A1(new_n485), .A2(new_n471), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT13), .Z(new_n638));
  OR2_X1    g213(.A1(new_n638), .A2(G2100), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n489), .A2(G123), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n470), .A2(G135), .ZN(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n482), .A2(G111), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n640), .B(new_n641), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(G2096), .Z(new_n645));
  NAND2_X1  g220(.A1(new_n638), .A2(G2100), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n639), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT86), .Z(G156));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT15), .ZN(new_n653));
  INV_X1    g228(.A(G2435), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(KEYINPUT14), .ZN(new_n656));
  XOR2_X1   g231(.A(G2443), .B(G2446), .Z(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1341), .B(G1348), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n657), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n655), .A2(KEYINPUT14), .A3(new_n662), .ZN(new_n663));
  AND3_X1   g238(.A1(new_n658), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n661), .B1(new_n658), .B2(new_n663), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n650), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n658), .A2(new_n663), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(new_n660), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n658), .A2(new_n661), .A3(new_n663), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(new_n649), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n666), .A2(new_n670), .A3(G14), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(KEYINPUT87), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT87), .ZN(new_n673));
  NAND4_X1  g248(.A1(new_n666), .A2(new_n670), .A3(new_n673), .A4(G14), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(G401));
  XOR2_X1   g251(.A(G2084), .B(G2090), .Z(new_n677));
  XNOR2_X1  g252(.A(G2072), .B(G2078), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2067), .B(G2678), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT18), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n678), .B(KEYINPUT17), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(new_n677), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n678), .A2(new_n679), .ZN(new_n685));
  AOI211_X1 g260(.A(new_n677), .B(new_n685), .C1(new_n682), .C2(new_n679), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n686), .A2(KEYINPUT88), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(KEYINPUT88), .ZN(new_n688));
  OAI221_X1 g263(.A(new_n681), .B1(new_n679), .B2(new_n684), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT89), .ZN(new_n690));
  XNOR2_X1  g265(.A(G2096), .B(G2100), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(G227));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  INV_X1    g268(.A(G1981), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(G1991), .ZN(new_n696));
  INV_X1    g271(.A(G1996), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G1971), .B(G1976), .Z(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(G1956), .B(G2474), .Z(new_n702));
  XOR2_X1   g277(.A(G1961), .B(G1966), .Z(new_n703));
  AND2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT20), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n702), .A2(new_n703), .ZN(new_n707));
  AOI22_X1  g282(.A1(new_n705), .A2(new_n706), .B1(new_n701), .B2(new_n707), .ZN(new_n708));
  OR3_X1    g283(.A1(new_n701), .A2(new_n704), .A3(new_n707), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n708), .B(new_n709), .C1(new_n706), .C2(new_n705), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n698), .B(new_n710), .Z(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT91), .B(G1986), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(G229));
  INV_X1    g289(.A(G16), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G6), .ZN(new_n716));
  INV_X1    g291(.A(G305), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n716), .B1(new_n717), .B2(new_n715), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT32), .B(G1981), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT95), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n718), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n715), .A2(G23), .ZN(new_n722));
  INV_X1    g297(.A(new_n595), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n723), .B2(new_n715), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT33), .B(G1976), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G22), .ZN(new_n727));
  OAI21_X1  g302(.A(KEYINPUT96), .B1(new_n727), .B2(G16), .ZN(new_n728));
  OR3_X1    g303(.A1(new_n727), .A2(KEYINPUT96), .A3(G16), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n728), .B(new_n729), .C1(G166), .C2(new_n715), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT97), .B(G1971), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n721), .A2(new_n726), .A3(new_n732), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT34), .Z(new_n734));
  NOR2_X1   g309(.A1(G16), .A2(G24), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(new_n608), .B2(G16), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT94), .B(G1986), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G29), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G25), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n489), .A2(G119), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT92), .Z(new_n742));
  INV_X1    g317(.A(G131), .ZN(new_n743));
  OAI21_X1  g318(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n482), .A2(G107), .ZN(new_n745));
  OAI22_X1  g320(.A1(new_n486), .A2(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n740), .B1(new_n747), .B2(new_n739), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT35), .B(G1991), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT93), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n748), .B(new_n750), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n734), .A2(new_n738), .A3(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT36), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT99), .B(KEYINPUT25), .Z(new_n755));
  NAND2_X1  g330(.A1(new_n471), .A2(G103), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n470), .A2(G139), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n485), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n757), .B(new_n758), .C1(new_n482), .C2(new_n759), .ZN(new_n760));
  MUX2_X1   g335(.A(G33), .B(new_n760), .S(G29), .Z(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT100), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(G2072), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT101), .ZN(new_n764));
  AOI22_X1  g339(.A1(G129), .A2(new_n489), .B1(new_n470), .B2(G141), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n471), .A2(G105), .ZN(new_n766));
  NAND3_X1  g341(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT26), .Z(new_n768));
  NAND3_X1  g343(.A1(new_n765), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT102), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n770), .A2(G29), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G29), .B2(G32), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT27), .B(G1996), .Z(new_n774));
  NOR2_X1   g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT103), .ZN(new_n776));
  AOI211_X1 g351(.A(new_n764), .B(new_n776), .C1(new_n773), .C2(new_n774), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n644), .A2(new_n739), .ZN(new_n778));
  INV_X1    g353(.A(G11), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n778), .B1(KEYINPUT31), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(KEYINPUT31), .B2(new_n779), .ZN(new_n781));
  NAND2_X1  g356(.A1(G168), .A2(G16), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G16), .B2(G21), .ZN(new_n783));
  INV_X1    g358(.A(G1966), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(G29), .A2(G35), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G162), .B2(G29), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT105), .B(KEYINPUT29), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(G2090), .ZN(new_n790));
  AOI211_X1 g365(.A(new_n781), .B(new_n785), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(G171), .A2(G16), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G5), .B2(G16), .ZN(new_n793));
  INV_X1    g368(.A(G1961), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n791), .A2(new_n795), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n793), .A2(new_n794), .B1(new_n784), .B2(new_n783), .ZN(new_n797));
  NOR2_X1   g372(.A1(G27), .A2(G29), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G164), .B2(G29), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G2078), .ZN(new_n800));
  NAND2_X1  g375(.A1(G299), .A2(G16), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n715), .A2(KEYINPUT23), .A3(G20), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT23), .ZN(new_n803));
  INV_X1    g378(.A(G20), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(G16), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n801), .A2(new_n802), .A3(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G1956), .ZN(new_n807));
  INV_X1    g382(.A(G28), .ZN(new_n808));
  AOI21_X1  g383(.A(G29), .B1(new_n808), .B2(KEYINPUT30), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n808), .A2(KEYINPUT30), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT104), .ZN(new_n811));
  AOI211_X1 g386(.A(new_n800), .B(new_n807), .C1(new_n809), .C2(new_n811), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n777), .A2(new_n796), .A3(new_n797), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n715), .A2(G19), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n569), .B2(new_n715), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(G1341), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT28), .ZN(new_n817));
  INV_X1    g392(.A(G26), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(G29), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n818), .A2(G29), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n489), .A2(G128), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n470), .A2(G140), .ZN(new_n822));
  OAI21_X1  g397(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n482), .A2(G116), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n821), .B(new_n822), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n820), .B1(new_n825), .B2(G29), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n819), .B1(new_n826), .B2(new_n817), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n815), .A2(G1341), .B1(G2067), .B2(new_n827), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n827), .A2(G2067), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n715), .A2(G4), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n629), .B2(new_n715), .ZN(new_n831));
  INV_X1    g406(.A(G1348), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n816), .A2(new_n828), .A3(new_n829), .A4(new_n833), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT98), .Z(new_n835));
  NOR3_X1   g410(.A1(new_n754), .A2(new_n813), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n789), .A2(new_n790), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT106), .Z(new_n838));
  OR2_X1    g413(.A1(new_n762), .A2(G2072), .ZN(new_n839));
  AND2_X1   g414(.A1(KEYINPUT24), .A2(G34), .ZN(new_n840));
  NOR2_X1   g415(.A1(KEYINPUT24), .A2(G34), .ZN(new_n841));
  NOR3_X1   g416(.A1(new_n840), .A2(new_n841), .A3(G29), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n842), .B1(new_n479), .B2(G29), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(G2084), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n836), .A2(new_n838), .A3(new_n839), .A4(new_n844), .ZN(G150));
  INV_X1    g420(.A(G150), .ZN(G311));
  INV_X1    g421(.A(G93), .ZN(new_n847));
  INV_X1    g422(.A(G55), .ZN(new_n848));
  OAI22_X1  g423(.A1(new_n514), .A2(new_n847), .B1(new_n516), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(G67), .B1(new_n543), .B2(new_n545), .ZN(new_n850));
  NAND2_X1  g425(.A1(G80), .A2(G543), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n849), .B1(new_n852), .B2(new_n549), .ZN(new_n853));
  INV_X1    g428(.A(G860), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT37), .ZN(new_n856));
  OAI21_X1  g431(.A(KEYINPUT77), .B1(new_n556), .B2(new_n559), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n564), .B1(new_n529), .B2(G56), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n561), .B(new_n566), .C1(new_n858), .C2(new_n510), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n853), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n849), .ZN(new_n861));
  AOI22_X1  g436(.A1(new_n529), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n861), .B1(new_n862), .B2(new_n510), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n554), .A2(new_n555), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n559), .B1(new_n864), .B2(new_n549), .ZN(new_n865));
  OAI21_X1  g440(.A(KEYINPUT107), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n860), .A2(new_n866), .ZN(new_n867));
  AOI211_X1 g442(.A(KEYINPUT107), .B(new_n853), .C1(new_n857), .C2(new_n859), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n621), .A2(new_n630), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT38), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n869), .B(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT39), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT108), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n854), .B1(new_n872), .B2(new_n873), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n856), .B1(new_n875), .B2(new_n876), .ZN(G145));
  XNOR2_X1  g452(.A(new_n760), .B(new_n637), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n825), .B(KEYINPUT109), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n470), .A2(G142), .ZN(new_n881));
  OAI21_X1  g456(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n482), .A2(G118), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n884), .B1(G130), .B2(new_n489), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n747), .B(new_n885), .Z(new_n886));
  XNOR2_X1  g461(.A(new_n880), .B(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n479), .B(new_n644), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(new_n492), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n770), .B(new_n501), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n890), .A2(new_n891), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n888), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n892), .A2(new_n893), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(new_n887), .ZN(new_n896));
  INV_X1    g471(.A(G37), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n894), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g474(.A1(new_n853), .A2(G868), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n608), .B(KEYINPUT110), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n595), .B(G166), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(G305), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n904), .A2(G305), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n903), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n907), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n909), .A2(new_n902), .A3(new_n905), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT42), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n869), .B(new_n633), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n629), .A2(new_n585), .A3(new_n584), .A4(new_n589), .ZN(new_n914));
  NAND2_X1  g489(.A1(G299), .A2(new_n621), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n914), .A2(new_n915), .A3(KEYINPUT41), .ZN(new_n918));
  AOI21_X1  g493(.A(KEYINPUT41), .B1(new_n914), .B2(new_n915), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n917), .B1(new_n913), .B2(new_n920), .ZN(new_n921));
  XOR2_X1   g496(.A(new_n912), .B(new_n921), .Z(new_n922));
  OAI21_X1  g497(.A(new_n901), .B1(new_n922), .B2(new_n622), .ZN(G331));
  XOR2_X1   g498(.A(G331), .B(KEYINPUT111), .Z(G295));
  XOR2_X1   g499(.A(KEYINPUT112), .B(KEYINPUT43), .Z(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n863), .B1(new_n560), .B2(new_n567), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT107), .ZN(new_n928));
  INV_X1    g503(.A(new_n865), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n928), .B1(new_n929), .B2(new_n853), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n860), .A2(new_n928), .ZN(new_n932));
  AOI22_X1  g507(.A1(new_n529), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT75), .B1(new_n933), .B2(new_n510), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n548), .A2(new_n542), .A3(new_n549), .ZN(new_n935));
  AOI22_X1  g510(.A1(new_n934), .A2(new_n935), .B1(G52), .B2(new_n540), .ZN(new_n936));
  AOI21_X1  g511(.A(G168), .B1(new_n936), .B2(new_n539), .ZN(new_n937));
  NOR2_X1   g512(.A1(G301), .A2(G286), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n931), .B(new_n932), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(G301), .A2(G286), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n936), .A2(G168), .A3(new_n539), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n940), .B(new_n941), .C1(new_n867), .C2(new_n868), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n939), .A2(new_n942), .A3(new_n920), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT113), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n939), .A2(new_n942), .ZN(new_n946));
  INV_X1    g521(.A(new_n916), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n939), .A2(new_n942), .A3(KEYINPUT113), .A4(new_n920), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n945), .A2(new_n948), .A3(new_n911), .A4(new_n949), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n950), .A2(new_n897), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n945), .A2(new_n948), .A3(new_n949), .ZN(new_n952));
  INV_X1    g527(.A(new_n911), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n926), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n948), .A2(new_n943), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n953), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n957), .A2(new_n950), .A3(new_n897), .A4(new_n926), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  NOR3_X1   g534(.A1(new_n955), .A2(KEYINPUT44), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n951), .A2(new_n957), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT43), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n951), .A2(new_n954), .A3(new_n926), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n960), .B1(KEYINPUT44), .B2(new_n964), .ZN(G397));
  INV_X1    g540(.A(G1384), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n501), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI211_X1 g544(.A(G40), .B(new_n472), .C1(new_n477), .C2(new_n478), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n825), .B(G2067), .ZN(new_n973));
  INV_X1    g548(.A(new_n770), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n973), .B1(new_n974), .B2(G1996), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n971), .A2(new_n697), .ZN(new_n977));
  XOR2_X1   g552(.A(new_n977), .B(KEYINPUT114), .Z(new_n978));
  AOI21_X1  g553(.A(new_n976), .B1(new_n978), .B2(new_n770), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n747), .B(new_n749), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n979), .B1(new_n972), .B2(new_n980), .ZN(new_n981));
  OR2_X1    g556(.A1(G290), .A2(G1986), .ZN(new_n982));
  NAND2_X1  g557(.A1(G290), .A2(G1986), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n972), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n967), .A2(new_n970), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(G8), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(G1976), .B2(new_n723), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n990));
  OR2_X1    g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(G305), .B(KEYINPUT49), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT116), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n694), .B1(new_n599), .B2(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n992), .B(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n995), .A2(G8), .A3(new_n987), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n596), .A2(G1976), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n989), .A2(new_n990), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n991), .B(new_n996), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n970), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n966), .ZN(new_n1001));
  AND3_X1   g576(.A1(new_n969), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(KEYINPUT56), .B(G2072), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g579(.A(G299), .B(KEYINPUT57), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n967), .A2(KEYINPUT50), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT50), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n501), .A2(new_n1008), .A3(new_n966), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n1007), .A2(new_n1000), .A3(new_n1009), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1004), .B(new_n1006), .C1(G1956), .C2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1011), .A2(KEYINPUT61), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT60), .ZN(new_n1013));
  OAI22_X1  g588(.A1(new_n1010), .A2(G1348), .B1(G2067), .B2(new_n987), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT119), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1007), .A2(new_n1000), .A3(new_n1009), .ZN(new_n1017));
  INV_X1    g592(.A(G2067), .ZN(new_n1018));
  AOI22_X1  g593(.A1(new_n1017), .A2(new_n832), .B1(new_n1018), .B2(new_n986), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT119), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1013), .B1(new_n1016), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1012), .B1(new_n1021), .B2(new_n621), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1020), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1019), .A2(KEYINPUT119), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT60), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1016), .A2(new_n1013), .A3(new_n1020), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(new_n629), .A3(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n969), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1028));
  XNOR2_X1  g603(.A(KEYINPUT58), .B(G1341), .ZN(new_n1029));
  OAI22_X1  g604(.A1(new_n1028), .A2(G1996), .B1(new_n986), .B2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1030), .A2(KEYINPUT120), .A3(KEYINPUT59), .A4(new_n569), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT61), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT121), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1030), .A2(new_n569), .ZN(new_n1034));
  XOR2_X1   g609(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n1035));
  AOI22_X1  g610(.A1(new_n1011), .A2(new_n1033), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1022), .A2(new_n1027), .A3(new_n1031), .A4(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1004), .B1(G1956), .B2(new_n1010), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n1005), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1011), .A2(new_n1016), .A3(new_n629), .A4(new_n1020), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1037), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1042), .B1(new_n1028), .B2(G2078), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1017), .A2(new_n794), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OR3_X1    g620(.A1(new_n1028), .A2(new_n1042), .A3(G2078), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1045), .A2(G301), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n472), .ZN(new_n1048));
  NOR3_X1   g623(.A1(new_n1048), .A2(new_n1042), .A3(G2078), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n476), .A2(G40), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n969), .A2(new_n1001), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n1045), .A2(new_n1051), .ZN(new_n1052));
  OAI211_X1 g627(.A(KEYINPUT54), .B(new_n1047), .C1(new_n1052), .C2(G301), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT122), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT51), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(G286), .A2(G8), .ZN(new_n1058));
  INV_X1    g633(.A(G2084), .ZN(new_n1059));
  AOI22_X1  g634(.A1(new_n1010), .A2(new_n1059), .B1(new_n1028), .B2(new_n784), .ZN(new_n1060));
  INV_X1    g635(.A(G8), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1057), .B(new_n1058), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1062));
  OAI22_X1  g637(.A1(new_n1002), .A2(G1966), .B1(G2084), .B2(new_n1017), .ZN(new_n1063));
  OAI211_X1 g638(.A(G8), .B(new_n1056), .C1(new_n1063), .C2(G286), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1062), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1063), .A2(G8), .A3(G286), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(G303), .A2(G8), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n1069), .B(KEYINPUT55), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1010), .A2(new_n790), .ZN(new_n1071));
  INV_X1    g646(.A(G1971), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1028), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1071), .A2(KEYINPUT118), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(G8), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT118), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1070), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n1079));
  AOI21_X1  g654(.A(G301), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1080));
  AND4_X1   g655(.A1(G301), .A2(new_n1043), .A3(new_n1044), .A4(new_n1051), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1079), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT123), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  OAI211_X1 g659(.A(KEYINPUT123), .B(new_n1079), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1078), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1041), .A2(new_n1053), .A3(new_n1068), .A4(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1070), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT115), .B1(new_n1028), .B2(new_n1072), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT115), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1071), .B1(new_n1090), .B2(new_n1073), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1088), .B(G8), .C1(new_n1089), .C2(new_n1091), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n1092), .A2(new_n1077), .A3(new_n1080), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1066), .A2(KEYINPUT62), .A3(new_n1067), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT62), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1093), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT63), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1060), .A2(new_n1061), .A3(G286), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1077), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1096), .A2(new_n1099), .A3(new_n1092), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n999), .B1(new_n1087), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1098), .ZN(new_n1102));
  OAI21_X1  g677(.A(G8), .B1(new_n1091), .B2(new_n1089), .ZN(new_n1103));
  AOI211_X1 g678(.A(new_n1102), .B(new_n999), .C1(new_n1070), .C2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(G288), .A2(G1976), .ZN(new_n1105));
  XOR2_X1   g680(.A(new_n1105), .B(KEYINPUT117), .Z(new_n1106));
  AOI22_X1  g681(.A1(new_n1106), .A2(new_n996), .B1(new_n694), .B2(new_n717), .ZN(new_n1107));
  OAI22_X1  g682(.A1(new_n1104), .A2(new_n1097), .B1(new_n988), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n985), .B1(new_n1101), .B2(new_n1108), .ZN(new_n1109));
  XOR2_X1   g684(.A(new_n978), .B(KEYINPUT46), .Z(new_n1110));
  OAI21_X1  g685(.A(new_n971), .B1(new_n974), .B2(new_n973), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1112), .B(KEYINPUT47), .ZN(new_n1113));
  INV_X1    g688(.A(new_n749), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n979), .A2(new_n747), .A3(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n825), .A2(G2067), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n971), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n982), .A2(new_n972), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1118), .B(KEYINPUT124), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n1119), .B(KEYINPUT48), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1113), .B(new_n1117), .C1(new_n981), .C2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1109), .A2(new_n1122), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g698(.A1(G227), .A2(new_n463), .ZN(new_n1125));
  INV_X1    g699(.A(KEYINPUT125), .ZN(new_n1126));
  OAI21_X1  g700(.A(new_n713), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g701(.A(new_n1127), .ZN(new_n1128));
  NAND2_X1  g702(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1129));
  AND3_X1   g703(.A1(new_n675), .A2(new_n898), .A3(new_n1129), .ZN(new_n1130));
  OAI211_X1 g704(.A(new_n1128), .B(new_n1130), .C1(new_n955), .C2(new_n959), .ZN(new_n1131));
  INV_X1    g705(.A(KEYINPUT126), .ZN(new_n1132));
  NOR2_X1   g706(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  AND2_X1   g707(.A1(new_n952), .A2(new_n953), .ZN(new_n1134));
  NAND2_X1  g708(.A1(new_n950), .A2(new_n897), .ZN(new_n1135));
  OAI21_X1  g709(.A(new_n925), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g710(.A(new_n1127), .B1(new_n1136), .B2(new_n958), .ZN(new_n1137));
  AOI21_X1  g711(.A(KEYINPUT126), .B1(new_n1137), .B2(new_n1130), .ZN(new_n1138));
  OAI21_X1  g712(.A(KEYINPUT127), .B1(new_n1133), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g713(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1140));
  NAND3_X1  g714(.A1(new_n1137), .A2(KEYINPUT126), .A3(new_n1130), .ZN(new_n1141));
  INV_X1    g715(.A(KEYINPUT127), .ZN(new_n1142));
  NAND3_X1  g716(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g717(.A1(new_n1139), .A2(new_n1143), .ZN(G308));
  NAND2_X1  g718(.A1(new_n1140), .A2(new_n1141), .ZN(G225));
endmodule


