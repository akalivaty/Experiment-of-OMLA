//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 1 1 0 1 1 1 1 1 1 1 0 0 1 0 1 0 1 0 0 0 1 0 1 0 1 1 1 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1286, new_n1287, new_n1288, new_n1289, new_n1291,
    new_n1292, new_n1293, new_n1294, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT65), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND3_X1  g0013(.A1(new_n211), .A2(G20), .A3(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  INV_X1    g0021(.A(G77), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  INV_X1    g0023(.A(G107), .ZN(new_n224));
  INV_X1    g0024(.A(G264), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n206), .B1(new_n220), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n209), .B(new_n214), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  INV_X1    g0037(.A(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n234), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XOR2_X1   g0043(.A(G50), .B(G58), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(KEYINPUT10), .ZN(new_n247));
  INV_X1    g0047(.A(G1), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n248), .B1(G41), .B2(G45), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G1), .A3(G13), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n250), .A2(new_n252), .A3(G274), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n249), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n254), .B1(G226), .B2(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT3), .B(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G222), .A2(G1698), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(G223), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n258), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n252), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n262), .B(new_n263), .C1(G77), .C2(new_n258), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n257), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G190), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G200), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n268), .B1(new_n257), .B2(new_n264), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  XOR2_X1   g0070(.A(KEYINPUT8), .B(G58), .Z(new_n271));
  INV_X1    g0071(.A(G20), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G33), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(G20), .A2(G33), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n271), .A2(new_n274), .B1(G150), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n203), .A2(G20), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n212), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n248), .A2(G13), .A3(G20), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(new_n280), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n248), .A2(G20), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G50), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n284), .A2(new_n288), .B1(new_n287), .B2(new_n283), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n281), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(KEYINPUT9), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT9), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n281), .A2(new_n292), .A3(new_n289), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n247), .B1(new_n270), .B2(new_n294), .ZN(new_n295));
  NOR3_X1   g0095(.A1(new_n267), .A2(KEYINPUT10), .A3(new_n269), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT67), .ZN(new_n297));
  AND3_X1   g0097(.A1(new_n291), .A2(new_n297), .A3(new_n293), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n297), .B1(new_n291), .B2(new_n293), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n296), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT68), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI211_X1 g0102(.A(KEYINPUT68), .B(new_n296), .C1(new_n298), .C2(new_n299), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n295), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT18), .ZN(new_n305));
  OAI21_X1  g0105(.A(KEYINPUT7), .B1(new_n258), .B2(G20), .ZN(new_n306));
  INV_X1    g0106(.A(G33), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT3), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT3), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G33), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT73), .B(KEYINPUT7), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n311), .A2(new_n312), .A3(new_n272), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n306), .A2(new_n313), .A3(G68), .ZN(new_n314));
  INV_X1    g0114(.A(G58), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n315), .A2(new_n216), .ZN(new_n316));
  OAI21_X1  g0116(.A(G20), .B1(new_n316), .B2(new_n202), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n275), .A2(G159), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n314), .A2(new_n320), .A3(KEYINPUT16), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT74), .ZN(new_n322));
  AOI21_X1  g0122(.A(G20), .B1(new_n308), .B2(new_n310), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n216), .B1(new_n323), .B2(new_n312), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n319), .B1(new_n324), .B2(new_n306), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT74), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n325), .A2(new_n326), .A3(KEYINPUT16), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n322), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n280), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n311), .A2(new_n272), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT75), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(new_n309), .B2(G33), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n307), .A2(KEYINPUT75), .A3(KEYINPUT3), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n332), .A2(new_n310), .A3(new_n333), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n272), .A2(KEYINPUT7), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n330), .A2(new_n312), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n320), .B1(new_n336), .B2(new_n216), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT16), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n329), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n328), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n271), .A2(new_n285), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n271), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n342), .A2(new_n284), .B1(new_n343), .B2(new_n283), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  OR2_X1    g0145(.A1(G223), .A2(G1698), .ZN(new_n346));
  INV_X1    g0146(.A(G226), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G1698), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n349), .A2(new_n258), .B1(G33), .B2(G87), .ZN(new_n350));
  OAI21_X1  g0150(.A(KEYINPUT76), .B1(new_n350), .B2(new_n252), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n252), .A2(G274), .ZN(new_n352));
  OAI22_X1  g0152(.A1(new_n231), .A2(new_n255), .B1(new_n352), .B2(new_n249), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n353), .A2(G179), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n346), .A2(new_n348), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n355), .A2(new_n311), .B1(new_n307), .B2(new_n218), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT76), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n356), .A2(new_n357), .A3(new_n263), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n351), .A2(new_n354), .A3(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G169), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n350), .A2(new_n252), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n360), .B1(new_n361), .B2(new_n353), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n305), .B1(new_n345), .B2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n344), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n366), .B1(new_n328), .B2(new_n339), .ZN(new_n367));
  NOR3_X1   g0167(.A1(new_n367), .A2(KEYINPUT18), .A3(new_n363), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n353), .A2(G190), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n351), .A2(new_n370), .A3(new_n358), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n268), .B1(new_n361), .B2(new_n353), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT77), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n374), .A2(KEYINPUT17), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n374), .A2(KEYINPUT17), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n367), .B(new_n373), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  AOI221_X4 g0177(.A(new_n366), .B1(new_n371), .B2(new_n372), .C1(new_n328), .C2(new_n339), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n377), .B1(new_n378), .B2(new_n376), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n369), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT66), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n282), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n248), .A2(KEYINPUT66), .A3(G13), .A4(G20), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n384), .A2(G68), .A3(new_n329), .A4(new_n285), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT12), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n382), .A2(new_n383), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n386), .B1(new_n387), .B2(new_n216), .ZN(new_n388));
  INV_X1    g0188(.A(G13), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n389), .A2(G1), .ZN(new_n390));
  AND4_X1   g0190(.A1(new_n386), .A2(new_n390), .A3(G20), .A4(new_n216), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n385), .B1(new_n388), .B2(new_n391), .ZN(new_n392));
  OAI22_X1  g0192(.A1(new_n273), .A2(new_n222), .B1(new_n272), .B2(G68), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT71), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n275), .A2(G50), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n393), .B2(new_n394), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n280), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT11), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI211_X1 g0200(.A(KEYINPUT11), .B(new_n280), .C1(new_n395), .C2(new_n397), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n392), .B1(new_n402), .B2(KEYINPUT72), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT72), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n400), .A2(new_n404), .A3(new_n401), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n231), .A2(G1698), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n258), .B(new_n407), .C1(G226), .C2(G1698), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G33), .A2(G97), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n252), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n253), .B1(new_n255), .B2(new_n217), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(new_n413), .A3(KEYINPUT13), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT13), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n410), .B2(new_n412), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n414), .A2(G169), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT14), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n411), .A2(new_n413), .B1(KEYINPUT70), .B2(KEYINPUT13), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT70), .ZN(new_n420));
  NOR4_X1   g0220(.A1(new_n410), .A2(new_n412), .A3(new_n420), .A4(new_n415), .ZN(new_n421));
  OAI21_X1  g0221(.A(G179), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n417), .A2(KEYINPUT14), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n406), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n414), .A2(G200), .A3(new_n416), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT69), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n414), .A2(new_n416), .A3(KEYINPUT69), .A4(G200), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(G190), .B1(new_n419), .B2(new_n421), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n430), .A2(new_n405), .A3(new_n403), .A4(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n253), .B1(new_n255), .B2(new_n223), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n258), .A2(G238), .A3(G1698), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n258), .A2(new_n260), .ZN(new_n435));
  OAI221_X1 g0235(.A(new_n434), .B1(new_n224), .B2(new_n258), .C1(new_n435), .C2(new_n231), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n433), .B1(new_n436), .B2(new_n263), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(G190), .ZN(new_n438));
  NOR4_X1   g0238(.A1(new_n387), .A2(new_n222), .A3(new_n280), .A4(new_n286), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n271), .A2(new_n275), .B1(G20), .B2(G77), .ZN(new_n440));
  XOR2_X1   g0240(.A(KEYINPUT15), .B(G87), .Z(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n274), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n329), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n384), .A2(G77), .ZN(new_n444));
  NOR3_X1   g0244(.A1(new_n439), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n438), .B(new_n445), .C1(new_n268), .C2(new_n437), .ZN(new_n446));
  INV_X1    g0246(.A(new_n437), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n445), .B1(new_n447), .B2(new_n360), .ZN(new_n448));
  INV_X1    g0248(.A(G179), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n437), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n425), .A2(new_n432), .A3(new_n446), .A4(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n290), .ZN(new_n453));
  INV_X1    g0253(.A(new_n265), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(G169), .ZN(new_n455));
  AOI211_X1 g0255(.A(new_n453), .B(new_n455), .C1(new_n449), .C2(new_n454), .ZN(new_n456));
  NOR4_X1   g0256(.A1(new_n304), .A2(new_n380), .A3(new_n452), .A4(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n258), .A2(new_n272), .A3(G87), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT22), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT22), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n258), .A2(new_n460), .A3(new_n272), .A4(G87), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT24), .ZN(new_n463));
  INV_X1    g0263(.A(G116), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n307), .A2(new_n464), .A3(G20), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT23), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n466), .B1(new_n272), .B2(G107), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n224), .A2(KEYINPUT23), .A3(G20), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n462), .A2(new_n463), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n463), .B1(new_n462), .B2(new_n469), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n280), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n282), .A2(G107), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n473), .A2(KEYINPUT88), .ZN(new_n474));
  XNOR2_X1  g0274(.A(KEYINPUT87), .B(KEYINPUT25), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n475), .B1(new_n473), .B2(KEYINPUT88), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  AND2_X1   g0277(.A1(new_n474), .A2(new_n476), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n248), .A2(G33), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n282), .A2(new_n479), .A3(new_n212), .A4(new_n279), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT80), .ZN(new_n481));
  XNOR2_X1  g0281(.A(new_n480), .B(new_n481), .ZN(new_n482));
  AOI211_X1 g0282(.A(new_n477), .B(new_n478), .C1(G107), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n472), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n308), .A2(new_n310), .A3(G257), .A4(G1698), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n308), .A2(new_n310), .A3(G250), .A4(new_n260), .ZN(new_n486));
  INV_X1    g0286(.A(G294), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n485), .B(new_n486), .C1(new_n307), .C2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n263), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT89), .ZN(new_n490));
  XNOR2_X1  g0290(.A(KEYINPUT5), .B(G41), .ZN(new_n491));
  INV_X1    g0291(.A(G45), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n492), .A2(G1), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n491), .A2(new_n493), .B1(new_n213), .B2(new_n251), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n490), .B1(new_n494), .B2(G264), .ZN(new_n495));
  AND2_X1   g0295(.A1(KEYINPUT5), .A2(G41), .ZN(new_n496));
  NOR2_X1   g0296(.A1(KEYINPUT5), .A2(G41), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n493), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AND4_X1   g0298(.A1(new_n490), .A2(new_n498), .A3(G264), .A4(new_n252), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n489), .B1(new_n495), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT90), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n491), .A2(new_n252), .A3(G274), .A4(new_n493), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n498), .A2(new_n252), .ZN(new_n504));
  OAI21_X1  g0304(.A(KEYINPUT89), .B1(new_n504), .B2(new_n225), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n494), .A2(new_n490), .A3(G264), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n507), .A2(KEYINPUT90), .A3(new_n489), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n502), .A2(new_n503), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n268), .ZN(new_n510));
  INV_X1    g0310(.A(new_n503), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n500), .A2(G190), .A3(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n484), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n502), .A2(G179), .A3(new_n503), .A4(new_n508), .ZN(new_n515));
  OAI21_X1  g0315(.A(G169), .B1(new_n500), .B2(new_n511), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n515), .A2(new_n516), .B1(new_n472), .B2(new_n483), .ZN(new_n517));
  OAI21_X1  g0317(.A(KEYINPUT91), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n515), .A2(new_n516), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n484), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT91), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n512), .B1(new_n509), .B2(new_n268), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n520), .B(new_n521), .C1(new_n484), .C2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(G257), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n503), .B1(new_n504), .B2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G33), .A2(G283), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n308), .A2(new_n310), .A3(G250), .A4(G1698), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n308), .A2(new_n310), .A3(G244), .A4(new_n260), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT4), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n527), .B(new_n528), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n530), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT81), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n529), .A2(KEYINPUT81), .A3(new_n530), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n531), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n526), .B1(new_n536), .B2(new_n252), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(G200), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT78), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT6), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT6), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT78), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n540), .B(new_n542), .C1(G97), .C2(new_n224), .ZN(new_n543));
  INV_X1    g0343(.A(G97), .ZN(new_n544));
  OAI21_X1  g0344(.A(KEYINPUT79), .B1(new_n544), .B2(G107), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT79), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n546), .A2(new_n224), .A3(G97), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n543), .A2(new_n548), .ZN(new_n549));
  AOI22_X1  g0349(.A1(KEYINPUT78), .A2(new_n541), .B1(new_n544), .B2(G107), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n550), .A2(new_n540), .A3(new_n545), .A4(new_n547), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n551), .A3(G20), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n275), .A2(G77), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n334), .A2(new_n335), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n312), .B1(new_n258), .B2(G20), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n224), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n280), .B1(new_n554), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n282), .A2(G97), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n559), .B1(new_n482), .B2(G97), .ZN(new_n560));
  OAI211_X1 g0360(.A(G190), .B(new_n526), .C1(new_n536), .C2(new_n252), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n538), .A2(new_n558), .A3(new_n560), .A4(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n482), .A2(new_n441), .ZN(new_n563));
  INV_X1    g0363(.A(new_n441), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n387), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n308), .A2(new_n310), .A3(new_n272), .A4(G68), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT19), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n273), .B2(new_n544), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n272), .B1(new_n409), .B2(new_n567), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n218), .A2(new_n544), .A3(new_n224), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(KEYINPUT82), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT82), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n570), .A2(new_n574), .A3(new_n571), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n569), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT83), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n280), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n570), .A2(new_n574), .A3(new_n571), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n574), .B1(new_n570), .B2(new_n571), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n566), .B(new_n568), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n581), .A2(KEYINPUT83), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n563), .B(new_n565), .C1(new_n578), .C2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n493), .A2(new_n219), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n252), .ZN(new_n585));
  INV_X1    g0385(.A(new_n493), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n585), .B1(new_n352), .B2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n308), .A2(new_n310), .A3(G244), .A4(G1698), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n308), .A2(new_n310), .A3(G238), .A4(new_n260), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n588), .B(new_n589), .C1(new_n307), .C2(new_n464), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n587), .B1(new_n263), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n449), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n263), .ZN(new_n593));
  INV_X1    g0393(.A(new_n352), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n594), .A2(new_n493), .B1(new_n252), .B2(new_n584), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n360), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n583), .A2(new_n592), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n537), .A2(new_n360), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n449), .B(new_n526), .C1(new_n536), .C2(new_n252), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n558), .A2(new_n560), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n593), .A2(new_n266), .A3(new_n595), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(new_n591), .B2(G200), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n581), .A2(KEYINPUT83), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n576), .A2(new_n577), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(new_n606), .A3(new_n280), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n482), .A2(G87), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n604), .A2(new_n607), .A3(new_n565), .A4(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n562), .A2(new_n598), .A3(new_n602), .A4(new_n609), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n527), .B(new_n272), .C1(G33), .C2(new_n544), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT20), .ZN(new_n612));
  AOI22_X1  g0412(.A1(KEYINPUT86), .A2(new_n612), .B1(new_n464), .B2(G20), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n611), .A2(new_n613), .A3(new_n280), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n612), .A2(KEYINPUT86), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n611), .A2(new_n613), .A3(new_n280), .A4(new_n615), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n384), .A2(new_n329), .A3(G116), .A4(new_n479), .ZN(new_n620));
  AOI21_X1  g0420(.A(KEYINPUT85), .B1(new_n387), .B2(new_n464), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT85), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n384), .A2(new_n622), .A3(G116), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n619), .B(new_n620), .C1(new_n621), .C2(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n308), .A2(new_n310), .A3(G264), .A4(G1698), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(KEYINPUT84), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT84), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n258), .A2(new_n627), .A3(G264), .A4(G1698), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n311), .A2(G303), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n258), .A2(G257), .A3(new_n260), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n626), .A2(new_n628), .A3(new_n629), .A4(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n263), .ZN(new_n632));
  INV_X1    g0432(.A(G270), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n503), .B1(new_n504), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n624), .B1(new_n636), .B2(G200), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n634), .B1(new_n631), .B2(new_n263), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(G190), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n636), .A2(new_n624), .A3(G169), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT21), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n624), .A2(new_n638), .A3(G179), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n636), .A2(new_n624), .A3(KEYINPUT21), .A4(G169), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n640), .A2(new_n643), .A3(new_n644), .A4(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n610), .A2(new_n646), .ZN(new_n647));
  AND4_X1   g0447(.A1(new_n457), .A2(new_n518), .A3(new_n523), .A4(new_n647), .ZN(G372));
  INV_X1    g0448(.A(new_n456), .ZN(new_n649));
  INV_X1    g0449(.A(new_n369), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n425), .A2(new_n451), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n651), .A2(new_n432), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n650), .B1(new_n652), .B2(new_n379), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n649), .B1(new_n653), .B2(new_n304), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT92), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n645), .A2(new_n644), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n638), .A2(new_n360), .ZN(new_n657));
  AOI21_X1  g0457(.A(KEYINPUT21), .B1(new_n657), .B2(new_n624), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n655), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n643), .A2(KEYINPUT92), .A3(new_n644), .A4(new_n645), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n520), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n610), .A2(new_n514), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n598), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT26), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n598), .A2(new_n609), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n666), .B1(new_n667), .B2(new_n602), .ZN(new_n668));
  INV_X1    g0468(.A(new_n602), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n669), .A2(KEYINPUT26), .A3(new_n598), .A4(new_n609), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n665), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n664), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n654), .B1(new_n457), .B2(new_n672), .ZN(new_n673));
  XOR2_X1   g0473(.A(new_n673), .B(KEYINPUT93), .Z(G369));
  NAND2_X1  g0474(.A1(new_n390), .A2(new_n272), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G213), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(G343), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n484), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n518), .A2(new_n523), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n517), .A2(new_n680), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g0484(.A(KEYINPUT94), .B(G330), .Z(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n656), .A2(new_n658), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n624), .A2(new_n680), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(new_n640), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n661), .B2(new_n688), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n684), .A2(new_n686), .A3(new_n690), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n691), .A2(KEYINPUT95), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(KEYINPUT95), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n520), .A2(new_n680), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n697));
  INV_X1    g0497(.A(new_n680), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(KEYINPUT96), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(KEYINPUT96), .B1(new_n697), .B2(new_n698), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n696), .B1(new_n684), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n695), .A2(new_n704), .ZN(G399));
  INV_X1    g0505(.A(new_n207), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G41), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n571), .A2(G116), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(G1), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n210), .B2(new_n708), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT29), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n672), .A2(new_n713), .A3(new_n698), .ZN(new_n714));
  INV_X1    g0514(.A(new_n610), .ZN(new_n715));
  INV_X1    g0515(.A(new_n514), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n520), .A2(new_n687), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n680), .B1(new_n671), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n714), .B1(new_n713), .B2(new_n719), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n518), .A2(new_n647), .A3(new_n523), .A4(new_n698), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  INV_X1    g0522(.A(new_n531), .ZN(new_n723));
  AOI21_X1  g0523(.A(KEYINPUT81), .B1(new_n529), .B2(new_n530), .ZN(new_n724));
  INV_X1    g0524(.A(new_n535), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n525), .B1(new_n726), .B2(new_n263), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n727), .A2(new_n502), .A3(new_n508), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n638), .A2(G179), .A3(new_n591), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n722), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n500), .A2(new_n501), .ZN(new_n731));
  AOI21_X1  g0531(.A(KEYINPUT90), .B1(new_n507), .B2(new_n489), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n729), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n733), .A2(KEYINPUT30), .A3(new_n734), .A4(new_n727), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n638), .A2(new_n591), .A3(G179), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n509), .A2(new_n537), .A3(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n730), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(new_n680), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT31), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n738), .A2(KEYINPUT31), .A3(new_n680), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n721), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(new_n685), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n720), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n712), .B1(new_n746), .B2(G1), .ZN(G364));
  NOR2_X1   g0547(.A1(new_n389), .A2(G20), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n248), .B1(new_n748), .B2(G45), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n707), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n751), .B1(new_n690), .B2(new_n686), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(new_n686), .B2(new_n690), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT97), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n258), .A2(new_n207), .ZN(new_n755));
  INV_X1    g0555(.A(G355), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n755), .A2(new_n756), .B1(G116), .B2(new_n207), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n245), .A2(G45), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n706), .A2(new_n258), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n760), .B1(new_n211), .B2(new_n492), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n757), .B1(new_n758), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n212), .B1(G20), .B2(new_n360), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n763), .A2(KEYINPUT98), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(KEYINPUT98), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G13), .A2(G33), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(G20), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n751), .B1(new_n762), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n272), .A2(new_n449), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n773), .A2(G190), .A3(new_n268), .ZN(new_n774));
  INV_X1    g0574(.A(G322), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G190), .A2(G200), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n773), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G311), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n311), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n272), .A2(G179), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(new_n777), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n776), .B(new_n780), .C1(G329), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n773), .A2(G200), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n266), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G326), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n785), .A2(G190), .ZN(new_n788));
  XNOR2_X1  g0588(.A(KEYINPUT33), .B(G317), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n781), .A2(G190), .A3(G200), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n788), .A2(new_n789), .B1(new_n791), .B2(G303), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n266), .A2(G179), .A3(G200), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n272), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n781), .A2(new_n266), .A3(G200), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n795), .A2(G294), .B1(new_n797), .B2(G283), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n784), .A2(new_n787), .A3(new_n792), .A4(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n790), .A2(new_n218), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n783), .A2(G159), .ZN(new_n802));
  INV_X1    g0602(.A(new_n788), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n801), .B1(new_n802), .B2(KEYINPUT32), .C1(new_n803), .C2(new_n216), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n802), .A2(KEYINPUT32), .B1(G107), .B2(new_n797), .ZN(new_n805));
  INV_X1    g0605(.A(new_n786), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n805), .B1(new_n287), .B2(new_n806), .C1(new_n544), .C2(new_n794), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n258), .B1(new_n778), .B2(new_n222), .C1(new_n315), .C2(new_n774), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n799), .B1(new_n804), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n772), .B1(new_n810), .B2(new_n766), .ZN(new_n811));
  INV_X1    g0611(.A(new_n769), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n690), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n754), .A2(new_n813), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n814), .A2(KEYINPUT99), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n814), .A2(KEYINPUT99), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(G396));
  INV_X1    g0618(.A(new_n751), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n672), .A2(new_n698), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT101), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n448), .A2(new_n450), .A3(new_n698), .ZN(new_n822));
  OR2_X1    g0622(.A1(new_n445), .A2(new_n698), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n446), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n451), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n821), .B(new_n822), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n446), .A2(new_n823), .B1(new_n448), .B2(new_n450), .ZN(new_n827));
  INV_X1    g0627(.A(new_n822), .ZN(new_n828));
  OAI21_X1  g0628(.A(KEYINPUT101), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n820), .B(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n745), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n819), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n835), .A2(KEYINPUT102), .B1(new_n834), .B2(new_n833), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(KEYINPUT102), .B2(new_n835), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n766), .A2(new_n767), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n751), .B1(new_n839), .B2(G77), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n796), .A2(new_n218), .B1(new_n782), .B2(new_n779), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(KEYINPUT100), .ZN(new_n842));
  INV_X1    g0642(.A(G283), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n803), .A2(new_n843), .B1(new_n544), .B2(new_n794), .ZN(new_n844));
  INV_X1    g0644(.A(G303), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n806), .A2(new_n845), .B1(new_n790), .B2(new_n224), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n311), .B1(new_n778), .B2(new_n464), .C1(new_n487), .C2(new_n774), .ZN(new_n847));
  OR4_X1    g0647(.A1(new_n842), .A2(new_n844), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n774), .ZN(new_n849));
  INV_X1    g0649(.A(new_n778), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n849), .A2(G143), .B1(new_n850), .B2(G159), .ZN(new_n851));
  INV_X1    g0651(.A(G150), .ZN(new_n852));
  INV_X1    g0652(.A(G137), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n851), .B1(new_n803), .B2(new_n852), .C1(new_n853), .C2(new_n806), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT34), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n796), .A2(new_n216), .ZN(new_n857));
  INV_X1    g0657(.A(G132), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n258), .B1(new_n782), .B2(new_n858), .C1(new_n287), .C2(new_n790), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n857), .B(new_n859), .C1(G58), .C2(new_n795), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n854), .A2(new_n855), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n848), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n840), .B1(new_n863), .B2(new_n766), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n831), .B2(new_n768), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n837), .A2(new_n865), .ZN(G384));
  NOR3_X1   g0666(.A1(new_n212), .A2(new_n272), .A3(new_n464), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n549), .A2(new_n551), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT35), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n869), .B2(new_n868), .ZN(new_n871));
  XOR2_X1   g0671(.A(new_n871), .B(KEYINPUT36), .Z(new_n872));
  AND2_X1   g0672(.A1(new_n201), .A2(G68), .ZN(new_n873));
  NOR3_X1   g0673(.A1(new_n316), .A2(new_n210), .A3(new_n222), .ZN(new_n874));
  OAI211_X1 g0674(.A(G1), .B(new_n389), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n876), .B(KEYINPUT103), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n406), .A2(new_n680), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n425), .A2(new_n432), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n425), .A2(new_n432), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n880), .A2(new_n406), .A3(new_n680), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n830), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n882), .A2(new_n743), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n345), .A2(new_n364), .ZN(new_n884));
  INV_X1    g0684(.A(new_n678), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n216), .B1(new_n555), .B2(new_n556), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n338), .B1(new_n886), .B2(new_n319), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n280), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n888), .B1(new_n327), .B2(new_n322), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n885), .B1(new_n889), .B2(new_n366), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT37), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n367), .A2(new_n373), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n884), .A2(new_n890), .A3(new_n891), .A4(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT104), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n885), .B1(new_n359), .B2(new_n362), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n314), .A2(new_n320), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n329), .B1(new_n896), .B2(new_n338), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n326), .B1(new_n325), .B2(KEYINPUT16), .ZN(new_n898));
  AND4_X1   g0698(.A1(new_n326), .A2(new_n314), .A3(KEYINPUT16), .A4(new_n320), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n895), .B1(new_n900), .B2(new_n344), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n894), .B(KEYINPUT37), .C1(new_n378), .C2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n893), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n900), .A2(new_n344), .ZN(new_n904));
  INV_X1    g0704(.A(new_n895), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n892), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n894), .B1(new_n907), .B2(KEYINPUT37), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT105), .B1(new_n903), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n378), .A2(new_n901), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT104), .B1(new_n910), .B2(new_n891), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT105), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n911), .A2(new_n912), .A3(new_n893), .A4(new_n902), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n909), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n904), .A2(new_n885), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n369), .B2(new_n379), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT38), .B1(new_n914), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT38), .ZN(new_n919));
  AOI211_X1 g0719(.A(new_n919), .B(new_n916), .C1(new_n909), .C2(new_n913), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n883), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT40), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n914), .A2(KEYINPUT38), .A3(new_n917), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n380), .A2(new_n345), .A3(new_n885), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n884), .A2(new_n890), .A3(new_n892), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(KEYINPUT37), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n893), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n919), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n924), .A2(new_n930), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n882), .A2(KEYINPUT40), .A3(new_n743), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n923), .A2(new_n933), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n457), .A2(new_n743), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n686), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(new_n934), .B2(new_n935), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n914), .A2(new_n917), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n919), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n924), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n881), .A2(new_n879), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n672), .A2(new_n831), .A3(new_n698), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n942), .B1(new_n943), .B2(new_n822), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n940), .A2(new_n944), .B1(new_n650), .B2(new_n678), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n939), .A2(KEYINPUT39), .A3(new_n924), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n425), .A2(new_n680), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT39), .ZN(new_n948));
  AOI21_X1  g0748(.A(KEYINPUT38), .B1(new_n925), .B2(new_n928), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n948), .B1(new_n920), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n946), .A2(new_n947), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n945), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n654), .B1(new_n720), .B2(new_n457), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n952), .B(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n937), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n937), .A2(new_n954), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT106), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n955), .B1(new_n248), .B2(new_n748), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n956), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n959), .A2(KEYINPUT106), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n877), .B1(new_n958), .B2(new_n960), .ZN(G367));
  NOR2_X1   g0761(.A1(new_n238), .A2(new_n760), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n771), .B1(new_n706), .B2(new_n441), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(G159), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n803), .A2(new_n965), .B1(new_n201), .B2(new_n778), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT114), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n258), .B1(new_n774), .B2(new_n852), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(G137), .B2(new_n783), .ZN(new_n969));
  AOI22_X1  g0769(.A1(G68), .A2(new_n795), .B1(new_n786), .B2(G143), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n796), .A2(new_n222), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(G58), .B2(new_n791), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n967), .A2(new_n969), .A3(new_n970), .A4(new_n972), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n803), .A2(new_n487), .B1(new_n796), .B2(new_n544), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n806), .A2(new_n779), .B1(new_n224), .B2(new_n794), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n311), .B1(new_n778), .B2(new_n843), .ZN(new_n977));
  INV_X1    g0777(.A(G317), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n774), .A2(new_n845), .B1(new_n782), .B2(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n790), .A2(new_n464), .ZN(new_n980));
  AOI211_X1 g0780(.A(new_n977), .B(new_n979), .C1(KEYINPUT46), .C2(new_n980), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n976), .B(new_n981), .C1(KEYINPUT46), .C2(new_n980), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n973), .A2(KEYINPUT47), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n766), .ZN(new_n984));
  AOI21_X1  g0784(.A(KEYINPUT47), .B1(new_n973), .B2(new_n982), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n751), .B1(new_n962), .B2(new_n964), .C1(new_n984), .C2(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n607), .A2(new_n565), .A3(new_n608), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n987), .A2(new_n680), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n665), .A2(new_n988), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n989), .A2(KEYINPUT107), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n989), .B(KEYINPUT107), .C1(new_n667), .C2(new_n988), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n986), .B1(new_n992), .B2(new_n769), .ZN(new_n993));
  XNOR2_X1  g0793(.A(KEYINPUT111), .B(KEYINPUT45), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n601), .A2(new_n680), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n562), .A2(new_n602), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(KEYINPUT108), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n669), .A2(new_n680), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT108), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n562), .A2(new_n602), .A3(new_n999), .A4(new_n995), .ZN(new_n1000));
  AND3_X1   g0800(.A1(new_n997), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n704), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(KEYINPUT112), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT112), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n704), .A2(new_n1005), .A3(new_n1002), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n994), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1005), .B1(new_n704), .B2(new_n1002), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n702), .B1(new_n682), .B2(new_n683), .ZN(new_n1009));
  NOR4_X1   g0809(.A1(new_n1009), .A2(KEYINPUT112), .A3(new_n1001), .A4(new_n696), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n994), .ZN(new_n1011));
  NOR3_X1   g0811(.A1(new_n1008), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1007), .A2(new_n1012), .ZN(new_n1013));
  OAI211_X1 g0813(.A(KEYINPUT44), .B(new_n1001), .C1(new_n1009), .C2(new_n696), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(KEYINPUT113), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT44), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1001), .B1(new_n1009), .B2(new_n696), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1016), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1019), .A2(KEYINPUT113), .A3(new_n1014), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n694), .B1(new_n1013), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n690), .A2(new_n686), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n684), .B(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1024), .A2(new_n702), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1024), .A2(new_n702), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n746), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1015), .B(new_n1019), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1004), .A2(new_n1006), .A3(new_n994), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1011), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1031), .A2(new_n1034), .A3(new_n695), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1022), .A2(new_n1030), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n746), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n707), .B(KEYINPUT41), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n749), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n695), .A2(new_n1001), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n997), .A2(new_n1000), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n602), .B1(new_n1042), .B2(new_n520), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1009), .A2(new_n1002), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n1043), .A2(new_n698), .B1(new_n1044), .B2(KEYINPUT42), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1044), .A2(KEYINPUT42), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT43), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n992), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n990), .A2(new_n991), .A3(KEYINPUT43), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1047), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1045), .A2(new_n1046), .A3(new_n1048), .A4(new_n992), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1041), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT109), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1053), .B(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1041), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT110), .ZN(new_n1057));
  AND2_X1   g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1059));
  NOR3_X1   g0859(.A1(new_n1055), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n993), .B1(new_n1040), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(G387));
  OAI211_X1 g0862(.A(new_n1026), .B(new_n1027), .C1(new_n745), .C2(new_n720), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1029), .A2(new_n707), .A3(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n682), .A2(new_n683), .A3(new_n769), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n755), .A2(new_n709), .B1(G107), .B2(new_n207), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n234), .A2(new_n492), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n271), .A2(new_n287), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT50), .Z(new_n1069));
  INV_X1    g0869(.A(new_n709), .ZN(new_n1070));
  AOI211_X1 g0870(.A(G45), .B(new_n1070), .C1(G68), .C2(G77), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n760), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1066), .B1(new_n1067), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n751), .B1(new_n1073), .B2(new_n771), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n778), .A2(new_n216), .B1(new_n782), .B2(new_n852), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n311), .B(new_n1075), .C1(G50), .C2(new_n849), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n791), .A2(G77), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n564), .A2(new_n794), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n271), .B2(new_n788), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n786), .A2(G159), .B1(new_n797), .B2(G97), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1076), .A2(new_n1077), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n258), .B1(new_n783), .B2(G326), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n794), .A2(new_n843), .B1(new_n790), .B2(new_n487), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n849), .A2(G317), .B1(new_n850), .B2(G303), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n1084), .B1(new_n803), .B2(new_n779), .C1(new_n775), .C2(new_n806), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT48), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1083), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n1086), .B2(new_n1085), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT49), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1082), .B1(new_n464), .B2(new_n796), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1081), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1074), .B1(new_n1092), .B2(new_n766), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1028), .A2(new_n750), .B1(new_n1065), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1064), .A2(new_n1094), .ZN(G393));
  NAND3_X1  g0895(.A1(new_n1022), .A2(new_n750), .A3(new_n1035), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n766), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n794), .A2(new_n222), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n271), .B2(new_n850), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n201), .B2(new_n803), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT115), .Z(new_n1101));
  OAI22_X1  g0901(.A1(new_n806), .A2(new_n852), .B1(new_n965), .B2(new_n774), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT51), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n796), .A2(new_n218), .ZN(new_n1104));
  INV_X1    g0904(.A(G143), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n258), .B1(new_n782), .B2(new_n1105), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1104), .B(new_n1106), .C1(G68), .C2(new_n791), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1101), .A2(new_n1103), .A3(new_n1107), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(G317), .A2(new_n786), .B1(new_n849), .B2(G311), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT52), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n311), .B1(new_n782), .B2(new_n775), .C1(new_n487), .C2(new_n778), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n803), .A2(new_n845), .B1(new_n796), .B2(new_n224), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n794), .A2(new_n464), .B1(new_n790), .B2(new_n843), .ZN(new_n1113));
  OR4_X1    g0913(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1097), .B1(new_n1108), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n242), .A2(new_n759), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n771), .B1(G97), .B2(new_n706), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n819), .B(new_n1115), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  XOR2_X1   g0918(.A(new_n1118), .B(KEYINPUT116), .Z(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n812), .B2(new_n1002), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n1096), .A2(KEYINPUT117), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(KEYINPUT117), .B1(new_n1096), .B2(new_n1120), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1036), .A2(new_n707), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1031), .A2(new_n1034), .A3(new_n695), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n695), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(KEYINPUT118), .B1(new_n1127), .B2(new_n1030), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1022), .A2(new_n1035), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT118), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1129), .A2(new_n1130), .A3(new_n1029), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1124), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1123), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(G390));
  INV_X1    g0934(.A(G330), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n738), .A2(KEYINPUT31), .A3(new_n680), .ZN(new_n1136));
  AOI21_X1  g0936(.A(KEYINPUT31), .B1(new_n738), .B2(new_n680), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1135), .B1(new_n1138), .B2(new_n721), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n882), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n943), .A2(new_n822), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n947), .B1(new_n1142), .B2(new_n941), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(new_n946), .B2(new_n950), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n828), .B1(new_n719), .B2(new_n831), .ZN(new_n1145));
  OR2_X1    g0945(.A1(new_n1145), .A2(new_n942), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n947), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1146), .A2(new_n1147), .A3(new_n931), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1141), .B1(new_n1144), .B2(new_n1149), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n943), .A2(new_n822), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1147), .B1(new_n1151), .B2(new_n942), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n918), .A2(new_n920), .A3(new_n948), .ZN(new_n1153));
  AOI21_X1  g0953(.A(KEYINPUT39), .B1(new_n924), .B2(new_n930), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1152), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n743), .A2(new_n686), .A3(new_n831), .A4(new_n941), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1155), .A2(new_n1148), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1150), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n767), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n751), .B1(new_n839), .B2(new_n271), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n774), .A2(new_n464), .B1(new_n782), .B2(new_n487), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n258), .B(new_n1162), .C1(G97), .C2(new_n850), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n788), .A2(G107), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1098), .B1(G283), .B2(new_n786), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n800), .A2(new_n857), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(G125), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n258), .B1(new_n782), .B2(new_n1168), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n803), .A2(new_n853), .B1(new_n796), .B2(new_n201), .ZN(new_n1170));
  INV_X1    g0970(.A(G128), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n806), .A2(new_n1171), .B1(new_n965), .B2(new_n794), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT54), .B(G143), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n774), .A2(new_n858), .B1(new_n778), .B2(new_n1173), .ZN(new_n1174));
  OR4_X1    g0974(.A1(new_n1169), .A2(new_n1170), .A3(new_n1172), .A4(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n791), .A2(G150), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT53), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1167), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1161), .B1(new_n1178), .B2(new_n766), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1159), .A2(new_n750), .B1(new_n1160), .B2(new_n1179), .ZN(new_n1180));
  AOI211_X1 g0980(.A(KEYINPUT29), .B(new_n680), .C1(new_n664), .C2(new_n671), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n671), .A2(new_n718), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n713), .B1(new_n1182), .B2(new_n698), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n457), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n652), .A2(new_n379), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n369), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n302), .A2(new_n303), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n295), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n456), .B1(new_n1186), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1139), .A2(new_n457), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1184), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(KEYINPUT119), .ZN(new_n1193));
  AND4_X1   g0993(.A1(new_n518), .A2(new_n647), .A3(new_n523), .A4(new_n698), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n741), .A2(new_n742), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n686), .B(new_n831), .C1(new_n1194), .C2(new_n1195), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n1196), .A2(new_n942), .B1(new_n1139), .B2(new_n882), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1156), .A2(new_n1145), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n941), .B1(new_n1139), .B2(new_n831), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n1197), .A2(new_n1151), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT119), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1184), .A2(new_n1190), .A3(new_n1201), .A4(new_n1191), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1193), .A2(new_n1200), .A3(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1158), .A2(new_n1203), .ZN(new_n1204));
  AND3_X1   g1004(.A1(new_n1193), .A2(new_n1200), .A3(new_n1202), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1150), .A2(new_n1157), .A3(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1204), .A2(new_n707), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1180), .A2(new_n1207), .ZN(G378));
  AOI21_X1  g1008(.A(new_n819), .B1(new_n838), .B2(new_n201), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n796), .A2(new_n315), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1211), .B1(new_n803), .B2(new_n544), .C1(new_n464), .C2(new_n806), .ZN(new_n1212));
  INV_X1    g1012(.A(G41), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1213), .B(new_n311), .C1(new_n782), .C2(new_n843), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n564), .A2(new_n778), .B1(new_n224), .B2(new_n774), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1077), .B1(new_n216), .B2(new_n794), .ZN(new_n1216));
  OR4_X1    g1016(.A1(new_n1212), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT58), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1220));
  AOI21_X1  g1020(.A(G50), .B1(new_n307), .B2(new_n1213), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n258), .B2(G41), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1220), .A2(new_n1222), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n1168), .A2(new_n806), .B1(new_n803), .B2(new_n858), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n849), .A2(G128), .B1(new_n850), .B2(G137), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n790), .B2(new_n1173), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1224), .B(new_n1226), .C1(G150), .C2(new_n795), .ZN(new_n1227));
  XOR2_X1   g1027(.A(new_n1227), .B(KEYINPUT120), .Z(new_n1228));
  OR2_X1    g1028(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1229));
  AOI211_X1 g1029(.A(G33), .B(G41), .C1(new_n783), .C2(G124), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n965), .B2(new_n796), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n1228), .B2(KEYINPUT59), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n1219), .B(new_n1223), .C1(new_n1229), .C2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1209), .B1(new_n1233), .B2(new_n1097), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1189), .B(new_n649), .C1(new_n453), .C2(new_n678), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n290), .B(new_n885), .C1(new_n304), .C2(new_n456), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1237), .B(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1234), .B1(new_n1241), .B2(new_n767), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT40), .B1(new_n940), .B2(new_n883), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n933), .A2(G330), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1241), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1135), .B1(new_n931), .B2(new_n932), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n923), .A2(new_n1240), .A3(new_n1246), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1245), .A2(new_n951), .A3(new_n945), .A4(new_n1247), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n923), .A2(new_n1246), .A3(new_n1240), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1240), .B1(new_n923), .B2(new_n1246), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n952), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1248), .A2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1242), .B1(new_n1252), .B2(new_n750), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n1249), .A2(new_n952), .A3(new_n1250), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n1245), .A2(new_n1247), .B1(new_n951), .B2(new_n945), .ZN(new_n1255));
  OAI21_X1  g1055(.A(KEYINPUT57), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1201), .B1(new_n953), .B2(new_n1191), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1202), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1206), .A2(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n707), .B1(new_n1256), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1206), .A2(new_n1259), .ZN(new_n1262));
  AOI21_X1  g1062(.A(KEYINPUT57), .B1(new_n1262), .B2(new_n1252), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1253), .B1(new_n1261), .B2(new_n1263), .ZN(G375));
  AOI21_X1  g1064(.A(new_n819), .B1(new_n838), .B2(new_n216), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n788), .A2(G116), .B1(new_n786), .B2(G294), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1266), .B1(new_n544), .B2(new_n790), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n258), .B1(new_n783), .B2(G303), .ZN(new_n1268));
  OAI221_X1 g1068(.A(new_n1268), .B1(new_n224), .B2(new_n778), .C1(new_n843), .C2(new_n774), .ZN(new_n1269));
  NOR4_X1   g1069(.A1(new_n1267), .A2(new_n1269), .A3(new_n971), .A4(new_n1078), .ZN(new_n1270));
  OAI221_X1 g1070(.A(new_n258), .B1(new_n782), .B2(new_n1171), .C1(new_n852), .C2(new_n778), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1211), .B1(new_n287), .B2(new_n794), .ZN(new_n1272));
  AOI211_X1 g1072(.A(new_n1271), .B(new_n1272), .C1(G159), .C2(new_n791), .ZN(new_n1273));
  XOR2_X1   g1073(.A(new_n1273), .B(KEYINPUT121), .Z(new_n1274));
  NAND2_X1  g1074(.A1(new_n786), .A2(G132), .ZN(new_n1275));
  OAI221_X1 g1075(.A(new_n1275), .B1(new_n853), .B2(new_n774), .C1(new_n803), .C2(new_n1173), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1270), .B1(new_n1274), .B2(new_n1277), .ZN(new_n1278));
  OAI221_X1 g1078(.A(new_n1265), .B1(new_n1097), .B2(new_n1278), .C1(new_n941), .C2(new_n768), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1200), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1279), .B1(new_n1280), .B2(new_n749), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1203), .A2(new_n1038), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1200), .B1(new_n1193), .B2(new_n1202), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1282), .B1(new_n1283), .B2(new_n1284), .ZN(G381));
  INV_X1    g1085(.A(G375), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(G393), .A2(G396), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  NOR4_X1   g1088(.A1(G378), .A2(new_n1288), .A3(G384), .A4(G381), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1286), .A2(new_n1061), .A3(new_n1289), .A4(new_n1133), .ZN(G407));
  INV_X1    g1090(.A(G378), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n679), .A2(G213), .ZN(new_n1292));
  XOR2_X1   g1092(.A(new_n1292), .B(KEYINPUT122), .Z(new_n1293));
  NAND2_X1  g1093(.A1(new_n1291), .A2(new_n1293), .ZN(new_n1294));
  OAI211_X1 g1094(.A(G407), .B(G213), .C1(G375), .C2(new_n1294), .ZN(G409));
  AOI21_X1  g1095(.A(new_n817), .B1(new_n1064), .B2(new_n1094), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1287), .A2(new_n1296), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1297), .B1(new_n1123), .B2(new_n1132), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1122), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1096), .A2(KEYINPUT117), .A3(new_n1120), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1297), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n708), .B1(new_n1127), .B2(new_n1030), .ZN(new_n1303));
  AOI211_X1 g1103(.A(KEYINPUT118), .B(new_n1030), .C1(new_n1022), .C2(new_n1035), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1130), .B1(new_n1129), .B2(new_n1029), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1303), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1301), .A2(new_n1302), .A3(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1298), .A2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(G387), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1298), .A2(new_n1307), .A3(new_n1061), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT61), .ZN(new_n1312));
  XNOR2_X1  g1112(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1203), .A2(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1280), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(KEYINPUT124), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT124), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1314), .A2(new_n1315), .A3(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n708), .B1(new_n1284), .B2(KEYINPUT60), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1317), .A2(new_n1319), .A3(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(G384), .B1(new_n1321), .B2(new_n1282), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1321), .A2(G384), .A3(new_n1282), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1325), .A2(G2897), .A3(new_n1293), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1323), .A2(KEYINPUT125), .A3(new_n1324), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT125), .ZN(new_n1328));
  AND3_X1   g1128(.A1(new_n1321), .A2(G384), .A3(new_n1282), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1328), .B1(new_n1329), .B2(new_n1322), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1327), .A2(new_n1330), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n679), .A2(G213), .A3(G2897), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1332), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1326), .B1(new_n1331), .B2(new_n1333), .ZN(new_n1334));
  OAI211_X1 g1134(.A(G378), .B(new_n1253), .C1(new_n1261), .C2(new_n1263), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1262), .A2(new_n1252), .A3(new_n1038), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1253), .A2(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1291), .A2(new_n1337), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1293), .B1(new_n1335), .B2(new_n1338), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1312), .B1(new_n1334), .B2(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT62), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1335), .A2(new_n1338), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1342), .A2(new_n1327), .A3(new_n1292), .A4(new_n1330), .ZN(new_n1343));
  AOI211_X1 g1143(.A(new_n1341), .B(new_n1293), .C1(new_n1335), .C2(new_n1338), .ZN(new_n1344));
  AND2_X1   g1144(.A1(new_n1327), .A2(new_n1330), .ZN(new_n1345));
  AOI22_X1  g1145(.A1(new_n1341), .A2(new_n1343), .B1(new_n1344), .B2(new_n1345), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1311), .B1(new_n1340), .B2(new_n1346), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1311), .A2(KEYINPUT61), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1342), .A2(new_n1292), .ZN(new_n1349));
  OAI211_X1 g1149(.A(new_n1349), .B(new_n1326), .C1(new_n1331), .C2(new_n1333), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT63), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1343), .A2(new_n1351), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1345), .A2(KEYINPUT63), .A3(new_n1339), .ZN(new_n1353));
  NAND4_X1  g1153(.A1(new_n1348), .A2(new_n1350), .A3(new_n1352), .A4(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1347), .A2(new_n1354), .ZN(G405));
  NAND2_X1  g1155(.A1(G375), .A2(new_n1291), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1356), .A2(new_n1325), .A3(new_n1335), .ZN(new_n1357));
  INV_X1    g1157(.A(new_n1335), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1262), .A2(new_n1252), .A3(KEYINPUT57), .ZN(new_n1359));
  AOI22_X1  g1159(.A1(new_n1248), .A2(new_n1251), .B1(new_n1206), .B2(new_n1259), .ZN(new_n1360));
  OAI211_X1 g1160(.A(new_n1359), .B(new_n707), .C1(KEYINPUT57), .C2(new_n1360), .ZN(new_n1361));
  AOI21_X1  g1161(.A(G378), .B1(new_n1361), .B2(new_n1253), .ZN(new_n1362));
  NOR2_X1   g1162(.A1(new_n1358), .A2(new_n1362), .ZN(new_n1363));
  OAI211_X1 g1163(.A(KEYINPUT126), .B(new_n1357), .C1(new_n1363), .C2(new_n1331), .ZN(new_n1364));
  INV_X1    g1164(.A(KEYINPUT126), .ZN(new_n1365));
  NAND3_X1  g1165(.A1(new_n1363), .A2(new_n1365), .A3(new_n1325), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1364), .A2(new_n1366), .ZN(new_n1367));
  INV_X1    g1167(.A(KEYINPUT127), .ZN(new_n1368));
  AND3_X1   g1168(.A1(new_n1298), .A2(new_n1307), .A3(new_n1061), .ZN(new_n1369));
  AOI21_X1  g1169(.A(new_n1061), .B1(new_n1298), .B2(new_n1307), .ZN(new_n1370));
  OAI21_X1  g1170(.A(new_n1368), .B1(new_n1369), .B2(new_n1370), .ZN(new_n1371));
  NAND3_X1  g1171(.A1(new_n1309), .A2(KEYINPUT127), .A3(new_n1310), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1371), .A2(new_n1372), .ZN(new_n1373));
  XNOR2_X1  g1173(.A(new_n1367), .B(new_n1373), .ZN(G402));
endmodule


