

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U554 ( .A1(G1384), .A2(G164), .ZN(n682) );
  INV_X1 U555 ( .A(n708), .ZN(n726) );
  XNOR2_X1 U556 ( .A(n707), .B(n706), .ZN(n712) );
  INV_X1 U557 ( .A(KEYINPUT17), .ZN(n524) );
  XOR2_X1 U558 ( .A(n749), .B(KEYINPUT64), .Z(n522) );
  XNOR2_X1 U559 ( .A(KEYINPUT94), .B(KEYINPUT30), .ZN(n716) );
  XNOR2_X1 U560 ( .A(n717), .B(n716), .ZN(n718) );
  INV_X1 U561 ( .A(KEYINPUT29), .ZN(n706) );
  INV_X1 U562 ( .A(KEYINPUT31), .ZN(n722) );
  INV_X1 U563 ( .A(KEYINPUT95), .ZN(n732) );
  NAND2_X1 U564 ( .A1(n882), .A2(G138), .ZN(n527) );
  AND2_X1 U565 ( .A1(n528), .A2(G2104), .ZN(n881) );
  NOR2_X1 U566 ( .A1(G651), .A2(n624), .ZN(n639) );
  INV_X1 U567 ( .A(KEYINPUT86), .ZN(n535) );
  INV_X1 U568 ( .A(G2104), .ZN(n597) );
  AND2_X1 U569 ( .A1(n597), .A2(G126), .ZN(n523) );
  NAND2_X1 U570 ( .A1(n523), .A2(G2105), .ZN(n533) );
  NOR2_X1 U571 ( .A1(G2104), .A2(G2105), .ZN(n525) );
  XNOR2_X2 U572 ( .A(n525), .B(n524), .ZN(n882) );
  AND2_X1 U573 ( .A1(G2104), .A2(G2105), .ZN(n885) );
  NAND2_X1 U574 ( .A1(G114), .A2(n885), .ZN(n526) );
  NAND2_X1 U575 ( .A1(n527), .A2(n526), .ZN(n531) );
  INV_X1 U576 ( .A(G2105), .ZN(n528) );
  NAND2_X1 U577 ( .A1(G102), .A2(n881), .ZN(n529) );
  XNOR2_X1 U578 ( .A(KEYINPUT85), .B(n529), .ZN(n530) );
  NOR2_X1 U579 ( .A1(n531), .A2(n530), .ZN(n532) );
  NAND2_X1 U580 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U581 ( .A(n535), .B(n534), .ZN(G164) );
  INV_X1 U582 ( .A(G651), .ZN(n540) );
  NOR2_X1 U583 ( .A1(G543), .A2(n540), .ZN(n536) );
  XOR2_X1 U584 ( .A(KEYINPUT1), .B(n536), .Z(n634) );
  NAND2_X1 U585 ( .A1(G64), .A2(n634), .ZN(n538) );
  XOR2_X1 U586 ( .A(KEYINPUT0), .B(G543), .Z(n624) );
  NAND2_X1 U587 ( .A1(G52), .A2(n639), .ZN(n537) );
  NAND2_X1 U588 ( .A1(n538), .A2(n537), .ZN(n546) );
  NOR2_X1 U589 ( .A1(G651), .A2(G543), .ZN(n635) );
  NAND2_X1 U590 ( .A1(n635), .A2(G90), .ZN(n539) );
  XOR2_X1 U591 ( .A(KEYINPUT69), .B(n539), .Z(n543) );
  OR2_X1 U592 ( .A1(n540), .A2(n624), .ZN(n541) );
  XOR2_X1 U593 ( .A(KEYINPUT68), .B(n541), .Z(n636) );
  NAND2_X1 U594 ( .A1(G77), .A2(n636), .ZN(n542) );
  NAND2_X1 U595 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U596 ( .A(KEYINPUT9), .B(n544), .Z(n545) );
  NOR2_X1 U597 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U598 ( .A(KEYINPUT70), .B(n547), .ZN(G171) );
  INV_X1 U599 ( .A(G171), .ZN(G301) );
  AND2_X1 U600 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U601 ( .A(G57), .ZN(G237) );
  NAND2_X1 U602 ( .A1(G7), .A2(G661), .ZN(n548) );
  XNOR2_X1 U603 ( .A(n548), .B(KEYINPUT10), .ZN(n549) );
  XNOR2_X1 U604 ( .A(KEYINPUT72), .B(n549), .ZN(G223) );
  INV_X1 U605 ( .A(G223), .ZN(n824) );
  NAND2_X1 U606 ( .A1(n824), .A2(G567), .ZN(n550) );
  XOR2_X1 U607 ( .A(KEYINPUT11), .B(n550), .Z(G234) );
  NAND2_X1 U608 ( .A1(n635), .A2(G81), .ZN(n551) );
  XNOR2_X1 U609 ( .A(n551), .B(KEYINPUT12), .ZN(n553) );
  NAND2_X1 U610 ( .A1(G68), .A2(n636), .ZN(n552) );
  NAND2_X1 U611 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U612 ( .A(KEYINPUT13), .B(n554), .ZN(n560) );
  NAND2_X1 U613 ( .A1(G56), .A2(n634), .ZN(n555) );
  XOR2_X1 U614 ( .A(KEYINPUT14), .B(n555), .Z(n558) );
  NAND2_X1 U615 ( .A1(G43), .A2(n639), .ZN(n556) );
  XNOR2_X1 U616 ( .A(KEYINPUT73), .B(n556), .ZN(n557) );
  NOR2_X1 U617 ( .A1(n558), .A2(n557), .ZN(n559) );
  NAND2_X1 U618 ( .A1(n560), .A2(n559), .ZN(n1021) );
  INV_X1 U619 ( .A(G860), .ZN(n591) );
  OR2_X1 U620 ( .A1(n1021), .A2(n591), .ZN(G153) );
  NAND2_X1 U621 ( .A1(G301), .A2(G868), .ZN(n569) );
  NAND2_X1 U622 ( .A1(G92), .A2(n635), .ZN(n562) );
  NAND2_X1 U623 ( .A1(G79), .A2(n636), .ZN(n561) );
  NAND2_X1 U624 ( .A1(n562), .A2(n561), .ZN(n566) );
  NAND2_X1 U625 ( .A1(G66), .A2(n634), .ZN(n564) );
  NAND2_X1 U626 ( .A1(G54), .A2(n639), .ZN(n563) );
  NAND2_X1 U627 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U628 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U629 ( .A(KEYINPUT15), .B(n567), .Z(n911) );
  INV_X1 U630 ( .A(n911), .ZN(n1013) );
  INV_X1 U631 ( .A(G868), .ZN(n588) );
  NAND2_X1 U632 ( .A1(n1013), .A2(n588), .ZN(n568) );
  NAND2_X1 U633 ( .A1(n569), .A2(n568), .ZN(G284) );
  NAND2_X1 U634 ( .A1(G63), .A2(n634), .ZN(n571) );
  NAND2_X1 U635 ( .A1(G51), .A2(n639), .ZN(n570) );
  NAND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(KEYINPUT6), .B(n572), .ZN(n578) );
  NAND2_X1 U638 ( .A1(n635), .A2(G89), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(KEYINPUT4), .ZN(n575) );
  NAND2_X1 U640 ( .A1(G76), .A2(n636), .ZN(n574) );
  NAND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U642 ( .A(n576), .B(KEYINPUT5), .Z(n577) );
  NOR2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U644 ( .A(KEYINPUT74), .B(n579), .Z(n580) );
  XNOR2_X1 U645 ( .A(KEYINPUT7), .B(n580), .ZN(G168) );
  XOR2_X1 U646 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U647 ( .A1(n634), .A2(G65), .ZN(n582) );
  NAND2_X1 U648 ( .A1(G78), .A2(n636), .ZN(n581) );
  NAND2_X1 U649 ( .A1(n582), .A2(n581), .ZN(n585) );
  NAND2_X1 U650 ( .A1(G91), .A2(n635), .ZN(n583) );
  XNOR2_X1 U651 ( .A(KEYINPUT71), .B(n583), .ZN(n584) );
  NOR2_X1 U652 ( .A1(n585), .A2(n584), .ZN(n587) );
  NAND2_X1 U653 ( .A1(n639), .A2(G53), .ZN(n586) );
  NAND2_X1 U654 ( .A1(n587), .A2(n586), .ZN(G299) );
  NAND2_X1 U655 ( .A1(G868), .A2(G286), .ZN(n590) );
  NAND2_X1 U656 ( .A1(G299), .A2(n588), .ZN(n589) );
  NAND2_X1 U657 ( .A1(n590), .A2(n589), .ZN(G297) );
  NAND2_X1 U658 ( .A1(n591), .A2(G559), .ZN(n592) );
  NAND2_X1 U659 ( .A1(n592), .A2(n911), .ZN(n593) );
  XNOR2_X1 U660 ( .A(n593), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U661 ( .A1(G868), .A2(n1021), .ZN(n596) );
  NAND2_X1 U662 ( .A1(n911), .A2(G868), .ZN(n594) );
  NOR2_X1 U663 ( .A1(G559), .A2(n594), .ZN(n595) );
  NOR2_X1 U664 ( .A1(n596), .A2(n595), .ZN(G282) );
  AND2_X1 U665 ( .A1(n597), .A2(G2105), .ZN(n886) );
  NAND2_X1 U666 ( .A1(G123), .A2(n886), .ZN(n598) );
  XNOR2_X1 U667 ( .A(n598), .B(KEYINPUT18), .ZN(n600) );
  NAND2_X1 U668 ( .A1(n885), .A2(G111), .ZN(n599) );
  NAND2_X1 U669 ( .A1(n600), .A2(n599), .ZN(n604) );
  NAND2_X1 U670 ( .A1(G99), .A2(n881), .ZN(n602) );
  NAND2_X1 U671 ( .A1(G135), .A2(n882), .ZN(n601) );
  NAND2_X1 U672 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U673 ( .A1(n604), .A2(n603), .ZN(n926) );
  XNOR2_X1 U674 ( .A(n926), .B(G2096), .ZN(n606) );
  INV_X1 U675 ( .A(G2100), .ZN(n605) );
  NAND2_X1 U676 ( .A1(n606), .A2(n605), .ZN(G156) );
  NAND2_X1 U677 ( .A1(n639), .A2(G48), .ZN(n613) );
  NAND2_X1 U678 ( .A1(G86), .A2(n635), .ZN(n608) );
  NAND2_X1 U679 ( .A1(G61), .A2(n634), .ZN(n607) );
  NAND2_X1 U680 ( .A1(n608), .A2(n607), .ZN(n611) );
  NAND2_X1 U681 ( .A1(n636), .A2(G73), .ZN(n609) );
  XOR2_X1 U682 ( .A(KEYINPUT2), .B(n609), .Z(n610) );
  NOR2_X1 U683 ( .A1(n611), .A2(n610), .ZN(n612) );
  NAND2_X1 U684 ( .A1(n613), .A2(n612), .ZN(n614) );
  XOR2_X1 U685 ( .A(KEYINPUT79), .B(n614), .Z(G305) );
  NAND2_X1 U686 ( .A1(G88), .A2(n635), .ZN(n616) );
  NAND2_X1 U687 ( .A1(G75), .A2(n636), .ZN(n615) );
  NAND2_X1 U688 ( .A1(n616), .A2(n615), .ZN(n620) );
  NAND2_X1 U689 ( .A1(G62), .A2(n634), .ZN(n618) );
  NAND2_X1 U690 ( .A1(G50), .A2(n639), .ZN(n617) );
  NAND2_X1 U691 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U692 ( .A1(n620), .A2(n619), .ZN(G166) );
  NAND2_X1 U693 ( .A1(G49), .A2(n639), .ZN(n622) );
  NAND2_X1 U694 ( .A1(G74), .A2(G651), .ZN(n621) );
  NAND2_X1 U695 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U696 ( .A1(n634), .A2(n623), .ZN(n626) );
  NAND2_X1 U697 ( .A1(n624), .A2(G87), .ZN(n625) );
  NAND2_X1 U698 ( .A1(n626), .A2(n625), .ZN(G288) );
  NAND2_X1 U699 ( .A1(G60), .A2(n634), .ZN(n628) );
  NAND2_X1 U700 ( .A1(G47), .A2(n639), .ZN(n627) );
  NAND2_X1 U701 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U702 ( .A1(G85), .A2(n635), .ZN(n629) );
  XNOR2_X1 U703 ( .A(KEYINPUT67), .B(n629), .ZN(n630) );
  NOR2_X1 U704 ( .A1(n631), .A2(n630), .ZN(n633) );
  NAND2_X1 U705 ( .A1(G72), .A2(n636), .ZN(n632) );
  NAND2_X1 U706 ( .A1(n633), .A2(n632), .ZN(G290) );
  NAND2_X1 U707 ( .A1(G67), .A2(n634), .ZN(n644) );
  NAND2_X1 U708 ( .A1(G93), .A2(n635), .ZN(n638) );
  NAND2_X1 U709 ( .A1(G80), .A2(n636), .ZN(n637) );
  NAND2_X1 U710 ( .A1(n638), .A2(n637), .ZN(n642) );
  NAND2_X1 U711 ( .A1(G55), .A2(n639), .ZN(n640) );
  XNOR2_X1 U712 ( .A(KEYINPUT77), .B(n640), .ZN(n641) );
  NOR2_X1 U713 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U714 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U715 ( .A(n645), .B(KEYINPUT78), .Z(n832) );
  NOR2_X1 U716 ( .A1(G868), .A2(n832), .ZN(n646) );
  XNOR2_X1 U717 ( .A(n646), .B(KEYINPUT81), .ZN(n657) );
  XOR2_X1 U718 ( .A(KEYINPUT19), .B(KEYINPUT80), .Z(n647) );
  XNOR2_X1 U719 ( .A(G288), .B(n647), .ZN(n648) );
  XNOR2_X1 U720 ( .A(G166), .B(n648), .ZN(n650) );
  INV_X1 U721 ( .A(G299), .ZN(n701) );
  XNOR2_X1 U722 ( .A(G290), .B(n701), .ZN(n649) );
  XNOR2_X1 U723 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U724 ( .A(n832), .B(n651), .ZN(n652) );
  XNOR2_X1 U725 ( .A(G305), .B(n652), .ZN(n909) );
  XNOR2_X1 U726 ( .A(n1021), .B(KEYINPUT75), .ZN(n654) );
  NAND2_X1 U727 ( .A1(n911), .A2(G559), .ZN(n653) );
  XNOR2_X1 U728 ( .A(n654), .B(n653), .ZN(n830) );
  XNOR2_X1 U729 ( .A(n909), .B(n830), .ZN(n655) );
  NAND2_X1 U730 ( .A1(G868), .A2(n655), .ZN(n656) );
  NAND2_X1 U731 ( .A1(n657), .A2(n656), .ZN(G295) );
  NAND2_X1 U732 ( .A1(G2078), .A2(G2084), .ZN(n659) );
  XOR2_X1 U733 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n658) );
  XNOR2_X1 U734 ( .A(n659), .B(n658), .ZN(n660) );
  NAND2_X1 U735 ( .A1(n660), .A2(G2090), .ZN(n661) );
  XOR2_X1 U736 ( .A(KEYINPUT21), .B(n661), .Z(n662) );
  XNOR2_X1 U737 ( .A(KEYINPUT83), .B(n662), .ZN(n663) );
  NAND2_X1 U738 ( .A1(n663), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U739 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U740 ( .A1(G132), .A2(G82), .ZN(n664) );
  XNOR2_X1 U741 ( .A(n664), .B(KEYINPUT22), .ZN(n665) );
  XNOR2_X1 U742 ( .A(n665), .B(KEYINPUT84), .ZN(n666) );
  NOR2_X1 U743 ( .A1(G218), .A2(n666), .ZN(n667) );
  NAND2_X1 U744 ( .A1(G96), .A2(n667), .ZN(n828) );
  NAND2_X1 U745 ( .A1(n828), .A2(G2106), .ZN(n671) );
  NAND2_X1 U746 ( .A1(G69), .A2(G120), .ZN(n668) );
  NOR2_X1 U747 ( .A1(G237), .A2(n668), .ZN(n669) );
  NAND2_X1 U748 ( .A1(G108), .A2(n669), .ZN(n829) );
  NAND2_X1 U749 ( .A1(n829), .A2(G567), .ZN(n670) );
  NAND2_X1 U750 ( .A1(n671), .A2(n670), .ZN(n844) );
  NAND2_X1 U751 ( .A1(G483), .A2(G661), .ZN(n672) );
  NOR2_X1 U752 ( .A1(n844), .A2(n672), .ZN(n827) );
  NAND2_X1 U753 ( .A1(n827), .A2(G36), .ZN(G176) );
  NAND2_X1 U754 ( .A1(G113), .A2(n885), .ZN(n673) );
  XNOR2_X1 U755 ( .A(n673), .B(KEYINPUT66), .ZN(n676) );
  NAND2_X1 U756 ( .A1(G101), .A2(n881), .ZN(n674) );
  XOR2_X1 U757 ( .A(KEYINPUT23), .B(n674), .Z(n675) );
  NAND2_X1 U758 ( .A1(n676), .A2(n675), .ZN(n680) );
  NAND2_X1 U759 ( .A1(G137), .A2(n882), .ZN(n678) );
  NAND2_X1 U760 ( .A1(G125), .A2(n886), .ZN(n677) );
  NAND2_X1 U761 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U762 ( .A1(n680), .A2(n679), .ZN(G160) );
  INV_X1 U763 ( .A(G166), .ZN(G303) );
  XOR2_X1 U764 ( .A(KEYINPUT27), .B(KEYINPUT91), .Z(n684) );
  INV_X1 U765 ( .A(KEYINPUT65), .ZN(n681) );
  XNOR2_X2 U766 ( .A(n682), .B(n681), .ZN(n752) );
  NAND2_X1 U767 ( .A1(G160), .A2(G40), .ZN(n754) );
  NOR2_X4 U768 ( .A1(n752), .A2(n754), .ZN(n708) );
  NAND2_X1 U769 ( .A1(G2072), .A2(n708), .ZN(n683) );
  XNOR2_X1 U770 ( .A(n684), .B(n683), .ZN(n686) );
  INV_X1 U771 ( .A(G1956), .ZN(n981) );
  NOR2_X1 U772 ( .A1(n708), .A2(n981), .ZN(n685) );
  NOR2_X1 U773 ( .A1(n686), .A2(n685), .ZN(n700) );
  NOR2_X1 U774 ( .A1(n701), .A2(n700), .ZN(n687) );
  XOR2_X1 U775 ( .A(n687), .B(KEYINPUT28), .Z(n705) );
  XNOR2_X1 U776 ( .A(G1996), .B(KEYINPUT92), .ZN(n950) );
  NAND2_X1 U777 ( .A1(n950), .A2(n708), .ZN(n688) );
  XNOR2_X1 U778 ( .A(n688), .B(KEYINPUT26), .ZN(n690) );
  NAND2_X1 U779 ( .A1(n726), .A2(G1341), .ZN(n689) );
  NAND2_X1 U780 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U781 ( .A1(n1021), .A2(n691), .ZN(n697) );
  NAND2_X1 U782 ( .A1(n911), .A2(n697), .ZN(n696) );
  AND2_X1 U783 ( .A1(n726), .A2(G1348), .ZN(n692) );
  XNOR2_X1 U784 ( .A(n692), .B(KEYINPUT93), .ZN(n694) );
  NAND2_X1 U785 ( .A1(n708), .A2(G2067), .ZN(n693) );
  NAND2_X1 U786 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U787 ( .A1(n696), .A2(n695), .ZN(n699) );
  OR2_X1 U788 ( .A1(n911), .A2(n697), .ZN(n698) );
  NAND2_X1 U789 ( .A1(n699), .A2(n698), .ZN(n703) );
  NAND2_X1 U790 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U791 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U792 ( .A1(n705), .A2(n704), .ZN(n707) );
  XNOR2_X1 U793 ( .A(KEYINPUT25), .B(G2078), .ZN(n949) );
  NOR2_X1 U794 ( .A1(n726), .A2(n949), .ZN(n710) );
  INV_X1 U795 ( .A(G1961), .ZN(n986) );
  NOR2_X1 U796 ( .A1(n708), .A2(n986), .ZN(n709) );
  NOR2_X1 U797 ( .A1(n710), .A2(n709), .ZN(n719) );
  NAND2_X1 U798 ( .A1(G171), .A2(n719), .ZN(n711) );
  NAND2_X1 U799 ( .A1(n712), .A2(n711), .ZN(n725) );
  INV_X1 U800 ( .A(G8), .ZN(n713) );
  NOR2_X1 U801 ( .A1(n713), .A2(G1966), .ZN(n714) );
  AND2_X1 U802 ( .A1(n726), .A2(n714), .ZN(n739) );
  NOR2_X1 U803 ( .A1(G2084), .A2(n726), .ZN(n736) );
  NOR2_X1 U804 ( .A1(n739), .A2(n736), .ZN(n715) );
  NAND2_X1 U805 ( .A1(G8), .A2(n715), .ZN(n717) );
  NOR2_X1 U806 ( .A1(n718), .A2(G168), .ZN(n721) );
  NOR2_X1 U807 ( .A1(n719), .A2(G171), .ZN(n720) );
  NOR2_X1 U808 ( .A1(n721), .A2(n720), .ZN(n723) );
  XNOR2_X1 U809 ( .A(n723), .B(n722), .ZN(n724) );
  NAND2_X1 U810 ( .A1(n725), .A2(n724), .ZN(n737) );
  NAND2_X1 U811 ( .A1(G286), .A2(n737), .ZN(n731) );
  NAND2_X1 U812 ( .A1(G8), .A2(n726), .ZN(n797) );
  NOR2_X1 U813 ( .A1(G1971), .A2(n797), .ZN(n728) );
  NOR2_X1 U814 ( .A1(G2090), .A2(n726), .ZN(n727) );
  NOR2_X1 U815 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U816 ( .A1(n729), .A2(G303), .ZN(n730) );
  NAND2_X1 U817 ( .A1(n731), .A2(n730), .ZN(n733) );
  XNOR2_X1 U818 ( .A(n733), .B(n732), .ZN(n734) );
  NAND2_X1 U819 ( .A1(n734), .A2(G8), .ZN(n735) );
  XNOR2_X1 U820 ( .A(n735), .B(KEYINPUT32), .ZN(n790) );
  NAND2_X1 U821 ( .A1(G8), .A2(n736), .ZN(n741) );
  INV_X1 U822 ( .A(n737), .ZN(n738) );
  NOR2_X1 U823 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U824 ( .A1(n741), .A2(n740), .ZN(n791) );
  NAND2_X1 U825 ( .A1(G1976), .A2(G288), .ZN(n1009) );
  AND2_X1 U826 ( .A1(n791), .A2(n1009), .ZN(n742) );
  NAND2_X1 U827 ( .A1(n790), .A2(n742), .ZN(n748) );
  INV_X1 U828 ( .A(n1009), .ZN(n745) );
  NOR2_X1 U829 ( .A1(G1976), .A2(G288), .ZN(n1008) );
  NOR2_X1 U830 ( .A1(G1971), .A2(G303), .ZN(n743) );
  NOR2_X1 U831 ( .A1(n1008), .A2(n743), .ZN(n744) );
  OR2_X1 U832 ( .A1(n745), .A2(n744), .ZN(n746) );
  OR2_X1 U833 ( .A1(n797), .A2(n746), .ZN(n747) );
  NAND2_X1 U834 ( .A1(n748), .A2(n747), .ZN(n749) );
  INV_X1 U835 ( .A(KEYINPUT33), .ZN(n750) );
  NAND2_X1 U836 ( .A1(n522), .A2(n750), .ZN(n787) );
  NAND2_X1 U837 ( .A1(n1008), .A2(KEYINPUT33), .ZN(n751) );
  NOR2_X1 U838 ( .A1(n751), .A2(n797), .ZN(n785) );
  XOR2_X1 U839 ( .A(G1981), .B(G305), .Z(n1018) );
  INV_X1 U840 ( .A(n752), .ZN(n753) );
  NOR2_X1 U841 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U842 ( .A(n755), .B(KEYINPUT87), .ZN(n818) );
  XNOR2_X1 U843 ( .A(G1986), .B(G290), .ZN(n1015) );
  NAND2_X1 U844 ( .A1(G107), .A2(n885), .ZN(n757) );
  NAND2_X1 U845 ( .A1(G131), .A2(n882), .ZN(n756) );
  NAND2_X1 U846 ( .A1(n757), .A2(n756), .ZN(n761) );
  NAND2_X1 U847 ( .A1(G95), .A2(n881), .ZN(n759) );
  NAND2_X1 U848 ( .A1(G119), .A2(n886), .ZN(n758) );
  NAND2_X1 U849 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U850 ( .A1(n761), .A2(n760), .ZN(n898) );
  INV_X1 U851 ( .A(G1991), .ZN(n959) );
  NOR2_X1 U852 ( .A1(n898), .A2(n959), .ZN(n770) );
  NAND2_X1 U853 ( .A1(G105), .A2(n881), .ZN(n762) );
  XNOR2_X1 U854 ( .A(n762), .B(KEYINPUT38), .ZN(n764) );
  NAND2_X1 U855 ( .A1(n885), .A2(G117), .ZN(n763) );
  NAND2_X1 U856 ( .A1(n764), .A2(n763), .ZN(n768) );
  NAND2_X1 U857 ( .A1(G141), .A2(n882), .ZN(n766) );
  NAND2_X1 U858 ( .A1(G129), .A2(n886), .ZN(n765) );
  NAND2_X1 U859 ( .A1(n766), .A2(n765), .ZN(n767) );
  OR2_X1 U860 ( .A1(n768), .A2(n767), .ZN(n902) );
  AND2_X1 U861 ( .A1(G1996), .A2(n902), .ZN(n769) );
  NOR2_X1 U862 ( .A1(n770), .A2(n769), .ZN(n808) );
  XNOR2_X1 U863 ( .A(G2067), .B(KEYINPUT37), .ZN(n815) );
  NAND2_X1 U864 ( .A1(n881), .A2(G104), .ZN(n771) );
  XNOR2_X1 U865 ( .A(n771), .B(KEYINPUT88), .ZN(n773) );
  NAND2_X1 U866 ( .A1(G140), .A2(n882), .ZN(n772) );
  NAND2_X1 U867 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U868 ( .A(n774), .B(KEYINPUT89), .ZN(n775) );
  XNOR2_X1 U869 ( .A(n775), .B(KEYINPUT34), .ZN(n781) );
  XNOR2_X1 U870 ( .A(KEYINPUT90), .B(KEYINPUT35), .ZN(n779) );
  NAND2_X1 U871 ( .A1(G116), .A2(n885), .ZN(n777) );
  NAND2_X1 U872 ( .A1(G128), .A2(n886), .ZN(n776) );
  NAND2_X1 U873 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U874 ( .A(n779), .B(n778), .ZN(n780) );
  NAND2_X1 U875 ( .A1(n781), .A2(n780), .ZN(n782) );
  XOR2_X1 U876 ( .A(KEYINPUT36), .B(n782), .Z(n899) );
  OR2_X1 U877 ( .A1(n815), .A2(n899), .ZN(n813) );
  NAND2_X1 U878 ( .A1(n808), .A2(n813), .ZN(n939) );
  NOR2_X1 U879 ( .A1(n1015), .A2(n939), .ZN(n783) );
  OR2_X1 U880 ( .A1(n818), .A2(n783), .ZN(n801) );
  NAND2_X1 U881 ( .A1(n1018), .A2(n801), .ZN(n784) );
  NOR2_X1 U882 ( .A1(n785), .A2(n784), .ZN(n786) );
  NAND2_X1 U883 ( .A1(n787), .A2(n786), .ZN(n803) );
  NOR2_X1 U884 ( .A1(G2090), .A2(G303), .ZN(n788) );
  XNOR2_X1 U885 ( .A(n788), .B(KEYINPUT96), .ZN(n789) );
  NAND2_X1 U886 ( .A1(n789), .A2(G8), .ZN(n793) );
  NAND2_X1 U887 ( .A1(n791), .A2(n790), .ZN(n792) );
  NAND2_X1 U888 ( .A1(n793), .A2(n792), .ZN(n794) );
  NAND2_X1 U889 ( .A1(n794), .A2(n797), .ZN(n799) );
  NOR2_X1 U890 ( .A1(G1981), .A2(G305), .ZN(n795) );
  XOR2_X1 U891 ( .A(n795), .B(KEYINPUT24), .Z(n796) );
  OR2_X1 U892 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U893 ( .A1(n799), .A2(n798), .ZN(n800) );
  NAND2_X1 U894 ( .A1(n801), .A2(n800), .ZN(n802) );
  NAND2_X1 U895 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U896 ( .A(n804), .B(KEYINPUT97), .ZN(n822) );
  NOR2_X1 U897 ( .A1(n902), .A2(G1996), .ZN(n805) );
  XNOR2_X1 U898 ( .A(n805), .B(KEYINPUT98), .ZN(n932) );
  AND2_X1 U899 ( .A1(n959), .A2(n898), .ZN(n927) );
  NOR2_X1 U900 ( .A1(G1986), .A2(G290), .ZN(n806) );
  XOR2_X1 U901 ( .A(n806), .B(KEYINPUT99), .Z(n807) );
  NOR2_X1 U902 ( .A1(n927), .A2(n807), .ZN(n810) );
  INV_X1 U903 ( .A(n808), .ZN(n809) );
  NOR2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U905 ( .A1(n932), .A2(n811), .ZN(n812) );
  XNOR2_X1 U906 ( .A(n812), .B(KEYINPUT39), .ZN(n814) );
  NAND2_X1 U907 ( .A1(n814), .A2(n813), .ZN(n816) );
  NAND2_X1 U908 ( .A1(n815), .A2(n899), .ZN(n936) );
  NAND2_X1 U909 ( .A1(n816), .A2(n936), .ZN(n817) );
  XNOR2_X1 U910 ( .A(KEYINPUT100), .B(n817), .ZN(n820) );
  INV_X1 U911 ( .A(n818), .ZN(n819) );
  NAND2_X1 U912 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U913 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U914 ( .A(n823), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U915 ( .A1(G2106), .A2(n824), .ZN(G217) );
  AND2_X1 U916 ( .A1(G15), .A2(G2), .ZN(n825) );
  NAND2_X1 U917 ( .A1(G661), .A2(n825), .ZN(G259) );
  NAND2_X1 U918 ( .A1(G3), .A2(G1), .ZN(n826) );
  NAND2_X1 U919 ( .A1(n827), .A2(n826), .ZN(G188) );
  NOR2_X1 U920 ( .A1(n829), .A2(n828), .ZN(G325) );
  XOR2_X1 U921 ( .A(KEYINPUT102), .B(G325), .Z(G261) );
  XOR2_X1 U923 ( .A(n830), .B(KEYINPUT76), .Z(n831) );
  NOR2_X1 U924 ( .A1(G860), .A2(n831), .ZN(n833) );
  XNOR2_X1 U925 ( .A(n833), .B(n832), .ZN(G145) );
  INV_X1 U926 ( .A(G132), .ZN(G219) );
  INV_X1 U927 ( .A(G120), .ZN(G236) );
  INV_X1 U928 ( .A(G82), .ZN(G220) );
  INV_X1 U929 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U930 ( .A(G1348), .B(G2435), .ZN(n834) );
  XNOR2_X1 U931 ( .A(n834), .B(G2438), .ZN(n835) );
  XNOR2_X1 U932 ( .A(n835), .B(G1341), .ZN(n841) );
  XOR2_X1 U933 ( .A(G2451), .B(G2446), .Z(n837) );
  XNOR2_X1 U934 ( .A(G2427), .B(G2443), .ZN(n836) );
  XNOR2_X1 U935 ( .A(n837), .B(n836), .ZN(n839) );
  XOR2_X1 U936 ( .A(G2430), .B(G2454), .Z(n838) );
  XNOR2_X1 U937 ( .A(n839), .B(n838), .ZN(n840) );
  XNOR2_X1 U938 ( .A(n841), .B(n840), .ZN(n842) );
  NAND2_X1 U939 ( .A1(n842), .A2(G14), .ZN(n843) );
  XNOR2_X1 U940 ( .A(KEYINPUT101), .B(n843), .ZN(G401) );
  INV_X1 U941 ( .A(n844), .ZN(G319) );
  XOR2_X1 U942 ( .A(G2678), .B(KEYINPUT42), .Z(n846) );
  XNOR2_X1 U943 ( .A(KEYINPUT104), .B(KEYINPUT43), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U945 ( .A(KEYINPUT103), .B(G2090), .Z(n848) );
  XNOR2_X1 U946 ( .A(G2067), .B(G2072), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U948 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U949 ( .A(G2096), .B(G2100), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n852), .B(n851), .ZN(n854) );
  XOR2_X1 U951 ( .A(G2078), .B(G2084), .Z(n853) );
  XNOR2_X1 U952 ( .A(n854), .B(n853), .ZN(G227) );
  XOR2_X1 U953 ( .A(G1976), .B(G1971), .Z(n856) );
  XNOR2_X1 U954 ( .A(G1986), .B(G1961), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U956 ( .A(n857), .B(G2474), .Z(n859) );
  XNOR2_X1 U957 ( .A(G1966), .B(G1981), .ZN(n858) );
  XNOR2_X1 U958 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U959 ( .A(KEYINPUT41), .B(G1956), .Z(n861) );
  XNOR2_X1 U960 ( .A(G1996), .B(G1991), .ZN(n860) );
  XNOR2_X1 U961 ( .A(n861), .B(n860), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n863), .B(n862), .ZN(G229) );
  NAND2_X1 U963 ( .A1(G124), .A2(n886), .ZN(n864) );
  XNOR2_X1 U964 ( .A(n864), .B(KEYINPUT44), .ZN(n866) );
  NAND2_X1 U965 ( .A1(n885), .A2(G112), .ZN(n865) );
  NAND2_X1 U966 ( .A1(n866), .A2(n865), .ZN(n870) );
  NAND2_X1 U967 ( .A1(G100), .A2(n881), .ZN(n868) );
  NAND2_X1 U968 ( .A1(G136), .A2(n882), .ZN(n867) );
  NAND2_X1 U969 ( .A1(n868), .A2(n867), .ZN(n869) );
  NOR2_X1 U970 ( .A1(n870), .A2(n869), .ZN(G162) );
  XNOR2_X1 U971 ( .A(G162), .B(n926), .ZN(n880) );
  NAND2_X1 U972 ( .A1(G118), .A2(n885), .ZN(n872) );
  NAND2_X1 U973 ( .A1(G130), .A2(n886), .ZN(n871) );
  NAND2_X1 U974 ( .A1(n872), .A2(n871), .ZN(n878) );
  NAND2_X1 U975 ( .A1(n881), .A2(G106), .ZN(n873) );
  XOR2_X1 U976 ( .A(KEYINPUT105), .B(n873), .Z(n875) );
  NAND2_X1 U977 ( .A1(n882), .A2(G142), .ZN(n874) );
  NAND2_X1 U978 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U979 ( .A(KEYINPUT45), .B(n876), .Z(n877) );
  NOR2_X1 U980 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U981 ( .A(n880), .B(n879), .ZN(n897) );
  XOR2_X1 U982 ( .A(KEYINPUT108), .B(KEYINPUT46), .Z(n895) );
  NAND2_X1 U983 ( .A1(G103), .A2(n881), .ZN(n884) );
  NAND2_X1 U984 ( .A1(G139), .A2(n882), .ZN(n883) );
  NAND2_X1 U985 ( .A1(n884), .A2(n883), .ZN(n892) );
  NAND2_X1 U986 ( .A1(G115), .A2(n885), .ZN(n888) );
  NAND2_X1 U987 ( .A1(G127), .A2(n886), .ZN(n887) );
  NAND2_X1 U988 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U989 ( .A(KEYINPUT47), .B(n889), .Z(n890) );
  XNOR2_X1 U990 ( .A(KEYINPUT106), .B(n890), .ZN(n891) );
  NOR2_X1 U991 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U992 ( .A(KEYINPUT107), .B(n893), .Z(n922) );
  XNOR2_X1 U993 ( .A(n922), .B(KEYINPUT48), .ZN(n894) );
  XNOR2_X1 U994 ( .A(n895), .B(n894), .ZN(n896) );
  XOR2_X1 U995 ( .A(n897), .B(n896), .Z(n901) );
  XOR2_X1 U996 ( .A(n899), .B(n898), .Z(n900) );
  XNOR2_X1 U997 ( .A(n901), .B(n900), .ZN(n905) );
  XOR2_X1 U998 ( .A(G160), .B(n902), .Z(n903) );
  XNOR2_X1 U999 ( .A(G164), .B(n903), .ZN(n904) );
  XOR2_X1 U1000 ( .A(n905), .B(n904), .Z(n906) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n906), .ZN(G395) );
  XNOR2_X1 U1002 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n908) );
  XNOR2_X1 U1003 ( .A(n1021), .B(KEYINPUT109), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(n908), .B(n907), .ZN(n910) );
  XOR2_X1 U1005 ( .A(n910), .B(n909), .Z(n913) );
  XNOR2_X1 U1006 ( .A(G301), .B(n911), .ZN(n912) );
  XNOR2_X1 U1007 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1008 ( .A(n914), .B(G286), .ZN(n915) );
  NOR2_X1 U1009 ( .A1(G37), .A2(n915), .ZN(G397) );
  NOR2_X1 U1010 ( .A1(G227), .A2(G229), .ZN(n916) );
  XOR2_X1 U1011 ( .A(KEYINPUT49), .B(n916), .Z(n917) );
  NAND2_X1 U1012 ( .A1(G319), .A2(n917), .ZN(n918) );
  NOR2_X1 U1013 ( .A1(G401), .A2(n918), .ZN(n919) );
  XNOR2_X1 U1014 ( .A(KEYINPUT112), .B(n919), .ZN(n921) );
  NOR2_X1 U1015 ( .A1(G395), .A2(G397), .ZN(n920) );
  NAND2_X1 U1016 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1017 ( .A(G225), .ZN(G308) );
  INV_X1 U1018 ( .A(G96), .ZN(G221) );
  INV_X1 U1019 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1020 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n945) );
  XOR2_X1 U1021 ( .A(G2072), .B(n922), .Z(n924) );
  XOR2_X1 U1022 ( .A(G164), .B(G2078), .Z(n923) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  XOR2_X1 U1024 ( .A(KEYINPUT50), .B(n925), .Z(n942) );
  XNOR2_X1 U1025 ( .A(G160), .B(G2084), .ZN(n930) );
  NOR2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1027 ( .A(KEYINPUT113), .B(n928), .Z(n929) );
  NAND2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n935) );
  XOR2_X1 U1029 ( .A(G2090), .B(G162), .Z(n931) );
  NOR2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1031 ( .A(n933), .B(KEYINPUT51), .ZN(n934) );
  NOR2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n937) );
  NAND2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1035 ( .A(KEYINPUT114), .B(n940), .Z(n941) );
  NOR2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1037 ( .A(n943), .B(KEYINPUT52), .ZN(n944) );
  XNOR2_X1 U1038 ( .A(n945), .B(n944), .ZN(n947) );
  INV_X1 U1039 ( .A(KEYINPUT55), .ZN(n946) );
  NAND2_X1 U1040 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1041 ( .A1(n948), .A2(G29), .ZN(n1004) );
  XOR2_X1 U1042 ( .A(G2090), .B(G35), .Z(n966) );
  XNOR2_X1 U1043 ( .A(G27), .B(n949), .ZN(n958) );
  XNOR2_X1 U1044 ( .A(n950), .B(G32), .ZN(n956) );
  XOR2_X1 U1045 ( .A(G2072), .B(G33), .Z(n953) );
  XNOR2_X1 U1046 ( .A(G2067), .B(KEYINPUT117), .ZN(n951) );
  XNOR2_X1 U1047 ( .A(n951), .B(G26), .ZN(n952) );
  NAND2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1049 ( .A(n954), .B(KEYINPUT118), .ZN(n955) );
  NOR2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1051 ( .A1(n958), .A2(n957), .ZN(n962) );
  XNOR2_X1 U1052 ( .A(G25), .B(n959), .ZN(n960) );
  NAND2_X1 U1053 ( .A1(n960), .A2(G28), .ZN(n961) );
  NOR2_X1 U1054 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1055 ( .A(n963), .B(KEYINPUT119), .ZN(n964) );
  XNOR2_X1 U1056 ( .A(n964), .B(KEYINPUT53), .ZN(n965) );
  NAND2_X1 U1057 ( .A1(n966), .A2(n965), .ZN(n969) );
  XNOR2_X1 U1058 ( .A(G34), .B(G2084), .ZN(n967) );
  XNOR2_X1 U1059 ( .A(KEYINPUT54), .B(n967), .ZN(n968) );
  NOR2_X1 U1060 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1061 ( .A(KEYINPUT55), .B(n970), .ZN(n972) );
  INV_X1 U1062 ( .A(G29), .ZN(n971) );
  NAND2_X1 U1063 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1064 ( .A1(n973), .A2(G11), .ZN(n974) );
  XNOR2_X1 U1065 ( .A(n974), .B(KEYINPUT120), .ZN(n1002) );
  XOR2_X1 U1066 ( .A(KEYINPUT125), .B(G4), .Z(n976) );
  XNOR2_X1 U1067 ( .A(G1348), .B(KEYINPUT59), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(n976), .B(n975), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(G1341), .B(G19), .ZN(n978) );
  XNOR2_X1 U1070 ( .A(G1981), .B(G6), .ZN(n977) );
  NOR2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n984) );
  XOR2_X1 U1073 ( .A(G20), .B(n981), .Z(n982) );
  XNOR2_X1 U1074 ( .A(KEYINPUT124), .B(n982), .ZN(n983) );
  NOR2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1076 ( .A(KEYINPUT60), .B(n985), .ZN(n988) );
  XNOR2_X1 U1077 ( .A(n986), .B(G5), .ZN(n987) );
  NAND2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n995) );
  XNOR2_X1 U1079 ( .A(G1971), .B(G22), .ZN(n990) );
  XNOR2_X1 U1080 ( .A(G23), .B(G1976), .ZN(n989) );
  NOR2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n992) );
  XOR2_X1 U1082 ( .A(G1986), .B(G24), .Z(n991) );
  NAND2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(KEYINPUT58), .B(n993), .ZN(n994) );
  NOR2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n998) );
  XOR2_X1 U1086 ( .A(G1966), .B(G21), .Z(n996) );
  XNOR2_X1 U1087 ( .A(KEYINPUT126), .B(n996), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1089 ( .A(KEYINPUT61), .B(n999), .ZN(n1000) );
  NOR2_X1 U1090 ( .A1(n1000), .A2(G16), .ZN(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1032) );
  XNOR2_X1 U1093 ( .A(G16), .B(KEYINPUT121), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(n1005), .B(KEYINPUT56), .ZN(n1030) );
  XNOR2_X1 U1095 ( .A(G1971), .B(KEYINPUT122), .ZN(n1006) );
  XNOR2_X1 U1096 ( .A(n1006), .B(G303), .ZN(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1010) );
  NAND2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(G1956), .B(G299), .ZN(n1011) );
  NOR2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1017) );
  XNOR2_X1 U1101 ( .A(G1348), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1027) );
  XNOR2_X1 U1104 ( .A(G1966), .B(G168), .ZN(n1019) );
  NAND2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1106 ( .A(KEYINPUT57), .B(n1020), .ZN(n1025) );
  XNOR2_X1 U1107 ( .A(n1021), .B(G1341), .ZN(n1023) );
  XNOR2_X1 U1108 ( .A(G301), .B(G1961), .ZN(n1022) );
  NOR2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1111 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XOR2_X1 U1112 ( .A(KEYINPUT123), .B(n1028), .Z(n1029) );
  NOR2_X1 U1113 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NOR2_X1 U1114 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1115 ( .A(n1033), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1116 ( .A(G311), .ZN(G150) );
endmodule

