//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 1 1 0 1 0 1 1 1 1 0 0 0 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1281,
    new_n1282;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G58), .ZN(new_n211));
  INV_X1    g0011(.A(G232), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n209), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT1), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n209), .A2(G13), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n221), .B(G250), .C1(G257), .C2(G264), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT0), .Z(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(KEYINPUT64), .ZN(new_n225));
  INV_X1    g0025(.A(KEYINPUT64), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n226), .A2(G1), .A3(G13), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n228), .A2(new_n207), .ZN(new_n229));
  OAI21_X1  g0029(.A(G50), .B1(G58), .B2(G68), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n220), .B(new_n223), .C1(new_n229), .C2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n234), .B(new_n235), .Z(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT65), .B(KEYINPUT66), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n236), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XOR2_X1   g0045(.A(new_n245), .B(KEYINPUT67), .Z(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(KEYINPUT9), .ZN(new_n251));
  XOR2_X1   g0051(.A(KEYINPUT8), .B(G58), .Z(new_n252));
  NAND2_X1  g0052(.A1(new_n207), .A2(G33), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  AOI22_X1  g0055(.A1(new_n252), .A2(new_n254), .B1(G150), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n203), .A2(G20), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n228), .B1(new_n209), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n207), .A2(G1), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G13), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n202), .ZN(new_n265));
  AOI22_X1  g0065(.A1(G33), .A2(new_n208), .B1(new_n225), .B2(new_n227), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(G1), .B2(new_n207), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n261), .B(new_n265), .C1(new_n202), .C2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n269));
  INV_X1    g0069(.A(G274), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G41), .ZN(new_n273));
  OAI211_X1 g0073(.A(G1), .B(G13), .C1(new_n259), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n269), .ZN(new_n275));
  INV_X1    g0075(.A(G226), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n272), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT3), .B(G33), .ZN(new_n278));
  INV_X1    g0078(.A(G1698), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n278), .A2(G222), .A3(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G77), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n278), .A2(G1698), .ZN(new_n282));
  INV_X1    g0082(.A(G223), .ZN(new_n283));
  OAI221_X1 g0083(.A(new_n280), .B1(new_n281), .B2(new_n278), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n277), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n251), .A2(new_n268), .B1(new_n287), .B2(G200), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n265), .B1(new_n267), .B2(new_n202), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n289), .B1(new_n260), .B2(new_n258), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n290), .A2(KEYINPUT9), .B1(G190), .B2(new_n286), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT10), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT10), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n288), .A2(new_n291), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n268), .B1(new_n286), .B2(G169), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT68), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G179), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n286), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n297), .A2(new_n298), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n299), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT3), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G107), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n278), .A2(new_n279), .ZN(new_n309));
  OAI221_X1 g0109(.A(new_n308), .B1(new_n309), .B2(new_n212), .C1(new_n214), .C2(new_n282), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n285), .ZN(new_n311));
  INV_X1    g0111(.A(new_n275), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n271), .B1(new_n312), .B2(G244), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G169), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n264), .A2(new_n281), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(new_n267), .B2(new_n281), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n252), .A2(new_n255), .B1(G20), .B2(G77), .ZN(new_n319));
  XOR2_X1   g0119(.A(KEYINPUT15), .B(G87), .Z(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n254), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n266), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n316), .B(new_n324), .C1(G179), .C2(new_n314), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n314), .A2(G200), .ZN(new_n326));
  INV_X1    g0126(.A(G190), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n326), .B(new_n323), .C1(new_n327), .C2(new_n314), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  AND3_X1   g0129(.A1(new_n296), .A2(new_n303), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT13), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n304), .A2(new_n306), .A3(G226), .A4(new_n279), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT69), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT69), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n278), .A2(new_n334), .A3(G226), .A4(new_n279), .ZN(new_n335));
  INV_X1    g0135(.A(G97), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n259), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n278), .A2(G232), .A3(G1698), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n333), .A2(new_n335), .A3(new_n338), .A4(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n285), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n272), .B1(new_n275), .B2(new_n214), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n331), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  AOI211_X1 g0144(.A(KEYINPUT13), .B(new_n342), .C1(new_n340), .C2(new_n285), .ZN(new_n345));
  OAI21_X1  g0145(.A(G169), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT14), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n344), .A2(new_n345), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(G179), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT14), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n350), .B(G169), .C1(new_n344), .C2(new_n345), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n347), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n264), .A2(new_n213), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n353), .A2(KEYINPUT12), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT71), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT70), .ZN(new_n356));
  OR2_X1    g0156(.A1(new_n356), .A2(KEYINPUT12), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(KEYINPUT12), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n353), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n354), .B1(new_n355), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(new_n355), .B2(new_n359), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n260), .A2(new_n262), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G68), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n255), .A2(G50), .ZN(new_n364));
  OAI221_X1 g0164(.A(new_n364), .B1(new_n207), .B2(G68), .C1(new_n281), .C2(new_n253), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n260), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n366), .B(KEYINPUT11), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n361), .A2(new_n363), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n352), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n368), .ZN(new_n370));
  OAI21_X1  g0170(.A(G200), .B1(new_n344), .B2(new_n345), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n348), .A2(G190), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT18), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n278), .B2(G20), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n305), .A2(G33), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n380));
  OAI211_X1 g0180(.A(KEYINPUT7), .B(new_n207), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n213), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  AND2_X1   g0182(.A1(G58), .A2(G68), .ZN(new_n383));
  OAI21_X1  g0183(.A(G20), .B1(new_n383), .B2(new_n201), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT72), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI211_X1 g0186(.A(KEYINPUT72), .B(G20), .C1(new_n383), .C2(new_n201), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n255), .A2(G159), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NOR3_X1   g0189(.A1(new_n382), .A2(new_n389), .A3(KEYINPUT16), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n386), .A2(KEYINPUT73), .A3(new_n387), .A4(new_n388), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NOR3_X1   g0193(.A1(new_n278), .A2(new_n377), .A3(G20), .ZN(new_n394));
  AOI21_X1  g0194(.A(KEYINPUT7), .B1(new_n307), .B2(new_n207), .ZN(new_n395));
  OAI21_X1  g0195(.A(G68), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AND3_X1   g0196(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT16), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(KEYINPUT16), .B1(new_n382), .B2(new_n389), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n266), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NOR3_X1   g0201(.A1(new_n396), .A2(new_n391), .A3(new_n266), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n393), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n264), .A2(new_n252), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n404), .B1(new_n267), .B2(new_n252), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n278), .A2(G226), .A3(G1698), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G33), .A2(G87), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n408), .B(new_n409), .C1(new_n309), .C2(new_n283), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n285), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n271), .B1(new_n312), .B2(G232), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n315), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n411), .A2(new_n412), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n413), .B1(G179), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n376), .B1(new_n407), .B2(new_n416), .ZN(new_n417));
  AOI211_X1 g0217(.A(KEYINPUT18), .B(new_n415), .C1(new_n403), .C2(new_n406), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(G200), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n420), .B1(new_n411), .B2(new_n412), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n421), .B1(G190), .B2(new_n414), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n403), .A2(new_n406), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT17), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT17), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n403), .A2(new_n425), .A3(new_n406), .A4(new_n422), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n330), .A2(new_n375), .A3(new_n419), .A4(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT74), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n428), .B(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n278), .A2(G250), .A3(new_n279), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n304), .A2(new_n306), .A3(G257), .A4(G1698), .ZN(new_n433));
  NAND2_X1  g0233(.A1(G33), .A2(G294), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n285), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n206), .B(G45), .C1(new_n273), .C2(KEYINPUT5), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n273), .A2(KEYINPUT5), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n224), .B1(G33), .B2(G41), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(G264), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n439), .A2(G274), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n436), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(G169), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT83), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT83), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n444), .A2(new_n447), .A3(G169), .ZN(new_n448));
  INV_X1    g0248(.A(new_n444), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(G179), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n446), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n304), .A2(new_n306), .A3(new_n207), .A4(G87), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT22), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT22), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n278), .A2(new_n454), .A3(new_n207), .A4(G87), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G33), .A2(G116), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(G20), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT23), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n459), .B1(new_n207), .B2(G107), .ZN(new_n460));
  INV_X1    g0260(.A(G107), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n461), .A2(KEYINPUT23), .A3(G20), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n458), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n456), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT24), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT81), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT24), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n456), .A2(new_n466), .A3(new_n467), .A4(new_n463), .ZN(new_n468));
  AND2_X1   g0268(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT81), .B1(new_n464), .B2(KEYINPUT24), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n266), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n264), .A2(new_n461), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT82), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n472), .A2(new_n473), .A3(KEYINPUT25), .ZN(new_n474));
  XOR2_X1   g0274(.A(KEYINPUT82), .B(KEYINPUT25), .Z(new_n475));
  AOI22_X1  g0275(.A1(new_n262), .A2(G13), .B1(new_n206), .B2(G33), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n266), .A2(new_n476), .ZN(new_n477));
  OAI221_X1 g0277(.A(new_n474), .B1(new_n472), .B2(new_n475), .C1(new_n477), .C2(new_n461), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n451), .B1(new_n471), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n278), .A2(new_n207), .A3(G68), .ZN(new_n480));
  XNOR2_X1  g0280(.A(KEYINPUT78), .B(KEYINPUT19), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n253), .A2(new_n336), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NOR3_X1   g0283(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n481), .A2(new_n337), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n484), .B1(new_n485), .B2(new_n207), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n260), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n320), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n264), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n266), .A2(G87), .A3(new_n476), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n487), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n206), .A2(G45), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G250), .ZN(new_n494));
  OAI22_X1  g0294(.A1(new_n440), .A2(new_n494), .B1(new_n270), .B2(new_n493), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n278), .A2(G238), .A3(new_n279), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n278), .A2(G244), .A3(G1698), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n496), .A2(new_n497), .A3(new_n457), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n495), .B1(new_n498), .B2(new_n285), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G200), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n498), .A2(new_n285), .ZN(new_n502));
  INV_X1    g0302(.A(new_n495), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n502), .A2(G190), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT79), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n499), .A2(KEYINPUT79), .A3(G190), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n492), .A2(new_n501), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n487), .B(new_n489), .C1(new_n488), .C2(new_n477), .ZN(new_n509));
  AOI211_X1 g0309(.A(G179), .B(new_n495), .C1(new_n498), .C2(new_n285), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n509), .B(new_n511), .C1(G169), .C2(new_n499), .ZN(new_n512));
  AND2_X1   g0312(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n444), .A2(new_n327), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n514), .B1(G200), .B2(new_n444), .ZN(new_n515));
  INV_X1    g0315(.A(new_n470), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n465), .A2(new_n468), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n260), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n478), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n515), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n479), .A2(new_n513), .A3(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT21), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n266), .A2(G116), .A3(new_n476), .ZN(new_n523));
  INV_X1    g0323(.A(G116), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n264), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT20), .ZN(new_n528));
  AOI21_X1  g0328(.A(G20), .B1(G33), .B2(G283), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n259), .A2(G97), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n529), .A2(new_n530), .B1(G20), .B2(new_n524), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n528), .B1(new_n532), .B2(new_n266), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n260), .A2(KEYINPUT20), .A3(new_n531), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n527), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G169), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n441), .A2(G270), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n443), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n278), .A2(G257), .A3(new_n279), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n307), .A2(G303), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n304), .A2(new_n306), .A3(G264), .A4(G1698), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n285), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT80), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n543), .A2(KEYINPUT80), .A3(new_n285), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n539), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n522), .B1(new_n537), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n548), .A2(G179), .A3(new_n536), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n441), .A2(G270), .B1(G274), .B2(new_n439), .ZN(new_n551));
  INV_X1    g0351(.A(new_n547), .ZN(new_n552));
  AOI21_X1  g0352(.A(KEYINPUT80), .B1(new_n543), .B2(new_n285), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n315), .B1(new_n527), .B2(new_n535), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n554), .A2(new_n555), .A3(KEYINPUT21), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n549), .A2(new_n550), .A3(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n551), .B(G190), .C1(new_n552), .C2(new_n553), .ZN(new_n558));
  INV_X1    g0358(.A(new_n536), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n558), .B(new_n559), .C1(new_n548), .C2(new_n420), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n477), .A2(G97), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT76), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n264), .A2(G97), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n336), .B1(new_n266), .B2(new_n476), .ZN(new_n568));
  OAI21_X1  g0368(.A(KEYINPUT76), .B1(new_n568), .B2(new_n565), .ZN(new_n569));
  OAI21_X1  g0369(.A(G107), .B1(new_n394), .B2(new_n395), .ZN(new_n570));
  XNOR2_X1  g0370(.A(G97), .B(G107), .ZN(new_n571));
  OR2_X1    g0371(.A1(KEYINPUT75), .A2(KEYINPUT6), .ZN(new_n572));
  OR2_X1    g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n571), .A2(new_n572), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n336), .A2(KEYINPUT6), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n573), .A2(new_n574), .A3(G20), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n255), .A2(G77), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n570), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n567), .A2(new_n569), .B1(new_n578), .B2(new_n260), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n304), .A2(new_n306), .A3(G244), .A4(new_n279), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT4), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n278), .A2(KEYINPUT4), .A3(G244), .A4(new_n279), .ZN(new_n583));
  NAND2_X1  g0383(.A1(G33), .A2(G283), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n278), .A2(G250), .A3(G1698), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n582), .A2(new_n583), .A3(new_n584), .A4(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n285), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n441), .A2(G257), .B1(G274), .B2(new_n439), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n589), .A2(G179), .ZN(new_n590));
  AOI21_X1  g0390(.A(G169), .B1(new_n587), .B2(new_n588), .ZN(new_n591));
  NOR3_X1   g0391(.A1(new_n579), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n567), .A2(new_n569), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n578), .A2(new_n260), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n587), .A2(new_n588), .A3(G190), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n589), .A2(G200), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(KEYINPUT77), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT77), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n579), .A2(new_n600), .A3(new_n597), .A4(new_n595), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n592), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n562), .A2(new_n602), .ZN(new_n603));
  NOR3_X1   g0403(.A1(new_n431), .A2(new_n521), .A3(new_n603), .ZN(G372));
  INV_X1    g0404(.A(new_n303), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n369), .A2(new_n325), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n427), .A2(new_n373), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n419), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n605), .B1(new_n608), .B2(new_n296), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n499), .A2(new_n420), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n491), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n504), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n512), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n471), .A2(new_n478), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n613), .B1(new_n614), .B2(new_n515), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n445), .A2(KEYINPUT83), .B1(new_n449), .B2(G179), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n448), .A2(new_n616), .B1(new_n518), .B2(new_n519), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n615), .B(new_n602), .C1(new_n617), .C2(new_n557), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n508), .A2(new_n512), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n593), .A2(new_n594), .ZN(new_n620));
  INV_X1    g0420(.A(new_n591), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n620), .B(new_n621), .C1(G179), .C2(new_n589), .ZN(new_n622));
  OAI21_X1  g0422(.A(KEYINPUT26), .B1(new_n619), .B2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n510), .B1(new_n315), .B2(new_n500), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n504), .A2(new_n611), .B1(new_n624), .B2(new_n509), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT26), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(new_n626), .A3(new_n592), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n623), .A2(new_n627), .A3(new_n512), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n618), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n609), .B1(new_n431), .B2(new_n629), .ZN(G369));
  NAND2_X1  g0430(.A1(new_n479), .A2(new_n520), .ZN(new_n631));
  INV_X1    g0431(.A(G13), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n632), .A2(G1), .A3(G20), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT84), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n634), .A2(new_n635), .A3(KEYINPUT27), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n635), .B1(new_n634), .B2(KEYINPUT27), .ZN(new_n637));
  OAI221_X1 g0437(.A(G213), .B1(KEYINPUT27), .B2(new_n634), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(G343), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n557), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n631), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n617), .A2(new_n641), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT85), .ZN(new_n647));
  XNOR2_X1  g0447(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n641), .A2(new_n559), .ZN(new_n649));
  MUX2_X1   g0449(.A(new_n562), .B(new_n557), .S(new_n649), .Z(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(G330), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n614), .A2(new_n641), .ZN(new_n653));
  OAI22_X1  g0453(.A1(new_n631), .A2(new_n653), .B1(new_n479), .B2(new_n641), .ZN(new_n654));
  INV_X1    g0454(.A(new_n642), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n648), .A2(new_n657), .ZN(G399));
  INV_X1    g0458(.A(new_n221), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(G41), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n484), .A2(new_n524), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n661), .A2(G1), .A3(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n230), .B2(new_n661), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n665), .B(KEYINPUT28), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n640), .B1(new_n618), .B2(new_n628), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT29), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(KEYINPUT87), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT87), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n671), .B1(new_n667), .B2(KEYINPUT29), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT88), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n617), .B2(new_n557), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n554), .A2(new_n555), .A3(KEYINPUT21), .ZN(new_n675));
  AOI21_X1  g0475(.A(KEYINPUT21), .B1(new_n554), .B2(new_n555), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n479), .A2(new_n677), .A3(KEYINPUT88), .A4(new_n550), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n674), .A2(new_n678), .A3(new_n602), .A4(new_n615), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n513), .A2(new_n626), .A3(new_n592), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT26), .B1(new_n613), .B2(new_n622), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n680), .A2(new_n681), .A3(new_n512), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n683), .A2(KEYINPUT29), .A3(new_n641), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n670), .A2(new_n672), .A3(new_n684), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n479), .A2(new_n513), .A3(new_n520), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n686), .A2(new_n562), .A3(new_n602), .A4(new_n641), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT30), .ZN(new_n688));
  OAI211_X1 g0488(.A(new_n551), .B(G179), .C1(new_n552), .C2(new_n553), .ZN(new_n689));
  AOI22_X1  g0489(.A1(new_n435), .A2(new_n285), .B1(new_n441), .B2(G264), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n690), .A2(new_n499), .A3(new_n587), .A4(new_n588), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n688), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n499), .A2(G179), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n554), .A2(new_n444), .A3(new_n589), .A4(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n689), .A2(new_n691), .A3(new_n688), .ZN(new_n696));
  OAI211_X1 g0496(.A(KEYINPUT31), .B(new_n640), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(KEYINPUT86), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n640), .B1(new_n695), .B2(new_n696), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT31), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n699), .A2(KEYINPUT86), .A3(new_n700), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n687), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G330), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n685), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n666), .B1(new_n706), .B2(G1), .ZN(G364));
  INV_X1    g0507(.A(KEYINPUT90), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n632), .A2(G20), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n709), .B(KEYINPUT89), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n206), .B1(new_n710), .B2(G45), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n708), .B1(new_n712), .B2(new_n660), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n661), .A2(KEYINPUT90), .A3(new_n711), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n652), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(G330), .B2(new_n650), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n221), .A2(G355), .A3(new_n278), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(G116), .B2(new_n221), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n659), .A2(new_n278), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(G45), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n722), .B1(new_n723), .B2(new_n231), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n245), .A2(new_n723), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n720), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n228), .B1(G20), .B2(new_n315), .ZN(new_n727));
  NOR2_X1   g0527(.A1(G13), .A2(G33), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G20), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n716), .B1(new_n726), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n207), .A2(new_n327), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n300), .A2(G200), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(G322), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n307), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n207), .A2(G190), .ZN(new_n739));
  NOR2_X1   g0539(.A1(G179), .A2(G200), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G329), .ZN(new_n743));
  INV_X1    g0543(.A(G283), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n420), .A2(G179), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(new_n739), .ZN(new_n746));
  INV_X1    g0546(.A(G311), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n735), .A2(new_n739), .ZN(new_n748));
  OAI221_X1 g0548(.A(new_n743), .B1(new_n744), .B2(new_n746), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT91), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n327), .ZN(new_n752));
  AOI211_X1 g0552(.A(new_n738), .B(new_n749), .C1(G326), .C2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n734), .A2(new_n745), .ZN(new_n754));
  OR2_X1    g0554(.A1(new_n754), .A2(KEYINPUT92), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(KEYINPUT92), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT94), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G303), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n207), .B1(new_n740), .B2(G190), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n760), .A2(KEYINPUT93), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(KEYINPUT93), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n751), .A2(G190), .ZN(new_n765));
  XNOR2_X1  g0565(.A(KEYINPUT33), .B(G317), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n764), .A2(G294), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n753), .A2(new_n759), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n742), .A2(G159), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT32), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n278), .B1(new_n748), .B2(new_n281), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n736), .A2(new_n211), .B1(new_n746), .B2(new_n461), .ZN(new_n772));
  NOR3_X1   g0572(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n757), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G87), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n764), .A2(G97), .ZN(new_n776));
  AOI22_X1  g0576(.A1(G50), .A2(new_n752), .B1(new_n765), .B2(G68), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n773), .A2(new_n775), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n768), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n733), .B1(new_n779), .B2(new_n727), .ZN(new_n780));
  INV_X1    g0580(.A(new_n730), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n780), .B1(new_n650), .B2(new_n781), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n718), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(G396));
  OAI21_X1  g0584(.A(new_n328), .B1(new_n323), .B2(new_n641), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n785), .A2(new_n325), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n325), .A2(new_n640), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n667), .B(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n716), .B1(new_n789), .B2(new_n705), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(new_n705), .B2(new_n789), .ZN(new_n791));
  INV_X1    g0591(.A(new_n727), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n758), .A2(G107), .ZN(new_n793));
  INV_X1    g0593(.A(G294), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n307), .B1(new_n736), .B2(new_n794), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n748), .A2(new_n524), .B1(new_n741), .B2(new_n747), .ZN(new_n796));
  INV_X1    g0596(.A(new_n746), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n795), .B(new_n796), .C1(G87), .C2(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(G283), .A2(new_n765), .B1(new_n752), .B2(G303), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n793), .A2(new_n776), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n736), .ZN(new_n801));
  INV_X1    g0601(.A(new_n748), .ZN(new_n802));
  AOI22_X1  g0602(.A1(G143), .A2(new_n801), .B1(new_n802), .B2(G159), .ZN(new_n803));
  INV_X1    g0603(.A(new_n752), .ZN(new_n804));
  INV_X1    g0604(.A(G137), .ZN(new_n805));
  INV_X1    g0605(.A(G150), .ZN(new_n806));
  INV_X1    g0606(.A(new_n765), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n803), .B1(new_n804), .B2(new_n805), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n808), .B(KEYINPUT34), .Z(new_n809));
  NOR2_X1   g0609(.A1(new_n746), .A2(new_n213), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n307), .B(new_n810), .C1(G132), .C2(new_n742), .ZN(new_n811));
  INV_X1    g0611(.A(new_n758), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n811), .B1(new_n211), .B2(new_n763), .C1(new_n812), .C2(new_n202), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n800), .B1(new_n809), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT96), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n792), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n815), .B2(new_n814), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n727), .A2(new_n728), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n715), .B1(new_n281), .B2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT95), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n817), .B(new_n820), .C1(new_n788), .C2(new_n729), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n791), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(G384));
  XOR2_X1   g0623(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n824));
  NOR2_X1   g0624(.A1(new_n399), .A2(new_n391), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n398), .B1(new_n396), .B2(new_n397), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n260), .B1(new_n826), .B2(new_n390), .ZN(new_n827));
  INV_X1    g0627(.A(new_n402), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n825), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n416), .B1(new_n829), .B2(new_n405), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(KEYINPUT18), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n407), .A2(new_n376), .A3(new_n416), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n427), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n638), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n829), .B2(new_n405), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n830), .A2(new_n835), .A3(new_n423), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT100), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT37), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(new_n835), .B2(KEYINPUT99), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n830), .A2(new_n835), .A3(KEYINPUT100), .A4(new_n423), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n840), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n837), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n842), .B1(new_n840), .B2(new_n843), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n824), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n415), .A2(new_n638), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n827), .A2(new_n406), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n841), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n838), .A2(new_n841), .B1(new_n423), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n833), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n849), .A2(new_n834), .ZN(new_n853));
  OAI211_X1 g0653(.A(KEYINPUT38), .B(new_n851), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n847), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n370), .A2(new_n641), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n374), .A2(new_n856), .B1(new_n369), .B2(new_n641), .ZN(new_n857));
  NOR3_X1   g0657(.A1(new_n603), .A2(new_n521), .A3(new_n640), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n701), .A2(new_n697), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n857), .B(new_n788), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n855), .A2(KEYINPUT40), .A3(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT101), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT38), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n853), .B1(new_n419), .B2(new_n427), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n838), .A2(new_n841), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n850), .A2(new_n423), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n865), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n854), .A2(new_n870), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n701), .A2(new_n697), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n687), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n873), .A2(KEYINPUT101), .A3(new_n788), .A4(new_n857), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n864), .A2(new_n871), .A3(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT40), .ZN(new_n876));
  AND3_X1   g0676(.A1(new_n875), .A2(KEYINPUT102), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT102), .B1(new_n875), .B2(new_n876), .ZN(new_n878));
  OAI211_X1 g0678(.A(G330), .B(new_n862), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n430), .A2(G330), .A3(new_n873), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n875), .A2(new_n876), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT102), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n875), .A2(KEYINPUT102), .A3(new_n876), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n886), .A2(new_n430), .A3(new_n873), .A4(new_n862), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n881), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT39), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n847), .A2(new_n889), .A3(new_n854), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n871), .A2(KEYINPUT39), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n369), .A2(new_n640), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n638), .B1(new_n417), .B2(new_n418), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n787), .B1(new_n667), .B2(new_n788), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n857), .ZN(new_n899));
  INV_X1    g0699(.A(new_n871), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n896), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n895), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n888), .B(new_n903), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n430), .A2(new_n672), .A3(new_n670), .A4(new_n684), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n609), .ZN(new_n906));
  OR2_X1    g0706(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n904), .A2(new_n906), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n907), .B(new_n908), .C1(new_n206), .C2(new_n710), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT35), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n910), .A2(new_n911), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n912), .A2(G116), .A3(new_n229), .A4(new_n913), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT36), .ZN(new_n915));
  OAI21_X1  g0715(.A(G77), .B1(new_n211), .B2(new_n213), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n916), .A2(new_n230), .B1(G50), .B2(new_n213), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(G1), .A3(new_n632), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n918), .B(KEYINPUT97), .Z(new_n919));
  NAND3_X1  g0719(.A1(new_n909), .A2(new_n915), .A3(new_n919), .ZN(G367));
  NAND2_X1  g0720(.A1(new_n620), .A2(new_n640), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n602), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n622), .A2(new_n641), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n648), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n925), .B(KEYINPUT45), .Z(new_n926));
  NOR2_X1   g0726(.A1(new_n648), .A2(new_n924), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT44), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n926), .A2(new_n928), .A3(new_n657), .ZN(new_n929));
  INV_X1    g0729(.A(new_n657), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n652), .A2(new_n656), .ZN(new_n931));
  NOR3_X1   g0731(.A1(new_n930), .A2(new_n643), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n706), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n929), .A2(new_n934), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n935), .A2(new_n706), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n660), .B(KEYINPUT41), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n711), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n922), .A2(new_n617), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n640), .B1(new_n940), .B2(new_n622), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n924), .A2(new_n643), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n941), .B1(new_n942), .B2(KEYINPUT42), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(KEYINPUT42), .B2(new_n942), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT43), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n625), .B1(new_n492), .B2(new_n641), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n624), .A2(new_n509), .A3(new_n491), .A4(new_n640), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n944), .B1(new_n945), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n945), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n930), .A2(new_n924), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n952), .B(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n939), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n278), .B1(new_n736), .B2(new_n806), .ZN(new_n956));
  AOI22_X1  g0756(.A1(G77), .A2(new_n797), .B1(new_n742), .B2(G137), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n202), .B2(new_n748), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n956), .B(new_n958), .C1(G58), .C2(new_n774), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n752), .A2(G143), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n764), .A2(G68), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n765), .A2(G159), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n959), .A2(new_n960), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n758), .A2(KEYINPUT46), .A3(G116), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n801), .A2(G303), .B1(new_n742), .B2(G317), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n744), .B2(new_n748), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n746), .A2(new_n336), .ZN(new_n967));
  NOR3_X1   g0767(.A1(new_n966), .A2(new_n278), .A3(new_n967), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n964), .B(new_n968), .C1(new_n794), .C2(new_n807), .ZN(new_n969));
  XOR2_X1   g0769(.A(KEYINPUT104), .B(KEYINPUT46), .Z(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n757), .B2(new_n524), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n971), .B1(new_n461), .B2(new_n763), .C1(new_n747), .C2(new_n804), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n963), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT47), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n792), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n974), .B2(new_n973), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n241), .A2(new_n721), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n977), .B(new_n731), .C1(new_n221), .C2(new_n488), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n978), .A2(KEYINPUT103), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n978), .A2(KEYINPUT103), .ZN(new_n980));
  NOR3_X1   g0780(.A1(new_n979), .A2(new_n980), .A3(new_n715), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n976), .B(new_n981), .C1(new_n781), .C2(new_n948), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n955), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(G387));
  NOR2_X1   g0784(.A1(new_n934), .A2(new_n661), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n706), .B2(new_n932), .ZN(new_n986));
  AOI21_X1  g0786(.A(G45), .B1(G68), .B2(G77), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n252), .A2(new_n202), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n663), .B(new_n987), .C1(new_n988), .C2(KEYINPUT50), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(KEYINPUT50), .B2(new_n988), .ZN(new_n990));
  INV_X1    g0790(.A(new_n236), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n721), .B1(new_n991), .B2(new_n723), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n221), .A2(new_n278), .A3(new_n662), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n990), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n221), .A2(G107), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n731), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n716), .ZN(new_n997));
  AOI22_X1  g0797(.A1(G50), .A2(new_n801), .B1(new_n802), .B2(G68), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n806), .B2(new_n741), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n757), .A2(new_n281), .ZN(new_n1000));
  NOR4_X1   g0800(.A1(new_n999), .A2(new_n1000), .A3(new_n307), .A4(new_n967), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n752), .A2(G159), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n765), .A2(new_n252), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n764), .A2(new_n320), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n278), .B1(new_n742), .B2(G326), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(G317), .A2(new_n801), .B1(new_n802), .B2(G303), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1007), .B1(new_n804), .B2(new_n737), .C1(new_n747), .C2(new_n807), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(KEYINPUT48), .Z(new_n1009));
  OAI22_X1  g0809(.A1(new_n757), .A2(new_n794), .B1(new_n763), .B2(new_n744), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1006), .B1(new_n524), .B2(new_n746), .C1(new_n1011), .C2(KEYINPUT49), .ZN(new_n1012));
  AND2_X1   g0812(.A1(new_n1011), .A2(KEYINPUT49), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1005), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n997), .B1(new_n1014), .B2(new_n727), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n654), .B2(new_n781), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT105), .Z(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(new_n712), .B2(new_n932), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n986), .A2(new_n1018), .ZN(G393));
  NAND2_X1  g0819(.A1(new_n926), .A2(new_n928), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(new_n657), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1021), .A2(new_n934), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n935), .A2(new_n660), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1021), .A2(new_n712), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n307), .B1(new_n741), .B2(new_n737), .C1(new_n461), .C2(new_n746), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n774), .B2(G283), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT106), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n763), .A2(new_n524), .B1(new_n794), .B2(new_n748), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G303), .B2(new_n765), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n752), .A2(G317), .B1(G311), .B2(new_n801), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT52), .Z(new_n1033));
  NAND3_X1  g0833(.A1(new_n1029), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(G159), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n804), .A2(new_n806), .B1(new_n1035), .B2(new_n736), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT51), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n307), .B1(new_n797), .B2(G87), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n742), .A2(G143), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n252), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1039), .B(new_n1040), .C1(new_n1041), .C2(new_n748), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n757), .A2(new_n213), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1042), .B(new_n1043), .C1(G50), .C2(new_n765), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n764), .A2(G77), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1034), .B1(new_n1038), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT107), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n792), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n1049), .B2(new_n1048), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n731), .B1(new_n336), .B2(new_n221), .C1(new_n722), .C2(new_n249), .ZN(new_n1052));
  AND2_X1   g0852(.A1(new_n716), .A2(new_n1052), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1051), .B(new_n1053), .C1(new_n924), .C2(new_n781), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1026), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1025), .A2(new_n1056), .ZN(G390));
  NAND2_X1  g0857(.A1(new_n892), .A2(new_n728), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n715), .B1(new_n1041), .B2(new_n818), .ZN(new_n1059));
  INV_X1    g0859(.A(G87), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n307), .B1(new_n812), .B2(new_n1060), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1061), .A2(KEYINPUT111), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G107), .A2(new_n765), .B1(new_n752), .B2(G283), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n810), .B1(G294), .B2(new_n742), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G116), .A2(new_n801), .B1(new_n802), .B2(G97), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1046), .A2(new_n1063), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n1061), .B2(KEYINPUT111), .ZN(new_n1067));
  INV_X1    g0867(.A(G132), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n278), .B1(new_n736), .B2(new_n1068), .ZN(new_n1069));
  XOR2_X1   g0869(.A(KEYINPUT54), .B(G143), .Z(new_n1070));
  NAND2_X1  g0870(.A1(new_n802), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n742), .A2(G125), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1071), .B(new_n1072), .C1(new_n202), .C2(new_n746), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1069), .B(new_n1073), .C1(G159), .C2(new_n764), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT53), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(new_n774), .B2(G150), .ZN(new_n1076));
  INV_X1    g0876(.A(G128), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n1077), .A2(new_n804), .B1(new_n807), .B2(new_n805), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n757), .A2(KEYINPUT53), .A3(new_n806), .ZN(new_n1079));
  NOR3_X1   g0879(.A1(new_n1076), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n1062), .A2(new_n1067), .B1(new_n1074), .B2(new_n1080), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1058), .B(new_n1059), .C1(new_n792), .C2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n857), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n894), .B1(new_n897), .B2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n890), .A2(new_n891), .A3(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n704), .A2(G330), .A3(new_n788), .ZN(new_n1086));
  OR2_X1    g0886(.A1(new_n1086), .A2(new_n1083), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n640), .B(new_n786), .C1(new_n679), .C2(new_n682), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n857), .B1(new_n1088), .B2(new_n787), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n855), .A2(new_n894), .A3(new_n1089), .ZN(new_n1090));
  AND3_X1   g0890(.A1(new_n1085), .A2(new_n1087), .A3(new_n1090), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n873), .A2(G330), .A3(new_n788), .A4(new_n857), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n1085), .B2(new_n1090), .ZN(new_n1093));
  OAI21_X1  g0893(.A(KEYINPUT108), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1085), .A2(new_n1087), .A3(new_n1090), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT108), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1082), .B1(new_n1098), .B2(new_n711), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n905), .A2(new_n609), .A3(new_n880), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT109), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n861), .A2(G330), .B1(new_n1086), .B2(new_n1083), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1101), .B1(new_n1102), .B2(new_n897), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1086), .A2(new_n1083), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n1092), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1105), .A2(KEYINPUT109), .A3(new_n898), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1088), .A2(new_n787), .ZN(new_n1108));
  AND3_X1   g0908(.A1(new_n873), .A2(G330), .A3(new_n788), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1087), .B(new_n1108), .C1(new_n857), .C2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1100), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1094), .A2(new_n1097), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(KEYINPUT110), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT110), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1094), .A2(new_n1111), .A3(new_n1114), .A4(new_n1097), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1100), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n661), .B1(new_n1098), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1099), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(G378));
  NAND2_X1  g0922(.A1(new_n296), .A2(new_n303), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n290), .A2(new_n638), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1123), .B(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1126));
  XOR2_X1   g0926(.A(new_n1125), .B(new_n1126), .Z(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n728), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n727), .A2(G50), .A3(new_n728), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n961), .B1(new_n336), .B2(new_n807), .C1(new_n524), .C2(new_n804), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n273), .B(new_n307), .C1(new_n736), .C2(new_n461), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n320), .A2(new_n802), .B1(new_n797), .B2(G58), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n744), .B2(new_n741), .ZN(new_n1134));
  NOR4_X1   g0934(.A1(new_n1131), .A2(new_n1000), .A3(new_n1132), .A4(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT112), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(KEYINPUT113), .B(KEYINPUT58), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1136), .B(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(G50), .B1(new_n259), .B2(new_n273), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n278), .B2(G41), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n774), .A2(new_n1070), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT115), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n765), .A2(G132), .B1(G137), .B2(new_n802), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1143), .B(KEYINPUT114), .Z(new_n1144));
  OAI22_X1  g0944(.A1(new_n763), .A2(new_n806), .B1(new_n1077), .B2(new_n736), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(G125), .B2(new_n752), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1142), .A2(new_n1144), .A3(new_n1146), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1147), .A2(KEYINPUT59), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(KEYINPUT59), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n797), .A2(G159), .ZN(new_n1150));
  AOI211_X1 g0950(.A(G33), .B(G41), .C1(new_n742), .C2(G124), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1138), .B(new_n1140), .C1(new_n1148), .C2(new_n1152), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n715), .B(new_n1130), .C1(new_n1153), .C2(new_n727), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1129), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n879), .A2(new_n1128), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n886), .A2(G330), .A3(new_n862), .A4(new_n1127), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT116), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n903), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  AOI211_X1 g0960(.A(KEYINPUT116), .B(new_n902), .C1(new_n1156), .C2(new_n1157), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1155), .B1(new_n1162), .B2(new_n711), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT57), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1158), .A2(new_n903), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1156), .A2(new_n1157), .A3(new_n902), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1165), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n661), .B1(new_n1164), .B2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1100), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1165), .B1(new_n1162), .B2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1163), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(G375));
  NAND3_X1  g0973(.A1(new_n1107), .A2(new_n1100), .A3(new_n1110), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1119), .A2(new_n937), .A3(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT117), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1004), .B1(new_n744), .B2(new_n736), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT118), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n807), .A2(new_n524), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(G107), .A2(new_n802), .B1(new_n742), .B2(G303), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1180), .B(new_n307), .C1(new_n281), .C2(new_n746), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1179), .B(new_n1181), .C1(G294), .C2(new_n752), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1178), .B(new_n1182), .C1(new_n336), .C2(new_n812), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n278), .B1(new_n746), .B2(new_n211), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(G150), .A2(new_n802), .B1(new_n742), .B2(G128), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n805), .B2(new_n736), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1184), .B(new_n1186), .C1(new_n765), .C2(new_n1070), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n764), .A2(G50), .B1(G132), .B2(new_n752), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1187), .B(new_n1188), .C1(new_n1035), .C2(new_n812), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n792), .B1(new_n1183), .B2(new_n1189), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n715), .B(new_n1190), .C1(new_n213), .C2(new_n818), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT119), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n728), .B2(new_n1083), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n1117), .B2(new_n712), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1176), .A2(new_n1194), .ZN(G381));
  NAND3_X1  g0995(.A1(new_n986), .A2(new_n783), .A3(new_n1018), .ZN(new_n1196));
  NOR4_X1   g0996(.A1(G387), .A2(G384), .A3(G390), .A4(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT120), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1085), .A2(new_n1090), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1092), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1096), .B1(new_n1201), .B2(new_n1095), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1097), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1119), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(new_n660), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(new_n1115), .B2(new_n1113), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1198), .B1(new_n1206), .B2(new_n1099), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1121), .A2(KEYINPUT120), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(G375), .A2(new_n1210), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1197), .A2(new_n1211), .A3(new_n1194), .A4(new_n1176), .ZN(G407));
  NAND2_X1  g1012(.A1(new_n639), .A2(G213), .ZN(new_n1213));
  NOR3_X1   g1013(.A1(G375), .A2(new_n1210), .A3(new_n1213), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n1214), .A2(KEYINPUT121), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(KEYINPUT121), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1215), .A2(G213), .A3(G407), .A4(new_n1216), .ZN(G409));
  INV_X1    g1017(.A(KEYINPUT124), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1196), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n783), .B1(new_n986), .B2(new_n1018), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1025), .B(new_n1056), .C1(new_n1219), .C2(new_n1220), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n1024), .B2(new_n1055), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1221), .A2(new_n1223), .A3(new_n983), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n983), .B1(new_n1221), .B2(new_n1223), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1218), .B1(new_n1227), .B2(KEYINPUT61), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT61), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1226), .A2(KEYINPUT124), .A3(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1213), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT116), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1232), .B(new_n903), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1233), .A2(new_n1164), .A3(new_n937), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1155), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1235), .B1(new_n1236), .B2(new_n712), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1234), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1209), .A2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1235), .B1(new_n1233), .B2(new_n712), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT57), .B1(new_n1233), .B2(new_n1164), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1236), .A2(KEYINPUT57), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n660), .B1(new_n1242), .B2(new_n1170), .ZN(new_n1243));
  OAI211_X1 g1043(.A(G378), .B(new_n1240), .C1(new_n1241), .C2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1231), .B1(new_n1239), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT60), .ZN(new_n1247));
  OR2_X1    g1047(.A1(new_n1174), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1174), .A2(new_n1247), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1248), .A2(new_n660), .A3(new_n1119), .A4(new_n1249), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1250), .A2(G384), .A3(new_n1194), .ZN(new_n1251));
  AOI21_X1  g1051(.A(G384), .B1(new_n1250), .B2(new_n1194), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1231), .A2(G2897), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1254), .A2(KEYINPUT123), .A3(new_n1255), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1254), .A2(KEYINPUT123), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT123), .ZN(new_n1258));
  OAI211_X1 g1058(.A(G2897), .B(new_n1231), .C1(new_n1253), .C2(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1256), .B1(new_n1257), .B2(new_n1259), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n1228), .A2(new_n1230), .B1(new_n1246), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT125), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n1172), .A2(G378), .B1(new_n1209), .B2(new_n1238), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1262), .B1(new_n1263), .B2(new_n1231), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1239), .A2(new_n1244), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1265), .A2(KEYINPUT125), .A3(new_n1213), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1267), .A2(KEYINPUT63), .A3(new_n1253), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(KEYINPUT122), .B(KEYINPUT63), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n1246), .B2(new_n1254), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1261), .A2(new_n1268), .A3(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1264), .A2(new_n1266), .A3(new_n1260), .ZN(new_n1272));
  AND3_X1   g1072(.A1(new_n1272), .A2(KEYINPUT126), .A3(new_n1229), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT126), .B1(new_n1272), .B2(new_n1229), .ZN(new_n1274));
  AOI21_X1  g1074(.A(KEYINPUT62), .B1(new_n1245), .B2(new_n1253), .ZN(new_n1275));
  AND2_X1   g1075(.A1(new_n1253), .A2(KEYINPUT62), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1275), .B1(new_n1267), .B2(new_n1276), .ZN(new_n1277));
  NOR3_X1   g1077(.A1(new_n1273), .A2(new_n1274), .A3(new_n1277), .ZN(new_n1278));
  XOR2_X1   g1078(.A(new_n1226), .B(KEYINPUT127), .Z(new_n1279));
  OAI21_X1  g1079(.A(new_n1271), .B1(new_n1278), .B2(new_n1279), .ZN(G405));
  OAI21_X1  g1080(.A(new_n1244), .B1(new_n1210), .B2(new_n1172), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1281), .B(new_n1253), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(new_n1282), .B(new_n1227), .ZN(G402));
endmodule


