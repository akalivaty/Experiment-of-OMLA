//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 1 0 1 0 0 1 0 0 1 1 0 1 1 0 1 1 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 0 0 1 1 0 0 0 0 0 0 1 0 0 0 1 1 0 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1252, new_n1253, new_n1254, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(new_n204));
  NOR3_X1   g0004(.A1(new_n202), .A2(G77), .A3(new_n204), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(KEYINPUT65), .B(KEYINPUT0), .Z(new_n213));
  XNOR2_X1  g0013(.A(new_n212), .B(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n210), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT1), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(KEYINPUT66), .ZN(new_n224));
  INV_X1    g0024(.A(KEYINPUT66), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n225), .A2(G1), .A3(G13), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OR2_X1    g0030(.A1(new_n203), .A2(KEYINPUT67), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n203), .A2(KEYINPUT67), .ZN(new_n232));
  NAND3_X1  g0032(.A1(new_n231), .A2(G50), .A3(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n214), .B(new_n222), .C1(new_n230), .C2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT2), .B(G226), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XOR2_X1   g0045(.A(G50), .B(G58), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  NAND2_X1  g0051(.A1(G33), .A2(G41), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n252), .A2(G1), .A3(G13), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G274), .ZN(new_n254));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  INV_X1    g0055(.A(G45), .ZN(new_n256));
  AOI21_X1  g0056(.A(G1), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G226), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n258), .A2(new_n253), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT3), .B(G33), .ZN(new_n264));
  INV_X1    g0064(.A(G1698), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n264), .A2(G222), .A3(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G77), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n264), .A2(G1698), .ZN(new_n268));
  INV_X1    g0068(.A(G223), .ZN(new_n269));
  OAI221_X1 g0069(.A(new_n266), .B1(new_n267), .B2(new_n264), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  AND2_X1   g0070(.A1(new_n227), .A2(new_n252), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n263), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G169), .ZN(new_n273));
  INV_X1    g0073(.A(G179), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n273), .B1(new_n274), .B2(new_n272), .ZN(new_n275));
  NAND3_X1  g0075(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n224), .A2(new_n226), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n229), .B1(new_n201), .B2(new_n203), .ZN(new_n278));
  XNOR2_X1  g0078(.A(new_n278), .B(KEYINPUT70), .ZN(new_n279));
  NOR2_X1   g0079(.A1(KEYINPUT8), .A2(G58), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT68), .B(G58), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n280), .B1(new_n281), .B2(KEYINPUT8), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n229), .A2(G33), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G20), .A2(G33), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n282), .A2(new_n284), .B1(G150), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT69), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n279), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n286), .A2(new_n287), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n277), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G1), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(G13), .A3(G20), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n224), .A2(new_n226), .A3(new_n293), .A4(new_n276), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(G20), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G50), .ZN(new_n296));
  OAI22_X1  g0096(.A1(new_n294), .A2(new_n296), .B1(G50), .B2(new_n293), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n291), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n275), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT10), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n299), .B(KEYINPUT9), .ZN(new_n302));
  INV_X1    g0102(.A(G200), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n272), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n304), .B1(G190), .B2(new_n272), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n301), .B1(new_n302), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n299), .A2(KEYINPUT9), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT9), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n308), .B1(new_n291), .B2(new_n298), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n301), .B(new_n305), .C1(new_n307), .C2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n300), .B1(new_n306), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n227), .A2(new_n252), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n264), .A2(G232), .A3(G1698), .ZN(new_n314));
  NAND2_X1  g0114(.A1(G33), .A2(G97), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G33), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT3), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT3), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G33), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n318), .A2(new_n320), .A3(G226), .A4(new_n265), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT71), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT71), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n264), .A2(new_n323), .A3(G226), .A4(new_n265), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n313), .B1(new_n316), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G238), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n260), .B1(new_n327), .B2(new_n262), .ZN(new_n328));
  OAI21_X1  g0128(.A(KEYINPUT13), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT13), .ZN(new_n330));
  INV_X1    g0130(.A(new_n262), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n259), .B1(new_n331), .B2(G238), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n314), .A2(new_n315), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n333), .B1(new_n324), .B2(new_n322), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n330), .B(new_n332), .C1(new_n334), .C2(new_n313), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n329), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(G200), .ZN(new_n337));
  INV_X1    g0137(.A(G68), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n285), .A2(G50), .B1(G20), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n339), .B1(new_n267), .B2(new_n283), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n340), .A2(new_n277), .ZN(new_n341));
  OR2_X1    g0141(.A1(new_n341), .A2(KEYINPUT11), .ZN(new_n342));
  INV_X1    g0142(.A(new_n293), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n338), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n344), .B(KEYINPUT12), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n341), .A2(KEYINPUT11), .ZN(new_n346));
  INV_X1    g0146(.A(new_n294), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n347), .A2(G68), .A3(new_n295), .ZN(new_n348));
  AND4_X1   g0148(.A1(new_n342), .A2(new_n345), .A3(new_n346), .A4(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n329), .A2(new_n335), .A3(G190), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n337), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT72), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(new_n336), .B2(new_n274), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n329), .A2(new_n335), .A3(KEYINPUT72), .A4(G179), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n336), .A2(G169), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT14), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT14), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n336), .A2(new_n359), .A3(G169), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n356), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n349), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n352), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n203), .B1(new_n281), .B2(G68), .ZN(new_n365));
  INV_X1    g0165(.A(G159), .ZN(new_n366));
  INV_X1    g0166(.A(new_n285), .ZN(new_n367));
  OAI22_X1  g0167(.A1(new_n365), .A2(new_n229), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n318), .A2(new_n320), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n370), .A2(KEYINPUT7), .A3(new_n229), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT73), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n264), .A2(KEYINPUT73), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n374), .A2(new_n375), .A3(new_n229), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n372), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OAI211_X1 g0178(.A(KEYINPUT16), .B(new_n369), .C1(new_n378), .C2(new_n338), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT16), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n377), .B1(new_n264), .B2(G20), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n338), .B1(new_n381), .B2(new_n371), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n380), .B1(new_n368), .B2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n379), .A2(new_n383), .A3(new_n277), .ZN(new_n384));
  AND2_X1   g0184(.A1(new_n282), .A2(new_n295), .ZN(new_n385));
  INV_X1    g0185(.A(new_n282), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n385), .A2(new_n347), .B1(new_n343), .B2(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n318), .A2(new_n320), .A3(G223), .A4(new_n265), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n318), .A2(new_n320), .A3(G226), .A4(G1698), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G33), .A2(G87), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT74), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT74), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n388), .A2(new_n389), .A3(new_n393), .A4(new_n390), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n392), .A2(new_n271), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n259), .B1(new_n331), .B2(G232), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(G200), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n395), .A2(G190), .A3(new_n396), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n384), .A2(new_n387), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  XNOR2_X1  g0200(.A(new_n400), .B(KEYINPUT17), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n384), .A2(new_n387), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT75), .ZN(new_n403));
  AOI21_X1  g0203(.A(G169), .B1(new_n395), .B2(new_n396), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n395), .A2(new_n274), .A3(new_n396), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n403), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n406), .ZN(new_n408));
  NOR3_X1   g0208(.A1(new_n408), .A2(new_n404), .A3(KEYINPUT75), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n402), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT18), .ZN(new_n411));
  OAI21_X1  g0211(.A(KEYINPUT75), .B1(new_n408), .B2(new_n404), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n405), .A2(new_n403), .A3(new_n406), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n412), .A2(new_n413), .B1(new_n384), .B2(new_n387), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT18), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n401), .A2(new_n411), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n347), .A2(G77), .A3(new_n295), .ZN(new_n418));
  XOR2_X1   g0218(.A(KEYINPUT8), .B(G58), .Z(new_n419));
  AOI22_X1  g0219(.A1(new_n419), .A2(new_n285), .B1(G20), .B2(G77), .ZN(new_n420));
  XNOR2_X1  g0220(.A(KEYINPUT15), .B(G87), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n420), .B1(new_n283), .B2(new_n421), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n422), .A2(new_n277), .B1(new_n267), .B2(new_n343), .ZN(new_n423));
  OAI22_X1  g0223(.A1(new_n268), .A2(new_n327), .B1(new_n207), .B2(new_n264), .ZN(new_n424));
  NOR3_X1   g0224(.A1(new_n370), .A2(new_n237), .A3(G1698), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n271), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n259), .B1(new_n331), .B2(G244), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(G169), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n418), .A2(new_n423), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n428), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n274), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n431), .A2(new_n303), .ZN(new_n435));
  INV_X1    g0235(.A(G190), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n428), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n423), .A2(new_n418), .ZN(new_n438));
  NOR3_X1   g0238(.A1(new_n435), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NOR4_X1   g0241(.A1(new_n312), .A2(new_n364), .A3(new_n417), .A4(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT21), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n343), .A2(G116), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n292), .A2(G33), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n347), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n445), .B1(new_n447), .B2(G116), .ZN(new_n448));
  NAND2_X1  g0248(.A1(G33), .A2(G283), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n449), .B(new_n229), .C1(G33), .C2(new_n206), .ZN(new_n450));
  INV_X1    g0250(.A(G116), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(G20), .ZN(new_n452));
  AND3_X1   g0252(.A1(new_n277), .A2(KEYINPUT80), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT80), .B1(new_n277), .B2(new_n452), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n450), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT20), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI211_X1 g0257(.A(KEYINPUT20), .B(new_n450), .C1(new_n453), .C2(new_n454), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n448), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  XNOR2_X1  g0259(.A(KEYINPUT5), .B(G41), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n256), .A2(G1), .ZN(new_n461));
  INV_X1    g0261(.A(new_n223), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n460), .A2(new_n461), .B1(new_n462), .B2(new_n252), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n253), .A2(G274), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n292), .A2(G45), .ZN(new_n465));
  NOR2_X1   g0265(.A1(KEYINPUT5), .A2(G41), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(KEYINPUT5), .A2(G41), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n463), .A2(G270), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n319), .A2(G33), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n317), .A2(KEYINPUT3), .ZN(new_n472));
  OAI21_X1  g0272(.A(G303), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n318), .A2(new_n320), .A3(G264), .A4(G1698), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n318), .A2(new_n320), .A3(G257), .A4(new_n265), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n271), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n470), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(G169), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n444), .B1(new_n459), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT81), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI211_X1 g0282(.A(KEYINPUT81), .B(new_n444), .C1(new_n459), .C2(new_n479), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n457), .A2(new_n458), .ZN(new_n485));
  INV_X1    g0285(.A(new_n448), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI22_X1  g0287(.A1(new_n479), .A2(new_n444), .B1(new_n274), .B2(new_n478), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n478), .A2(G200), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n459), .B(new_n490), .C1(new_n436), .C2(new_n478), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n484), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(KEYINPUT23), .B1(new_n229), .B2(G107), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT23), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n495), .A2(new_n207), .A3(G20), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n229), .A2(G33), .A3(G116), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT82), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT24), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n494), .A2(new_n496), .A3(new_n497), .A4(new_n499), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n318), .A2(new_n320), .A3(new_n229), .A4(G87), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT22), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT22), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n264), .A2(new_n503), .A3(new_n229), .A4(G87), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n500), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  OR2_X1    g0305(.A1(new_n498), .A2(KEYINPUT24), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  AOI211_X1 g0308(.A(new_n506), .B(new_n500), .C1(new_n502), .C2(new_n504), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n277), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(KEYINPUT25), .B1(new_n343), .B2(new_n207), .ZN(new_n511));
  XNOR2_X1  g0311(.A(new_n511), .B(KEYINPUT84), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n343), .A2(KEYINPUT25), .A3(new_n207), .ZN(new_n513));
  XNOR2_X1  g0313(.A(new_n513), .B(KEYINPUT83), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n294), .B1(new_n292), .B2(G33), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n512), .A2(new_n514), .B1(G107), .B2(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n318), .A2(new_n320), .A3(G250), .A4(new_n265), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT85), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n264), .A2(KEYINPUT85), .A3(G250), .A4(new_n265), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G33), .A2(G294), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n264), .A2(G257), .A3(G1698), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n519), .A2(new_n520), .A3(new_n521), .A4(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n468), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n461), .B1(new_n524), .B2(new_n466), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n525), .A2(G264), .A3(new_n253), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(KEYINPUT86), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT86), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n525), .A2(new_n528), .A3(G264), .A4(new_n253), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n523), .A2(new_n271), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n460), .A2(new_n253), .A3(G274), .A4(new_n461), .ZN(new_n531));
  AOI21_X1  g0331(.A(G200), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n526), .A2(new_n531), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n533), .B1(new_n523), .B2(new_n271), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n534), .A2(new_n436), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n510), .B(new_n516), .C1(new_n532), .C2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n523), .A2(new_n271), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n527), .A2(new_n529), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(new_n531), .A3(new_n538), .ZN(new_n539));
  OAI22_X1  g0339(.A1(new_n539), .A2(new_n274), .B1(new_n429), .B2(new_n534), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n510), .A2(new_n516), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n536), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT6), .ZN(new_n544));
  NOR3_X1   g0344(.A1(new_n544), .A2(new_n206), .A3(G107), .ZN(new_n545));
  XNOR2_X1  g0345(.A(G97), .B(G107), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n545), .B1(new_n546), .B2(new_n544), .ZN(new_n547));
  OAI22_X1  g0347(.A1(new_n547), .A2(new_n229), .B1(new_n267), .B2(new_n367), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n207), .B1(new_n381), .B2(new_n371), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n277), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n293), .A2(G97), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n551), .B1(new_n515), .B2(G97), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n318), .A2(new_n320), .A3(G244), .A4(new_n265), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT4), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n264), .A2(KEYINPUT4), .A3(G244), .A4(new_n265), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n264), .A2(G250), .A3(G1698), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n555), .A2(new_n556), .A3(new_n449), .A4(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n271), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n525), .A2(G257), .A3(new_n253), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n531), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n550), .B(new_n552), .C1(new_n563), .C2(new_n436), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT76), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n561), .B1(new_n558), .B2(new_n271), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT76), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(G200), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n274), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n563), .A2(new_n429), .B1(new_n550), .B2(new_n552), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n565), .A2(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n253), .A2(G250), .A3(new_n465), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n254), .B2(new_n465), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n318), .A2(new_n320), .A3(G244), .A4(G1698), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT77), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT77), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n264), .A2(new_n578), .A3(G244), .A4(G1698), .ZN(new_n579));
  NAND2_X1  g0379(.A1(G33), .A2(G116), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n264), .A2(G238), .A3(new_n265), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n577), .A2(new_n579), .A3(new_n580), .A4(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n575), .B1(new_n582), .B2(new_n271), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n274), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT19), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n229), .B1(new_n315), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(G87), .B2(new_n208), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n318), .A2(new_n320), .A3(new_n229), .A4(G68), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n585), .B1(new_n283), .B2(new_n206), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n277), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT78), .ZN(new_n592));
  OR2_X1    g0392(.A1(new_n421), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n421), .A2(new_n592), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n347), .A2(new_n593), .A3(new_n446), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n421), .A2(new_n343), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n591), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n584), .B(new_n597), .C1(G169), .C2(new_n583), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n582), .A2(new_n271), .ZN(new_n599));
  INV_X1    g0399(.A(new_n575), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(G190), .A3(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n347), .A2(G87), .A3(new_n446), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n591), .A2(new_n596), .A3(new_n602), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n601), .B(new_n603), .C1(new_n303), .C2(new_n583), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n598), .A2(KEYINPUT79), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(KEYINPUT79), .B1(new_n598), .B2(new_n604), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n573), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NOR4_X1   g0407(.A1(new_n443), .A2(new_n493), .A3(new_n543), .A4(new_n607), .ZN(G372));
  XNOR2_X1  g0408(.A(new_n598), .B(KEYINPUT87), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n489), .A2(new_n542), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n611), .B1(new_n482), .B2(new_n483), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n601), .A2(new_n603), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n583), .A2(new_n303), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n597), .B1(new_n583), .B2(G169), .ZN(new_n615));
  AOI211_X1 g0415(.A(G179), .B(new_n575), .C1(new_n582), .C2(new_n271), .ZN(new_n616));
  OAI22_X1  g0416(.A1(new_n613), .A2(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n573), .A2(new_n536), .A3(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n610), .B1(new_n612), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n550), .A2(new_n552), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n621), .B(new_n571), .C1(G169), .C2(new_n568), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(KEYINPUT26), .B1(new_n618), .B2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT79), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n617), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n598), .A2(KEYINPUT79), .A3(new_n604), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n622), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n624), .B1(new_n628), .B2(KEYINPUT26), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n442), .B1(new_n620), .B2(new_n629), .ZN(new_n630));
  XNOR2_X1  g0430(.A(new_n630), .B(KEYINPUT88), .ZN(new_n631));
  OR2_X1    g0431(.A1(new_n306), .A2(new_n311), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n412), .A2(new_n413), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n633), .A2(new_n415), .A3(new_n402), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n415), .B1(new_n633), .B2(new_n402), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n361), .A2(new_n362), .B1(new_n351), .B2(new_n434), .ZN(new_n637));
  INV_X1    g0437(.A(new_n401), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n632), .A2(new_n639), .B1(new_n299), .B2(new_n275), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n631), .A2(new_n640), .ZN(G369));
  NAND3_X1  g0441(.A1(new_n292), .A2(new_n229), .A3(G13), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT27), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n644), .A2(new_n292), .A3(new_n229), .A4(G13), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n643), .A2(G213), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g0446(.A(new_n646), .B(KEYINPUT89), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(G343), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT90), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT90), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n647), .A2(new_n651), .A3(G343), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n492), .B1(new_n459), .B2(new_n654), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n487), .A2(new_n488), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n656), .B1(new_n482), .B2(new_n483), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n653), .A2(new_n487), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(G330), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n653), .A2(new_n541), .ZN(new_n662));
  OAI22_X1  g0462(.A1(new_n543), .A2(new_n662), .B1(new_n542), .B2(new_n654), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n657), .A2(new_n543), .A3(new_n653), .ZN(new_n665));
  INV_X1    g0465(.A(new_n542), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n665), .B1(new_n666), .B2(new_n654), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n664), .A2(new_n667), .ZN(G399));
  INV_X1    g0468(.A(KEYINPUT91), .ZN(new_n669));
  INV_X1    g0469(.A(new_n211), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n669), .B1(new_n670), .B2(G41), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n211), .A2(KEYINPUT91), .A3(new_n255), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n208), .A2(G87), .A3(G116), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G1), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n233), .B2(new_n673), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT28), .ZN(new_n677));
  INV_X1    g0477(.A(G330), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n470), .A2(new_n477), .A3(G179), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n679), .A2(new_n530), .A3(new_n568), .A4(new_n583), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT30), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT93), .ZN(new_n682));
  AOI21_X1  g0482(.A(G179), .B1(new_n470), .B2(new_n477), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n539), .A2(new_n563), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT92), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n583), .B(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n682), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n685), .B1(new_n599), .B2(new_n600), .ZN(new_n688));
  AOI211_X1 g0488(.A(KEYINPUT92), .B(new_n575), .C1(new_n582), .C2(new_n271), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n539), .A2(new_n563), .A3(new_n683), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n690), .A2(new_n691), .A3(KEYINPUT93), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n681), .B1(new_n687), .B2(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(KEYINPUT31), .B1(new_n693), .B2(new_n653), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n653), .A2(KEYINPUT31), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n684), .A2(new_n686), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n695), .B1(new_n681), .B2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(G200), .B1(new_n568), .B2(KEYINPUT76), .ZN(new_n699));
  AOI211_X1 g0499(.A(new_n566), .B(new_n561), .C1(new_n558), .C2(new_n271), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n622), .B1(new_n701), .B2(new_n564), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n702), .B1(new_n626), .B2(new_n627), .ZN(new_n703));
  AND3_X1   g0503(.A1(new_n536), .A2(new_n654), .A3(new_n542), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n703), .A2(new_n657), .A3(new_n491), .A4(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n678), .B1(new_n698), .B2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT95), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT26), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n617), .A2(new_n708), .A3(new_n622), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n623), .B1(new_n605), .B2(new_n606), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n709), .B1(new_n710), .B2(new_n708), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n654), .B1(new_n620), .B2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT29), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n707), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n611), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n484), .A2(new_n715), .ZN(new_n716));
  AOI22_X1  g0516(.A1(new_n539), .A2(new_n303), .B1(new_n436), .B2(new_n534), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(new_n541), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n702), .A2(new_n718), .A3(new_n617), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n609), .B1(new_n716), .B2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n709), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(new_n628), .B2(KEYINPUT26), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n653), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n723), .A2(KEYINPUT95), .A3(KEYINPUT29), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n714), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n654), .B1(new_n620), .B2(new_n629), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT94), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OAI211_X1 g0528(.A(KEYINPUT94), .B(new_n654), .C1(new_n620), .C2(new_n629), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n728), .A2(new_n713), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n706), .B1(new_n725), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n677), .B1(new_n731), .B2(G1), .ZN(G364));
  AOI21_X1  g0532(.A(new_n228), .B1(G20), .B2(new_n429), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n436), .A2(G179), .A3(G200), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n229), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n206), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n229), .A2(new_n274), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G200), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n436), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(G50), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n229), .A2(G179), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n743), .A2(new_n436), .A3(G200), .ZN(new_n744));
  OAI22_X1  g0544(.A1(new_n741), .A2(new_n742), .B1(new_n744), .B2(new_n207), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n739), .A2(G190), .ZN(new_n746));
  AOI211_X1 g0546(.A(new_n737), .B(new_n745), .C1(G68), .C2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G190), .A2(G200), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n743), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G159), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n751), .A2(KEYINPUT32), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n743), .A2(G190), .A3(G200), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n751), .A2(KEYINPUT32), .B1(new_n754), .B2(G87), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n738), .A2(new_n748), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n264), .B1(new_n756), .B2(new_n267), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n738), .A2(G190), .A3(new_n303), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n757), .B1(new_n281), .B2(new_n759), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n747), .A2(new_n752), .A3(new_n755), .A4(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G322), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n758), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G311), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n370), .B1(new_n756), .B2(new_n764), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n763), .B(new_n765), .C1(G329), .C2(new_n750), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n740), .A2(G326), .ZN(new_n767));
  XNOR2_X1  g0567(.A(KEYINPUT33), .B(G317), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n746), .A2(new_n768), .B1(new_n754), .B2(G303), .ZN(new_n769));
  INV_X1    g0569(.A(new_n736), .ZN(new_n770));
  INV_X1    g0570(.A(new_n744), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n770), .A2(G294), .B1(new_n771), .B2(G283), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n766), .A2(new_n767), .A3(new_n769), .A4(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n734), .B1(new_n761), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G13), .A2(G33), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G20), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n733), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n247), .A2(G45), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n374), .A2(new_n375), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n670), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n780), .B(new_n782), .C1(G45), .C2(new_n233), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n264), .A2(new_n211), .ZN(new_n784));
  INV_X1    g0584(.A(G355), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n784), .A2(new_n785), .B1(G116), .B2(new_n211), .ZN(new_n786));
  XOR2_X1   g0586(.A(new_n786), .B(KEYINPUT96), .Z(new_n787));
  AOI21_X1  g0587(.A(new_n779), .B1(new_n783), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n673), .ZN(new_n789));
  INV_X1    g0589(.A(G13), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(G20), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n292), .B1(new_n791), .B2(G45), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n789), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n774), .A2(new_n788), .A3(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n777), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n796), .B1(new_n659), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n660), .A2(new_n795), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n659), .A2(G330), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(G396));
  AND2_X1   g0601(.A1(new_n653), .A2(new_n438), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n433), .B1(new_n802), .B2(new_n439), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n434), .A2(new_n654), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n728), .A2(new_n729), .A3(new_n806), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n654), .B(new_n805), .C1(new_n620), .C2(new_n629), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n706), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n794), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n807), .A2(new_n706), .A3(new_n808), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n756), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n759), .A2(G143), .B1(new_n813), .B2(G159), .ZN(new_n814));
  INV_X1    g0614(.A(G137), .ZN(new_n815));
  INV_X1    g0615(.A(G150), .ZN(new_n816));
  INV_X1    g0616(.A(new_n746), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n814), .B1(new_n741), .B2(new_n815), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT34), .ZN(new_n819));
  AND2_X1   g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(G132), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n781), .B1(new_n821), .B2(new_n749), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n744), .A2(new_n338), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(new_n281), .B2(new_n770), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n742), .B2(new_n753), .ZN(new_n825));
  NOR3_X1   g0625(.A1(new_n820), .A2(new_n822), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n819), .B2(new_n818), .ZN(new_n827));
  INV_X1    g0627(.A(G283), .ZN(new_n828));
  INV_X1    g0628(.A(G303), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n828), .A2(new_n817), .B1(new_n741), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(G107), .B2(new_n754), .ZN(new_n831));
  INV_X1    g0631(.A(G294), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n758), .A2(new_n832), .B1(new_n749), .B2(new_n764), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n264), .B(new_n833), .C1(G116), .C2(new_n813), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n737), .B1(G87), .B2(new_n771), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n831), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n734), .B1(new_n827), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n733), .A2(new_n775), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n795), .B(new_n837), .C1(new_n267), .C2(new_n838), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n839), .B(KEYINPUT97), .Z(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n776), .B2(new_n805), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n812), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(G384));
  INV_X1    g0643(.A(new_n547), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n844), .A2(KEYINPUT35), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(KEYINPUT35), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n845), .A2(G116), .A3(new_n230), .A4(new_n846), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT36), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n201), .A2(G68), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n849), .B(KEYINPUT98), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n267), .B1(new_n281), .B2(G68), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n850), .B1(new_n234), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n790), .A2(G1), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n568), .A2(new_n583), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n854), .A2(KEYINPUT30), .A3(new_n679), .A4(new_n530), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT30), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n680), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(KEYINPUT93), .B1(new_n690), .B2(new_n691), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n684), .A2(new_n686), .A3(new_n682), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(KEYINPUT102), .B1(new_n861), .B2(new_n695), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT102), .ZN(new_n863));
  INV_X1    g0663(.A(new_n695), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n693), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n862), .A2(new_n865), .B1(new_n694), .B2(KEYINPUT101), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT101), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT31), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n861), .B2(new_n654), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n536), .A2(new_n654), .A3(new_n542), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n607), .A2(new_n870), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n867), .A2(new_n869), .B1(new_n871), .B2(new_n492), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n866), .A2(new_n872), .A3(KEYINPUT103), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT103), .ZN(new_n874));
  OAI211_X1 g0674(.A(KEYINPUT101), .B(new_n868), .C1(new_n861), .C2(new_n654), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n863), .B1(new_n693), .B2(new_n864), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n860), .A2(new_n859), .ZN(new_n877));
  AOI211_X1 g0677(.A(KEYINPUT102), .B(new_n695), .C1(new_n877), .C2(new_n681), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n875), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n705), .B1(new_n694), .B2(KEYINPUT101), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n874), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n873), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n387), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n379), .A2(new_n277), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n369), .B1(new_n378), .B2(new_n338), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n380), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n883), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n887), .A2(new_n648), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n417), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n400), .B1(new_n887), .B2(new_n648), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n884), .A2(new_n886), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n387), .A2(new_n891), .B1(new_n412), .B2(new_n413), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT37), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT37), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n402), .A2(new_n647), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n410), .A2(new_n894), .A3(new_n400), .A4(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n889), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT38), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n889), .A2(new_n897), .A3(KEYINPUT38), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n361), .A2(new_n362), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n654), .A2(new_n349), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n903), .A2(new_n351), .A3(new_n905), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n356), .A2(new_n351), .A3(new_n358), .A4(new_n360), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n904), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT99), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n907), .A2(KEYINPUT99), .A3(new_n904), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n906), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n805), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n882), .A2(new_n902), .A3(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT40), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n895), .B1(new_n636), .B2(new_n401), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n895), .A2(new_n400), .ZN(new_n919));
  OAI21_X1  g0719(.A(KEYINPUT37), .B1(new_n919), .B2(new_n414), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n896), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n899), .B1(new_n918), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n916), .B1(new_n923), .B2(new_n901), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n924), .A2(new_n882), .A3(new_n914), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n917), .A2(new_n925), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n882), .A2(new_n442), .ZN(new_n927));
  OAI21_X1  g0727(.A(G330), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT104), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n928), .A2(new_n929), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n926), .A2(new_n927), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n725), .A2(new_n730), .A3(new_n442), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n640), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT100), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT39), .ZN(new_n937));
  AND3_X1   g0737(.A1(new_n889), .A2(new_n897), .A3(KEYINPUT38), .ZN(new_n938));
  INV_X1    g0738(.A(new_n895), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n417), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(KEYINPUT38), .B1(new_n940), .B2(new_n921), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n937), .B1(new_n938), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n900), .A2(KEYINPUT39), .A3(new_n901), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n361), .A2(new_n362), .A3(new_n654), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n942), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n636), .A2(new_n647), .ZN(new_n947));
  INV_X1    g0747(.A(new_n908), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n948), .A2(KEYINPUT99), .B1(new_n363), .B2(new_n905), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n910), .A2(new_n949), .B1(new_n808), .B2(new_n804), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n947), .B1(new_n902), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n946), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n936), .B(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n933), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n292), .B2(new_n791), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n933), .A2(new_n953), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n848), .B1(new_n852), .B2(new_n853), .C1(new_n955), .C2(new_n956), .ZN(G367));
  AND2_X1   g0757(.A1(new_n653), .A2(new_n621), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n958), .A2(new_n702), .B1(new_n622), .B2(new_n654), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n665), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT106), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n961), .A2(KEYINPUT42), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n565), .A2(new_n570), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n622), .B1(new_n964), .B2(new_n542), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n961), .A2(KEYINPUT42), .B1(new_n654), .B2(new_n965), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n654), .A2(new_n603), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n618), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n968), .A2(KEYINPUT105), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n968), .B(KEYINPUT105), .C1(new_n610), .C2(new_n967), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n962), .A2(new_n966), .B1(KEYINPUT43), .B2(new_n972), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n973), .B(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n664), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n959), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n975), .A2(new_n977), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n673), .B(KEYINPUT41), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n667), .A2(new_n959), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(KEYINPUT107), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT107), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n667), .A2(new_n983), .A3(new_n959), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(KEYINPUT45), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n667), .A2(new_n959), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT44), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n986), .A2(KEYINPUT45), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n991), .A2(new_n664), .A3(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n976), .B1(new_n990), .B2(new_n992), .ZN(new_n995));
  INV_X1    g0795(.A(new_n657), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n663), .B1(new_n996), .B2(new_n654), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n997), .A2(new_n665), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n660), .B(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n731), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n994), .A2(new_n995), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n980), .B1(new_n1002), .B2(new_n731), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n978), .B(new_n979), .C1(new_n1003), .C2(new_n793), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n778), .B1(new_n211), .B2(new_n421), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n782), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1006), .A2(new_n243), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n794), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n758), .A2(new_n816), .B1(new_n749), .B2(new_n815), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n370), .B(new_n1009), .C1(new_n202), .C2(new_n813), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n281), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1011), .A2(new_n753), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n736), .A2(new_n338), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1012), .B(new_n1013), .C1(G159), .C2(new_n746), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n740), .A2(G143), .B1(new_n771), .B2(G77), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1010), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G283), .A2(new_n813), .B1(new_n750), .B2(G317), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n829), .B2(new_n758), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n781), .B(new_n1018), .C1(G294), .C2(new_n746), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n736), .A2(new_n207), .B1(new_n744), .B2(new_n206), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(G311), .B2(new_n740), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT46), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n754), .A2(G116), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1019), .B(new_n1021), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1022), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT108), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1016), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  XOR2_X1   g0827(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n1028));
  XNOR2_X1  g0828(.A(new_n1027), .B(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1008), .B1(new_n1029), .B2(new_n733), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n972), .B2(new_n797), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1004), .A2(new_n1031), .ZN(G387));
  OR2_X1    g0832(.A1(new_n663), .A2(new_n797), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n784), .A2(new_n674), .B1(G107), .B2(new_n211), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n240), .A2(new_n256), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n419), .A2(new_n742), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT50), .Z(new_n1037));
  INV_X1    g0837(.A(new_n674), .ZN(new_n1038));
  AOI211_X1 g0838(.A(G45), .B(new_n1038), .C1(G68), .C2(G77), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1006), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1034), .B1(new_n1035), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n794), .B1(new_n1041), .B2(new_n779), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n781), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n741), .A2(new_n366), .B1(new_n753), .B2(new_n267), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1043), .B(new_n1044), .C1(G97), .C2(new_n771), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G68), .A2(new_n813), .B1(new_n750), .B2(G150), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n742), .B2(new_n758), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n593), .A2(new_n594), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1047), .B1(new_n1048), .B2(new_n770), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1045), .B(new_n1049), .C1(new_n386), .C2(new_n817), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n759), .A2(G317), .B1(new_n813), .B2(G303), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1051), .A2(KEYINPUT110), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(KEYINPUT110), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G311), .A2(new_n746), .B1(new_n740), .B2(G322), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT48), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n736), .A2(new_n828), .B1(new_n753), .B2(new_n832), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1057), .A2(KEYINPUT49), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n781), .B1(G326), .B2(new_n750), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1060), .B(new_n1061), .C1(new_n451), .C2(new_n744), .ZN(new_n1062));
  AOI21_X1  g0862(.A(KEYINPUT49), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1050), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1042), .B1(new_n1064), .B2(new_n733), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n999), .A2(new_n793), .B1(new_n1033), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1000), .A2(new_n789), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n999), .A2(new_n731), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1066), .B1(new_n1067), .B2(new_n1068), .ZN(G393));
  INV_X1    g0869(.A(KEYINPUT111), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n994), .A2(new_n995), .A3(new_n1070), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n991), .A2(KEYINPUT111), .A3(new_n664), .A4(new_n993), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n789), .B(new_n1002), .C1(new_n1073), .C2(new_n1001), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n959), .A2(new_n797), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n817), .A2(new_n829), .B1(new_n451), .B2(new_n736), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1076), .A2(KEYINPUT113), .B1(G294), .B2(new_n813), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(KEYINPUT113), .B2(new_n1076), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT114), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G317), .A2(new_n740), .B1(new_n759), .B2(G311), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT52), .Z(new_n1081));
  OAI221_X1 g0881(.A(new_n370), .B1(new_n749), .B2(new_n762), .C1(new_n207), .C2(new_n744), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(G283), .B2(new_n754), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1079), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G150), .A2(new_n740), .B1(new_n759), .B2(G159), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1085), .B(new_n1086), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n419), .A2(new_n813), .B1(new_n750), .B2(G143), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n736), .A2(new_n267), .ZN(new_n1089));
  INV_X1    g0889(.A(G87), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n338), .A2(new_n753), .B1(new_n744), .B2(new_n1090), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n1089), .B(new_n1091), .C1(new_n202), .C2(new_n746), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1087), .A2(new_n781), .A3(new_n1088), .A4(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n734), .B1(new_n1084), .B2(new_n1093), .ZN(new_n1094));
  OR2_X1    g0894(.A1(new_n1006), .A2(new_n250), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n779), .B1(G97), .B2(new_n670), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n795), .B(new_n1094), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1073), .A2(new_n793), .B1(new_n1075), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1074), .A2(new_n1098), .ZN(G390));
  NAND2_X1  g0899(.A1(new_n808), .A2(new_n804), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n912), .B1(new_n706), .B2(new_n805), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n678), .B1(new_n873), .B2(new_n881), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1102), .B1(new_n1103), .B2(new_n914), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n912), .B1(new_n1103), .B2(new_n805), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n706), .A2(new_n805), .A3(new_n912), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n723), .A2(new_n803), .B1(new_n434), .B2(new_n654), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n1101), .A2(new_n1104), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1103), .A2(new_n442), .ZN(new_n1110));
  AND3_X1   g0910(.A1(new_n1110), .A2(new_n640), .A3(new_n934), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n882), .A2(G330), .A3(new_n914), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1100), .A2(new_n912), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n942), .A2(new_n943), .B1(new_n1114), .B2(new_n944), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n723), .A2(new_n803), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1116), .A2(new_n804), .B1(new_n910), .B2(new_n949), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n944), .B1(new_n938), .B2(new_n941), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1113), .B1(new_n1115), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(KEYINPUT38), .B1(new_n889), .B2(new_n897), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n938), .A2(new_n1121), .A3(new_n937), .ZN(new_n1122));
  AOI21_X1  g0922(.A(KEYINPUT39), .B1(new_n923), .B2(new_n901), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n1122), .A2(new_n1123), .B1(new_n945), .B2(new_n950), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n912), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n944), .B1(new_n938), .B2(new_n941), .C1(new_n1107), .C2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1124), .A2(new_n1106), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1120), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1112), .A2(new_n1128), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1109), .A2(new_n1111), .A3(new_n1127), .A4(new_n1120), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1129), .A2(new_n789), .A3(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1120), .A2(new_n1127), .A3(new_n793), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n775), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n838), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n794), .B1(new_n1134), .B2(new_n282), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n758), .A2(new_n451), .B1(new_n749), .B2(new_n832), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n264), .B(new_n1136), .C1(G97), .C2(new_n813), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n746), .A2(G107), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1089), .B1(G283), .B2(new_n740), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n823), .B1(G87), .B2(new_n754), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .A4(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(KEYINPUT54), .B(G143), .ZN(new_n1142));
  INV_X1    g0942(.A(G125), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n756), .A2(new_n1142), .B1(new_n749), .B2(new_n1143), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n370), .B(new_n1144), .C1(G132), .C2(new_n759), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(G128), .A2(new_n740), .B1(new_n202), .B2(new_n771), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(G159), .A2(new_n770), .B1(new_n746), .B2(G137), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n753), .A2(new_n816), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1149), .B(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1141), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1135), .B1(new_n1152), .B2(new_n733), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1133), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1132), .A2(new_n1154), .ZN(new_n1155));
  AND2_X1   g0955(.A1(new_n1155), .A2(KEYINPUT116), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1155), .A2(KEYINPUT116), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1131), .B1(new_n1156), .B2(new_n1157), .ZN(G378));
  AOI21_X1  g0958(.A(new_n913), .B1(new_n881), .B2(new_n873), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n678), .B1(new_n1159), .B2(new_n924), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n299), .A2(new_n647), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n312), .A2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n312), .A2(new_n1162), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  OR3_X1    g0966(.A1(new_n1163), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1166), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n917), .A2(new_n1160), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1169), .B1(new_n917), .B2(new_n1160), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n952), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n925), .A2(G330), .ZN(new_n1174));
  AOI21_X1  g0974(.A(KEYINPUT40), .B1(new_n1159), .B2(new_n902), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1173), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n952), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n917), .A2(new_n1160), .A3(new_n1169), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1172), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n793), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1173), .A2(new_n775), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n794), .B1(new_n1134), .B2(new_n202), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n1143), .A2(new_n741), .B1(new_n817), .B2(new_n821), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n759), .A2(G128), .B1(new_n813), .B2(G137), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n753), .B2(new_n1142), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1184), .B(new_n1186), .C1(G150), .C2(new_n770), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  OR2_X1    g0988(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n317), .A2(new_n255), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT117), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n744), .A2(new_n366), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(KEYINPUT118), .B(G124), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1192), .B(new_n1193), .C1(new_n750), .C2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1189), .A2(new_n1190), .A3(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1011), .A2(new_n744), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n206), .A2(new_n817), .B1(new_n741), .B2(new_n451), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1197), .B(new_n1198), .C1(G77), .C2(new_n754), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n758), .A2(new_n207), .B1(new_n749), .B2(new_n828), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1013), .B(new_n1200), .C1(new_n1048), .C2(new_n813), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1199), .A2(new_n255), .A3(new_n1201), .A4(new_n1043), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT58), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n742), .B(new_n1192), .C1(new_n781), .C2(G41), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1196), .A2(new_n1204), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1183), .B1(new_n1207), .B2(new_n733), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1182), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1181), .A2(new_n1209), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1179), .A2(new_n1172), .B1(new_n1130), .B2(new_n1111), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n673), .B1(new_n1211), .B2(KEYINPUT57), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n882), .A2(G330), .A3(new_n914), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1102), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1101), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n882), .A2(G330), .A3(new_n805), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1108), .B1(new_n1216), .B2(new_n1125), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1111), .B1(new_n1128), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1180), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT57), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1210), .B1(new_n1212), .B2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(G375));
  NAND2_X1  g1024(.A1(new_n1125), .A2(new_n775), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n794), .B1(new_n1134), .B2(G68), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n741), .A2(new_n821), .B1(new_n742), .B2(new_n736), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n817), .A2(new_n1142), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(new_n1227), .A2(new_n1228), .A3(new_n1197), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n754), .A2(G159), .B1(new_n750), .B2(G128), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT120), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n759), .A2(G137), .B1(new_n813), .B2(G150), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1229), .A2(new_n1231), .A3(new_n781), .A4(new_n1232), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1048), .A2(new_n770), .B1(G283), .B2(new_n759), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1234), .B(KEYINPUT119), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n451), .A2(new_n817), .B1(new_n741), .B2(new_n832), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n370), .B1(new_n749), .B2(new_n829), .C1(new_n207), .C2(new_n756), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n267), .A2(new_n744), .B1(new_n753), .B2(new_n206), .ZN(new_n1238));
  OR3_X1    g1038(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1233), .B1(new_n1235), .B2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1226), .B1(new_n1240), .B2(new_n733), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n1109), .A2(new_n793), .B1(new_n1225), .B2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n980), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1112), .A2(new_n1243), .ZN(new_n1244));
  NOR3_X1   g1044(.A1(new_n1111), .A2(new_n1215), .A3(new_n1217), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1242), .B1(new_n1244), .B2(new_n1245), .ZN(G381));
  OR4_X1    g1046(.A1(G396), .A2(G381), .A3(G384), .A4(G393), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1131), .A2(new_n1132), .A3(new_n1154), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1247), .A2(G390), .A3(new_n1249), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1250), .A2(new_n1004), .A3(new_n1031), .A4(new_n1223), .ZN(G407));
  NAND2_X1  g1051(.A1(new_n649), .A2(G213), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1223), .A2(new_n1248), .A3(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(G407), .A2(G213), .A3(new_n1254), .ZN(G409));
  INV_X1    g1055(.A(KEYINPUT126), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1253), .A2(G2897), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT123), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1245), .B1(KEYINPUT60), .B2(new_n1112), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1217), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1100), .B1(new_n1113), .B2(new_n1102), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1110), .A2(new_n640), .A3(new_n934), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1262), .A2(new_n1263), .A3(KEYINPUT60), .A4(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n789), .ZN(new_n1266));
  OAI211_X1 g1066(.A(KEYINPUT122), .B(new_n1242), .C1(new_n1261), .C2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n842), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1266), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1218), .A2(new_n1264), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1264), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT60), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1270), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1269), .A2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(KEYINPUT122), .B1(new_n1274), .B2(new_n1242), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1268), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1242), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(new_n1269), .B2(new_n1273), .ZN(new_n1278));
  NOR3_X1   g1078(.A1(new_n1278), .A2(KEYINPUT122), .A3(new_n842), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1260), .B1(new_n1276), .B2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(G384), .B1(new_n1278), .B2(KEYINPUT122), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT122), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1261), .A2(new_n1266), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1282), .B1(new_n1283), .B2(new_n1277), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1281), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1268), .A2(new_n1275), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(new_n1257), .B(new_n1258), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1285), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1280), .A2(new_n1288), .ZN(new_n1289));
  NOR3_X1   g1089(.A1(new_n1170), .A2(new_n1171), .A3(new_n952), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1177), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1219), .B(new_n1243), .C1(new_n1290), .C2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(KEYINPUT121), .ZN(new_n1293));
  AOI22_X1  g1093(.A1(new_n1180), .A2(new_n793), .B1(new_n1182), .B2(new_n1208), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT121), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1180), .A2(new_n1295), .A3(new_n1243), .A4(new_n1219), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1293), .A2(new_n1294), .A3(new_n1296), .ZN(new_n1297));
  AOI22_X1  g1097(.A1(new_n1223), .A2(G378), .B1(new_n1248), .B2(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(KEYINPUT125), .B1(new_n1298), .B2(new_n1253), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1297), .A2(new_n1248), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1180), .A2(KEYINPUT57), .A3(new_n1219), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n789), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1211), .A2(KEYINPUT57), .ZN(new_n1303));
  OAI211_X1 g1103(.A(G378), .B(new_n1294), .C1(new_n1302), .C2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1300), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT125), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1305), .A2(new_n1306), .A3(new_n1252), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1289), .B1(new_n1299), .B2(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1256), .B1(new_n1308), .B2(KEYINPUT61), .ZN(new_n1309));
  AND3_X1   g1109(.A1(new_n1285), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1259), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1306), .B1(new_n1305), .B2(new_n1252), .ZN(new_n1313));
  AOI211_X1 g1113(.A(KEYINPUT125), .B(new_n1253), .C1(new_n1300), .C2(new_n1304), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1312), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT61), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1315), .A2(KEYINPUT126), .A3(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1305), .A2(new_n1318), .A3(new_n1252), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1319), .A2(KEYINPUT62), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1299), .A2(new_n1318), .A3(new_n1307), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1320), .B1(new_n1321), .B2(KEYINPUT62), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1309), .A2(new_n1317), .A3(new_n1322), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(G387), .A2(new_n1074), .A3(new_n1098), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(G390), .A2(new_n1004), .A3(new_n1031), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  XOR2_X1   g1126(.A(G393), .B(G396), .Z(new_n1327));
  INV_X1    g1127(.A(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1326), .A2(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1324), .A2(new_n1327), .A3(new_n1325), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1323), .A2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT63), .ZN(new_n1333));
  AND2_X1   g1133(.A1(new_n1319), .A2(new_n1333), .ZN(new_n1334));
  NOR3_X1   g1134(.A1(new_n1331), .A2(new_n1334), .A3(KEYINPUT61), .ZN(new_n1335));
  OAI211_X1 g1135(.A(new_n1280), .B(new_n1288), .C1(new_n1298), .C2(new_n1253), .ZN(new_n1336));
  XNOR2_X1  g1136(.A(new_n1336), .B(KEYINPUT124), .ZN(new_n1337));
  OAI211_X1 g1137(.A(new_n1335), .B(new_n1337), .C1(new_n1333), .C2(new_n1321), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1332), .A2(new_n1338), .ZN(G405));
  INV_X1    g1139(.A(new_n1304), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1340), .B1(G375), .B2(new_n1248), .ZN(new_n1341));
  OR2_X1    g1141(.A1(new_n1341), .A2(KEYINPUT127), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1341), .A2(KEYINPUT127), .ZN(new_n1343));
  NAND4_X1  g1143(.A1(new_n1342), .A2(new_n1286), .A3(new_n1285), .A4(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1331), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1341), .A2(KEYINPUT127), .A3(new_n1318), .ZN(new_n1346));
  AND3_X1   g1146(.A1(new_n1344), .A2(new_n1345), .A3(new_n1346), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1345), .B1(new_n1344), .B2(new_n1346), .ZN(new_n1348));
  NOR2_X1   g1148(.A1(new_n1347), .A2(new_n1348), .ZN(G402));
endmodule


