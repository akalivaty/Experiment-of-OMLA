//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1 1 0 0 0 1 1 1 1 0 1 0 1 1 0 0 1 1 1 0 1 0 1 0 0 1 1 1 1 1 0 1 1 0 0 0 1 0 1 1 1 1 1 0 1 0 0 1 0 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n434, new_n437, new_n448, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n555, new_n557, new_n558, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n612, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1165, new_n1166;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(new_n434));
  INV_X1    g009(.A(new_n434), .ZN(G218));
  XOR2_X1   g010(.A(KEYINPUT65), .B(G132), .Z(G219));
  XOR2_X1   g011(.A(KEYINPUT0), .B(G82), .Z(new_n437));
  XNOR2_X1  g012(.A(new_n437), .B(KEYINPUT66), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  NAND2_X1  g032(.A1(KEYINPUT67), .A2(G2104), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g035(.A1(KEYINPUT67), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G137), .ZN(new_n463));
  NAND2_X1  g038(.A1(G101), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n465), .A2(new_n470), .ZN(G160));
  AOI21_X1  g046(.A(G2105), .B1(new_n460), .B2(new_n461), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G136), .ZN(new_n473));
  NOR2_X1   g048(.A1(G100), .A2(G2105), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n474), .B(KEYINPUT68), .ZN(new_n475));
  OAI21_X1  g050(.A(G2104), .B1(new_n466), .B2(G112), .ZN(new_n476));
  INV_X1    g051(.A(G124), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n462), .A2(G2105), .ZN(new_n478));
  OAI221_X1 g053(.A(new_n473), .B1(new_n475), .B2(new_n476), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G162));
  NAND3_X1  g055(.A1(new_n467), .A2(G138), .A3(new_n466), .ZN(new_n481));
  AND3_X1   g056(.A1(KEYINPUT67), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n482));
  AOI21_X1  g057(.A(KEYINPUT3), .B1(KEYINPUT67), .B2(G2104), .ZN(new_n483));
  OAI21_X1  g058(.A(G126), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(G114), .A2(G2104), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n466), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n481), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI211_X1 g063(.A(KEYINPUT4), .B(G138), .C1(new_n482), .C2(new_n483), .ZN(new_n489));
  NAND2_X1  g064(.A1(G102), .A2(G2104), .ZN(new_n490));
  AOI21_X1  g065(.A(G2105), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G164));
  INV_X1    g069(.A(G543), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT5), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT5), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G543), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G62), .ZN(new_n500));
  OR3_X1    g075(.A1(new_n499), .A2(KEYINPUT70), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(G75), .A2(G543), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT70), .B1(new_n499), .B2(new_n500), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT69), .B(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT69), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT69), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G651), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n507), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n508), .A2(KEYINPUT6), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(G50), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n515), .B1(new_n499), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n506), .A2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  INV_X1    g095(.A(new_n499), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n522));
  OAI21_X1  g097(.A(KEYINPUT71), .B1(new_n512), .B2(new_n513), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT71), .ZN(new_n524));
  INV_X1    g099(.A(new_n513), .ZN(new_n525));
  OAI211_X1 g100(.A(new_n524), .B(new_n525), .C1(new_n505), .C2(new_n507), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n523), .A2(G543), .A3(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G51), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n522), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT72), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n529), .B(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  INV_X1    g108(.A(G89), .ZN(new_n534));
  NOR3_X1   g109(.A1(new_n512), .A2(new_n513), .A3(new_n499), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  OAI211_X1 g111(.A(new_n531), .B(new_n533), .C1(new_n534), .C2(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  AOI22_X1  g113(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  INV_X1    g114(.A(new_n505), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT73), .ZN(new_n542));
  AND3_X1   g117(.A1(new_n523), .A2(G543), .A3(new_n526), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G52), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n535), .A2(G90), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n542), .A2(new_n544), .A3(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  NAND2_X1  g122(.A1(new_n543), .A2(G43), .ZN(new_n548));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G56), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n499), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n535), .A2(G81), .B1(new_n505), .B2(new_n551), .ZN(new_n552));
  AND2_X1   g127(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  AND3_X1   g129(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G36), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n555), .A2(new_n558), .ZN(G188));
  NAND3_X1  g134(.A1(new_n543), .A2(KEYINPUT9), .A3(G53), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n499), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n535), .A2(G91), .B1(G651), .B2(new_n563), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n523), .A2(G53), .A3(G543), .A4(new_n526), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n560), .A2(new_n564), .A3(new_n567), .ZN(G299));
  INV_X1    g143(.A(KEYINPUT74), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n543), .A2(new_n569), .A3(G49), .ZN(new_n570));
  INV_X1    g145(.A(G74), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n508), .B1(new_n499), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n572), .B1(new_n535), .B2(G87), .ZN(new_n573));
  INV_X1    g148(.A(G49), .ZN(new_n574));
  OAI21_X1  g149(.A(KEYINPUT74), .B1(new_n527), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n570), .A2(new_n573), .A3(new_n575), .ZN(G288));
  NAND2_X1  g151(.A1(new_n535), .A2(G86), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n514), .A2(G48), .A3(G543), .ZN(new_n578));
  INV_X1    g153(.A(G73), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT75), .B1(new_n579), .B2(new_n495), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT75), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n581), .A2(G73), .A3(G543), .ZN(new_n582));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n580), .B(new_n582), .C1(new_n499), .C2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(new_n505), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n577), .A2(new_n578), .A3(new_n585), .ZN(G305));
  AOI22_X1  g161(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n587), .A2(new_n540), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n535), .A2(G85), .ZN(new_n589));
  INV_X1    g164(.A(G47), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n527), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT76), .ZN(new_n592));
  AND2_X1   g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n591), .A2(new_n592), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n588), .B1(new_n593), .B2(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(G301), .A2(G868), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n535), .A2(G92), .ZN(new_n597));
  XOR2_X1   g172(.A(new_n597), .B(KEYINPUT10), .Z(new_n598));
  NAND2_X1  g173(.A1(new_n543), .A2(G54), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  XOR2_X1   g175(.A(KEYINPUT77), .B(G66), .Z(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(new_n499), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G651), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n598), .A2(new_n599), .A3(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n596), .B1(new_n605), .B2(G868), .ZN(G284));
  OAI21_X1  g181(.A(new_n596), .B1(new_n605), .B2(G868), .ZN(G321));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(G299), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G168), .B2(new_n608), .ZN(G297));
  XNOR2_X1  g185(.A(G297), .B(KEYINPUT78), .ZN(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n605), .B1(new_n612), .B2(G860), .ZN(G148));
  NAND2_X1  g188(.A1(new_n605), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G868), .B2(new_n553), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g192(.A(G123), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n478), .A2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT79), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n472), .A2(G135), .ZN(new_n622));
  NOR2_X1   g197(.A1(G99), .A2(G2105), .ZN(new_n623));
  OAI21_X1  g198(.A(G2104), .B1(new_n466), .B2(G111), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n621), .B(new_n622), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(G2096), .Z(new_n626));
  NAND3_X1  g201(.A1(new_n466), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT12), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2100), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n626), .A2(new_n630), .ZN(G156));
  XOR2_X1   g206(.A(KEYINPUT82), .B(G2438), .Z(new_n632));
  XNOR2_X1  g207(.A(G2427), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(KEYINPUT15), .B(G2435), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT81), .B(KEYINPUT14), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2451), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2454), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n638), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2443), .B(G2446), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G1341), .B(G1348), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(G14), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(KEYINPUT83), .ZN(new_n648));
  INV_X1    g223(.A(KEYINPUT83), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n646), .A2(new_n649), .A3(G14), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(G401));
  XNOR2_X1  g227(.A(G2084), .B(G2090), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT84), .ZN(new_n654));
  XOR2_X1   g229(.A(G2067), .B(G2678), .Z(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2072), .B(G2078), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT17), .Z(new_n658));
  AOI21_X1  g233(.A(new_n658), .B1(new_n654), .B2(new_n655), .ZN(new_n659));
  INV_X1    g234(.A(new_n655), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n660), .A2(new_n657), .ZN(new_n661));
  AOI211_X1 g236(.A(new_n656), .B(new_n659), .C1(new_n654), .C2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n656), .A2(new_n657), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT18), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2096), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(G2100), .Z(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(G227));
  XNOR2_X1  g243(.A(G1961), .B(G1966), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT85), .ZN(new_n670));
  XOR2_X1   g245(.A(G1956), .B(G2474), .Z(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n672), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(KEYINPUT87), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n673), .A2(new_n676), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(G1986), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1991), .B(G1996), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n685), .B(new_n686), .Z(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT22), .B(G1981), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(G229));
  NOR2_X1   g265(.A1(G16), .A2(G21), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(G168), .B2(G16), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G1966), .ZN(new_n693));
  NOR2_X1   g268(.A1(G4), .A2(G16), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n605), .B2(G16), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G1348), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(G5), .A2(G16), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(G171), .B2(G16), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G1961), .ZN(new_n701));
  OAI22_X1  g276(.A1(new_n700), .A2(new_n701), .B1(new_n695), .B2(G1348), .ZN(new_n702));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G26), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n472), .A2(G140), .ZN(new_n705));
  NOR2_X1   g280(.A1(G104), .A2(G2105), .ZN(new_n706));
  OAI21_X1  g281(.A(G2104), .B1(new_n466), .B2(G116), .ZN(new_n707));
  INV_X1    g282(.A(G128), .ZN(new_n708));
  OAI221_X1 g283(.A(new_n705), .B1(new_n706), .B2(new_n707), .C1(new_n708), .C2(new_n478), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT94), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n704), .B1(new_n710), .B2(new_n703), .ZN(new_n711));
  MUX2_X1   g286(.A(new_n704), .B(new_n711), .S(KEYINPUT28), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G2067), .ZN(new_n713));
  NOR3_X1   g288(.A1(new_n697), .A2(new_n702), .A3(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n692), .A2(G1966), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT31), .B(G11), .Z(new_n716));
  NAND2_X1  g291(.A1(new_n703), .A2(G35), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G162), .B2(new_n703), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT29), .Z(new_n719));
  INV_X1    g294(.A(G2090), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n716), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT97), .B(KEYINPUT24), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G34), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n723), .A2(G29), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G160), .B2(G29), .ZN(new_n725));
  INV_X1    g300(.A(G2084), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n625), .A2(new_n703), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT30), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n729), .A2(G28), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(G28), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n730), .A2(new_n731), .A3(new_n703), .ZN(new_n732));
  NAND4_X1  g307(.A1(new_n721), .A2(new_n727), .A3(new_n728), .A4(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n719), .A2(new_n720), .ZN(new_n734));
  NOR3_X1   g309(.A1(new_n715), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(G27), .A2(G29), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G164), .B2(G29), .ZN(new_n737));
  INV_X1    g312(.A(G2078), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G16), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G19), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n553), .B2(new_n740), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT93), .B(G1341), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n701), .B2(new_n700), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n714), .A2(new_n735), .A3(new_n739), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n740), .A2(G23), .ZN(new_n747));
  INV_X1    g322(.A(G288), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(new_n740), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT33), .B(G1976), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT91), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n749), .B(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n740), .A2(G22), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G166), .B2(new_n740), .ZN(new_n754));
  INV_X1    g329(.A(G1971), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  MUX2_X1   g332(.A(G6), .B(G305), .S(G16), .Z(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT90), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT32), .B(G1981), .Z(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT92), .ZN(new_n762));
  OAI22_X1  g337(.A1(new_n757), .A2(new_n761), .B1(new_n762), .B2(KEYINPUT34), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(KEYINPUT34), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g340(.A(G290), .B(KEYINPUT88), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(G16), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n740), .A2(G24), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT89), .B(G1986), .Z(new_n769));
  AND3_X1   g344(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n769), .B1(new_n767), .B2(new_n768), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n703), .A2(G25), .ZN(new_n772));
  INV_X1    g347(.A(new_n478), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G119), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n472), .A2(G131), .ZN(new_n775));
  OR2_X1    g350(.A1(G95), .A2(G2105), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n776), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n774), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n772), .B1(new_n779), .B2(new_n703), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT35), .B(G1991), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n770), .A2(new_n771), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n763), .A2(new_n764), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n765), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(KEYINPUT36), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT36), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n765), .A2(new_n787), .A3(new_n783), .A4(new_n784), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n746), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(G29), .A2(G33), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT25), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n793), .A2(new_n466), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT95), .Z(new_n795));
  AOI211_X1 g370(.A(new_n792), .B(new_n795), .C1(G139), .C2(new_n472), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n790), .B1(new_n796), .B2(G29), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT96), .B(G2072), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(G29), .A2(G32), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n773), .A2(G129), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n466), .A2(G105), .A3(G2104), .ZN(new_n802));
  NAND3_X1  g377(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT26), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n472), .A2(G141), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n801), .A2(new_n802), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT98), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n800), .B1(new_n808), .B2(G29), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT27), .B(G1996), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n740), .A2(KEYINPUT23), .A3(G20), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT23), .ZN(new_n813));
  INV_X1    g388(.A(G20), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(G16), .ZN(new_n815));
  INV_X1    g390(.A(G299), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n812), .B(new_n815), .C1(new_n816), .C2(new_n740), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT99), .B(G1956), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n789), .A2(new_n799), .A3(new_n811), .A4(new_n819), .ZN(G150));
  INV_X1    g395(.A(G150), .ZN(G311));
  NAND2_X1  g396(.A1(new_n535), .A2(G93), .ZN(new_n822));
  AOI22_X1  g397(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n823));
  INV_X1    g398(.A(G55), .ZN(new_n824));
  OAI221_X1 g399(.A(new_n822), .B1(new_n540), .B2(new_n823), .C1(new_n527), .C2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(G860), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT37), .Z(new_n827));
  OR2_X1    g402(.A1(new_n553), .A2(new_n825), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n553), .A2(new_n825), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XOR2_X1   g405(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n604), .A2(new_n612), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n827), .B1(new_n834), .B2(G860), .ZN(G145));
  INV_X1    g410(.A(new_n481), .ZN(new_n836));
  INV_X1    g411(.A(G126), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(new_n460), .B2(new_n461), .ZN(new_n838));
  INV_X1    g413(.A(new_n485), .ZN(new_n839));
  OAI21_X1  g414(.A(G2105), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n836), .B1(new_n840), .B2(KEYINPUT4), .ZN(new_n841));
  NOR3_X1   g416(.A1(new_n841), .A2(KEYINPUT100), .A3(new_n491), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT100), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(new_n488), .B2(new_n492), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n709), .B(KEYINPUT94), .Z(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n842), .A2(new_n844), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(new_n710), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n806), .B(KEYINPUT102), .Z(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n852), .A2(new_n796), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n850), .A2(KEYINPUT101), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT101), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n847), .A2(new_n855), .A3(new_n849), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(new_n808), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n854), .A2(new_n807), .A3(new_n856), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n858), .A2(new_n796), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n853), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n472), .A2(G142), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(KEYINPUT103), .Z(new_n863));
  INV_X1    g438(.A(G130), .ZN(new_n864));
  NOR2_X1   g439(.A1(G106), .A2(G2105), .ZN(new_n865));
  OAI21_X1  g440(.A(G2104), .B1(new_n466), .B2(G118), .ZN(new_n866));
  OAI22_X1  g441(.A1(new_n478), .A2(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n628), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n779), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n861), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n870), .B(KEYINPUT104), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n872), .A2(new_n860), .A3(new_n853), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n625), .B(G160), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(G162), .ZN(new_n876));
  OR3_X1    g451(.A1(new_n871), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  XOR2_X1   g452(.A(KEYINPUT105), .B(G37), .Z(new_n878));
  INV_X1    g453(.A(new_n872), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(new_n861), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(new_n873), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n878), .B1(new_n881), .B2(new_n876), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n877), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g459(.A1(new_n605), .A2(new_n816), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n604), .A2(G299), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT41), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT106), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT41), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n885), .A2(new_n890), .A3(new_n886), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n887), .A2(KEYINPUT106), .A3(KEYINPUT41), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n828), .A2(new_n829), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(new_n614), .ZN(new_n896));
  MUX2_X1   g471(.A(new_n894), .B(new_n887), .S(new_n896), .Z(new_n897));
  OR2_X1    g472(.A1(new_n897), .A2(KEYINPUT42), .ZN(new_n898));
  XNOR2_X1  g473(.A(G290), .B(G303), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(G288), .ZN(new_n900));
  XNOR2_X1  g475(.A(G290), .B(G166), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(new_n748), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  XOR2_X1   g478(.A(G305), .B(KEYINPUT107), .Z(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n900), .A2(new_n902), .A3(new_n904), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n897), .A2(KEYINPUT42), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n898), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n909), .B1(new_n898), .B2(new_n910), .ZN(new_n912));
  OAI21_X1  g487(.A(G868), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n825), .A2(new_n608), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(G295));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n914), .ZN(G331));
  NAND2_X1  g491(.A1(G168), .A2(new_n830), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n895), .A2(G286), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(new_n918), .A3(G171), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(G171), .B1(new_n917), .B2(new_n918), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n892), .B(new_n893), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n921), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n923), .A2(new_n919), .A3(new_n886), .A4(new_n885), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n909), .ZN(new_n926));
  INV_X1    g501(.A(G37), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n922), .A2(new_n924), .A3(new_n908), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(KEYINPUT109), .A3(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT109), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n932), .B1(new_n933), .B2(KEYINPUT43), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n920), .A2(new_n921), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n888), .A2(new_n891), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n924), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(new_n909), .ZN(new_n938));
  INV_X1    g513(.A(new_n878), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(new_n939), .A3(new_n928), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(KEYINPUT43), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n931), .A2(new_n934), .A3(KEYINPUT44), .A4(new_n941), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n938), .A2(new_n930), .A3(new_n939), .A4(new_n928), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n943), .B1(new_n929), .B2(new_n930), .ZN(new_n944));
  XNOR2_X1  g519(.A(KEYINPUT108), .B(KEYINPUT44), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n942), .A2(new_n946), .ZN(G397));
  NAND2_X1  g522(.A1(G160), .A2(G40), .ZN(new_n948));
  INV_X1    g523(.A(G1384), .ZN(new_n949));
  AOI211_X1 g524(.A(KEYINPUT45), .B(new_n948), .C1(new_n845), .C2(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n710), .B(G2067), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n806), .A2(G1996), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n951), .B(new_n952), .C1(G1996), .C2(new_n807), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n778), .A2(new_n781), .ZN(new_n954));
  OR2_X1    g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n778), .A2(new_n781), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n950), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(G1986), .ZN(new_n958));
  INV_X1    g533(.A(G290), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n950), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n950), .A2(G1986), .A3(G290), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  XOR2_X1   g537(.A(new_n962), .B(KEYINPUT110), .Z(new_n963));
  INV_X1    g538(.A(G8), .ZN(new_n964));
  AOI21_X1  g539(.A(G1384), .B1(new_n488), .B2(new_n492), .ZN(new_n965));
  INV_X1    g540(.A(G40), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n465), .A2(new_n470), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n964), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G1976), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n968), .B1(G288), .B2(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n970), .A2(KEYINPUT52), .ZN(new_n971));
  NAND2_X1  g546(.A1(G288), .A2(new_n969), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(G305), .A2(G1981), .ZN(new_n974));
  INV_X1    g549(.A(G1981), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n577), .A2(new_n578), .A3(new_n975), .A4(new_n585), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT114), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n976), .A2(new_n977), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n974), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT49), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI211_X1 g557(.A(KEYINPUT49), .B(new_n974), .C1(new_n978), .C2(new_n979), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n982), .A2(new_n968), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT113), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n985), .B1(new_n970), .B2(KEYINPUT52), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n970), .A2(new_n985), .A3(KEYINPUT52), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n973), .B(new_n984), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(G303), .A2(G8), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT112), .ZN(new_n991));
  NOR3_X1   g566(.A1(new_n990), .A2(new_n991), .A3(KEYINPUT55), .ZN(new_n992));
  XNOR2_X1  g567(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n992), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  OAI211_X1 g569(.A(KEYINPUT45), .B(new_n949), .C1(new_n842), .C2(new_n844), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n949), .B1(new_n841), .B2(new_n491), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n948), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT111), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT111), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n995), .A2(new_n1001), .A3(new_n998), .ZN(new_n1002));
  AOI21_X1  g577(.A(G1971), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n967), .B1(new_n965), .B2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n996), .A2(KEYINPUT50), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1008), .A2(G2090), .ZN(new_n1009));
  OAI211_X1 g584(.A(G8), .B(new_n994), .C1(new_n1003), .C2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1002), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1001), .B1(new_n995), .B2(new_n998), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n755), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n493), .A2(new_n1004), .A3(new_n949), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT116), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n948), .B1(new_n996), .B2(KEYINPUT50), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n965), .A2(new_n1017), .A3(new_n1004), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1015), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  OR2_X1    g594(.A1(new_n1019), .A2(G2090), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n964), .B1(new_n1013), .B2(new_n1020), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n989), .B(new_n1010), .C1(new_n1021), .C2(new_n994), .ZN(new_n1022));
  XOR2_X1   g597(.A(new_n1022), .B(KEYINPUT125), .Z(new_n1023));
  INV_X1    g598(.A(KEYINPUT117), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1024), .B1(new_n1007), .B2(new_n726), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1016), .A2(new_n1024), .A3(new_n726), .A4(new_n1014), .ZN(new_n1026));
  INV_X1    g601(.A(G1966), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n967), .B1(new_n965), .B2(KEYINPUT45), .ZN(new_n1028));
  AOI211_X1 g603(.A(new_n997), .B(G1384), .C1(new_n488), .C2(new_n492), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1026), .A2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(G8), .B1(new_n1025), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT51), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1033), .A2(KEYINPUT121), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(G286), .A2(G8), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1032), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1033), .A2(KEYINPUT121), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1016), .A2(new_n726), .A3(new_n1014), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT117), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1040), .A2(new_n1030), .A3(new_n1026), .ZN(new_n1041));
  OAI211_X1 g616(.A(G8), .B(new_n1034), .C1(new_n1041), .C2(G286), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1037), .A2(new_n1038), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1032), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(G286), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1043), .A2(KEYINPUT122), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT122), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT62), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT122), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT62), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1043), .A2(KEYINPUT122), .A3(new_n1045), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1000), .A2(new_n738), .A3(new_n1002), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1008), .A2(new_n701), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1029), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n998), .A2(new_n1059), .A3(new_n738), .ZN(new_n1060));
  OR2_X1    g635(.A1(new_n1060), .A2(KEYINPUT124), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(KEYINPUT124), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(KEYINPUT53), .A3(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1057), .A2(new_n1058), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(G171), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1048), .A2(new_n1054), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n845), .A2(new_n949), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1056), .B1(new_n1068), .B2(new_n997), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1069), .A2(new_n738), .A3(new_n967), .A4(new_n995), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1057), .A2(new_n1070), .A3(G301), .A4(new_n1058), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1065), .A2(new_n1071), .ZN(new_n1072));
  XOR2_X1   g647(.A(KEYINPUT123), .B(KEYINPUT54), .Z(new_n1073));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1057), .A2(new_n1058), .A3(new_n1070), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1074), .B1(new_n1075), .B2(G171), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1057), .A2(new_n1063), .A3(G301), .A4(new_n1058), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1072), .A2(new_n1073), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G1956), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1019), .A2(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g655(.A(KEYINPUT56), .B(G2072), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n995), .A2(new_n998), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n1084));
  NOR2_X1   g659(.A1(G299), .A2(KEYINPUT119), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT119), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n565), .B(KEYINPUT9), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1086), .B1(new_n1087), .B2(new_n564), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1084), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT120), .ZN(new_n1090));
  NAND2_X1  g665(.A1(G299), .A2(KEYINPUT119), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1087), .A2(new_n1086), .A3(new_n564), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1091), .A2(new_n1092), .A3(KEYINPUT57), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1089), .A2(new_n1090), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1090), .B1(new_n1089), .B2(new_n1093), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1083), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1089), .A2(new_n1080), .A3(new_n1082), .A4(new_n1093), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1096), .A2(KEYINPUT61), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT60), .ZN(new_n1099));
  AOI21_X1  g674(.A(G1348), .B1(new_n1016), .B2(new_n1014), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n965), .A2(new_n967), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1101), .A2(G2067), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1099), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  OR2_X1    g678(.A1(new_n1101), .A2(G2067), .ZN(new_n1104));
  OAI211_X1 g679(.A(KEYINPUT60), .B(new_n1104), .C1(new_n1007), .C2(G1348), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1103), .A2(new_n1105), .A3(new_n605), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1107), .A2(KEYINPUT60), .A3(new_n604), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1089), .A2(new_n1093), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n1083), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n1097), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT61), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1109), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1101), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT58), .B(G1341), .ZN(new_n1116));
  OAI22_X1  g691(.A1(new_n999), .A2(G1996), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n553), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1118), .B(KEYINPUT59), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1098), .A2(new_n1114), .A3(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1096), .B1(new_n604), .B2(new_n1107), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n1097), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1078), .B(new_n1123), .C1(new_n1047), .C2(new_n1046), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1023), .B1(new_n1067), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT118), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1032), .A2(G286), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1126), .B1(new_n1022), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT63), .ZN(new_n1130));
  OR2_X1    g705(.A1(new_n1021), .A2(new_n994), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1009), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n964), .B1(new_n1013), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n988), .B1(new_n1133), .B2(new_n994), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1131), .A2(new_n1134), .A3(KEYINPUT118), .A4(new_n1127), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1129), .A2(new_n1130), .A3(new_n1135), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n1133), .A2(new_n994), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1137), .A2(new_n1134), .A3(KEYINPUT63), .A4(new_n1127), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n989), .A2(new_n994), .A3(new_n1133), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n984), .A2(new_n969), .A3(new_n748), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1141), .B1(new_n978), .B2(new_n979), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n968), .B(KEYINPUT115), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1139), .A2(new_n1140), .A3(new_n1144), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n957), .B(new_n963), .C1(new_n1125), .C2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n956), .ZN(new_n1147));
  OAI22_X1  g722(.A1(new_n953), .A2(new_n1147), .B1(G2067), .B2(new_n846), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1148), .A2(new_n950), .ZN(new_n1149));
  INV_X1    g724(.A(G1996), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n950), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT46), .ZN(new_n1152));
  OR3_X1    g727(.A1(new_n1151), .A2(KEYINPUT126), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n806), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n951), .A2(new_n1154), .ZN(new_n1155));
  AOI22_X1  g730(.A1(new_n1155), .A2(new_n950), .B1(KEYINPUT126), .B2(new_n1152), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1151), .B1(KEYINPUT126), .B2(new_n1152), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1153), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  XOR2_X1   g733(.A(new_n1158), .B(KEYINPUT47), .Z(new_n1159));
  XNOR2_X1  g734(.A(new_n960), .B(KEYINPUT48), .ZN(new_n1160));
  XOR2_X1   g735(.A(new_n957), .B(KEYINPUT127), .Z(new_n1161));
  AOI211_X1 g736(.A(new_n1149), .B(new_n1159), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1146), .A2(new_n1162), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g738(.A1(new_n651), .A2(new_n667), .ZN(new_n1165));
  AOI21_X1  g739(.A(new_n1165), .B1(new_n882), .B2(new_n877), .ZN(new_n1166));
  AND4_X1   g740(.A1(G319), .A2(new_n1166), .A3(new_n944), .A4(new_n689), .ZN(G308));
  NAND4_X1  g741(.A1(new_n1166), .A2(new_n944), .A3(G319), .A4(new_n689), .ZN(G225));
endmodule


