//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 0 0 1 1 1 1 1 1 0 0 0 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n557,
    new_n558, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1188, new_n1189, new_n1190;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT66), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT67), .B(G69), .Z(G235));
  XNOR2_X1  g013(.A(KEYINPUT68), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT69), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G235), .A2(G236), .A3(G237), .A4(G238), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT70), .Z(G319));
  INV_X1    g036(.A(G137), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT72), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT72), .A2(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(KEYINPUT3), .A3(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT73), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n468), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n465), .A2(KEYINPUT73), .A3(KEYINPUT3), .A4(new_n466), .ZN(new_n472));
  AOI211_X1 g047(.A(new_n462), .B(G2105), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  AND2_X1   g049(.A1(KEYINPUT72), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(KEYINPUT72), .A2(G2104), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G101), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  OAI21_X1  g055(.A(KEYINPUT74), .B1(new_n473), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g056(.A(G2105), .B1(new_n471), .B2(new_n472), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G137), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT74), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n483), .A2(new_n484), .A3(new_n479), .ZN(new_n485));
  XNOR2_X1  g060(.A(KEYINPUT3), .B(G2104), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G125), .ZN(new_n487));
  INV_X1    g062(.A(G113), .ZN(new_n488));
  OAI21_X1  g063(.A(KEYINPUT71), .B1(new_n488), .B2(new_n464), .ZN(new_n489));
  OR3_X1    g064(.A1(new_n488), .A2(new_n464), .A3(KEYINPUT71), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n487), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  AND3_X1   g067(.A1(new_n481), .A2(new_n485), .A3(new_n492), .ZN(G160));
  AOI21_X1  g068(.A(new_n474), .B1(new_n471), .B2(new_n472), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G124), .ZN(new_n495));
  OR2_X1    g070(.A1(G100), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G112), .C2(new_n474), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n498), .B1(G136), .B2(new_n482), .ZN(G162));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n486), .A2(new_n500), .A3(G138), .A4(new_n474), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n475), .A2(new_n476), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n469), .B1(new_n503), .B2(KEYINPUT3), .ZN(new_n504));
  INV_X1    g079(.A(new_n472), .ZN(new_n505));
  OAI211_X1 g080(.A(G138), .B(new_n474), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n502), .B1(new_n506), .B2(KEYINPUT4), .ZN(new_n507));
  OR2_X1    g082(.A1(G102), .A2(G2105), .ZN(new_n508));
  OAI211_X1 g083(.A(new_n508), .B(G2104), .C1(G114), .C2(new_n474), .ZN(new_n509));
  XNOR2_X1  g084(.A(new_n509), .B(KEYINPUT75), .ZN(new_n510));
  OAI211_X1 g085(.A(G126), .B(G2105), .C1(new_n504), .C2(new_n505), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n507), .A2(new_n512), .ZN(G164));
  XNOR2_X1  g088(.A(KEYINPUT5), .B(G543), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT6), .B(G651), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n518), .A2(G50), .A3(G543), .ZN(new_n519));
  XOR2_X1   g094(.A(new_n519), .B(KEYINPUT76), .Z(new_n520));
  AND2_X1   g095(.A1(new_n518), .A2(new_n514), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G88), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT77), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n520), .A2(KEYINPUT77), .A3(new_n522), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n517), .B1(new_n525), .B2(new_n526), .ZN(G166));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n518), .A2(G543), .ZN(new_n530));
  INV_X1    g105(.A(G51), .ZN(new_n531));
  INV_X1    g106(.A(G89), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n518), .A2(new_n514), .ZN(new_n533));
  OAI221_X1 g108(.A(new_n529), .B1(new_n530), .B2(new_n531), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT78), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n534), .A2(new_n536), .ZN(G168));
  XOR2_X1   g112(.A(KEYINPUT79), .B(G90), .Z(new_n538));
  INV_X1    g113(.A(G52), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n533), .A2(new_n538), .B1(new_n530), .B2(new_n539), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n516), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n540), .A2(new_n542), .ZN(G171));
  INV_X1    g118(.A(G81), .ZN(new_n544));
  INV_X1    g119(.A(G43), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n533), .A2(new_n544), .B1(new_n530), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(new_n514), .ZN(new_n548));
  INV_X1    g123(.A(G56), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT80), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n516), .B1(new_n550), .B2(new_n551), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n546), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  NAND3_X1  g134(.A1(new_n518), .A2(G53), .A3(G543), .ZN(new_n560));
  XOR2_X1   g135(.A(new_n560), .B(KEYINPUT9), .Z(new_n561));
  AOI22_X1  g136(.A1(new_n514), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G91), .ZN(new_n563));
  OAI22_X1  g138(.A1(new_n562), .A2(new_n516), .B1(new_n533), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(G299));
  INV_X1    g141(.A(G171), .ZN(G301));
  INV_X1    g142(.A(G168), .ZN(G286));
  INV_X1    g143(.A(G166), .ZN(G303));
  AND2_X1   g144(.A1(new_n521), .A2(G87), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n571));
  INV_X1    g146(.A(G49), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n530), .B2(new_n572), .ZN(new_n573));
  OR2_X1    g148(.A1(new_n570), .A2(new_n573), .ZN(G288));
  INV_X1    g149(.A(G61), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT81), .B1(new_n548), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT81), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n514), .A2(new_n577), .A3(G61), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n576), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G651), .ZN(new_n581));
  INV_X1    g156(.A(new_n530), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G48), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n521), .A2(G86), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT82), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n586), .B(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n585), .A2(new_n588), .ZN(G305));
  INV_X1    g164(.A(G85), .ZN(new_n590));
  INV_X1    g165(.A(G47), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n533), .A2(new_n590), .B1(new_n530), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n593), .A2(new_n516), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G290));
  INV_X1    g171(.A(KEYINPUT83), .ZN(new_n597));
  NAND3_X1  g172(.A1(G301), .A2(new_n597), .A3(G868), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n548), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(G651), .B1(new_n582), .B2(G54), .ZN(new_n603));
  INV_X1    g178(.A(G92), .ZN(new_n604));
  XNOR2_X1  g179(.A(KEYINPUT84), .B(KEYINPUT10), .ZN(new_n605));
  OR3_X1    g180(.A1(new_n533), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n533), .B2(new_n604), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n603), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n597), .B1(G301), .B2(G868), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n599), .B1(new_n610), .B2(new_n611), .ZN(G284));
  AOI21_X1  g187(.A(new_n599), .B1(new_n610), .B2(new_n611), .ZN(G321));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(G868), .B2(new_n565), .ZN(G297));
  OAI21_X1  g190(.A(new_n614), .B1(G868), .B2(new_n565), .ZN(G280));
  INV_X1    g191(.A(new_n608), .ZN(new_n617));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND2_X1  g194(.A1(new_n552), .A2(new_n553), .ZN(new_n620));
  INV_X1    g195(.A(new_n546), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(new_n609), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n608), .A2(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(new_n609), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g201(.A(new_n486), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n627), .A2(new_n477), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT12), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2100), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n482), .A2(G135), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n494), .A2(G123), .ZN(new_n633));
  OR2_X1    g208(.A1(G99), .A2(G2105), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n634), .B(G2104), .C1(G111), .C2(new_n474), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n632), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n636), .A2(G2096), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(G2096), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n631), .A2(new_n637), .A3(new_n638), .ZN(G156));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(KEYINPUT14), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G1341), .B(G1348), .Z(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n645), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2451), .B(G2454), .Z(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(G14), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n649), .A2(new_n652), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(G401));
  XNOR2_X1  g231(.A(G2084), .B(G2090), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT86), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  AND2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(KEYINPUT88), .B(KEYINPUT18), .Z(new_n662));
  NOR2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2072), .B(G2078), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT87), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g241(.A(KEYINPUT17), .B1(new_n659), .B2(new_n660), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n662), .B1(new_n661), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n666), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2096), .B(G2100), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(G227));
  XNOR2_X1  g246(.A(G1956), .B(G2474), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT89), .ZN(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT90), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n673), .A2(KEYINPUT90), .A3(new_n674), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT19), .Z(new_n680));
  NAND3_X1  g255(.A1(new_n677), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT91), .B(KEYINPUT20), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n673), .A2(new_n674), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n680), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n685), .A2(new_n675), .A3(new_n686), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n683), .B(new_n687), .C1(new_n686), .C2(new_n685), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1991), .B(G1996), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1981), .B(G1986), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(G229));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G23), .ZN(new_n696));
  INV_X1    g271(.A(G288), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(new_n695), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT33), .ZN(new_n699));
  INV_X1    g274(.A(G1976), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n695), .A2(G22), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G166), .B2(new_n695), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G1971), .ZN(new_n704));
  NOR2_X1   g279(.A1(G6), .A2(G16), .ZN(new_n705));
  INV_X1    g280(.A(G305), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(G16), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT32), .B(G1981), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NOR3_X1   g284(.A1(new_n701), .A2(new_n704), .A3(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT34), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT92), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n714), .A2(G29), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(G29), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n718), .A2(G25), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n494), .A2(G119), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n482), .A2(G131), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n474), .A2(G107), .ZN(new_n722));
  OAI21_X1  g297(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n720), .B(new_n721), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n719), .B1(new_n724), .B2(new_n717), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT35), .B(G1991), .Z(new_n726));
  AND2_X1   g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n695), .A2(G24), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(new_n595), .B2(new_n695), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G1986), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n725), .A2(new_n726), .ZN(new_n731));
  NOR3_X1   g306(.A1(new_n727), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n712), .A2(new_n713), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT36), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n695), .A2(G20), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT23), .Z(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G299), .B2(G16), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G1956), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n695), .A2(G19), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n554), .B2(new_n695), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(G1341), .Z(new_n741));
  NAND2_X1  g316(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n718), .A2(G26), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT94), .Z(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT28), .ZN(new_n745));
  OR2_X1    g320(.A1(G104), .A2(G2105), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n746), .B(G2104), .C1(G116), .C2(new_n474), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT93), .Z(new_n748));
  NAND2_X1  g323(.A1(new_n482), .A2(G140), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n494), .A2(G128), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n745), .B1(new_n751), .B2(G29), .ZN(new_n752));
  INV_X1    g327(.A(G2067), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(G2072), .ZN(new_n755));
  INV_X1    g330(.A(G33), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n756), .A2(G29), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n482), .A2(G139), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n486), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT95), .B(KEYINPUT25), .Z(new_n760));
  NAND3_X1  g335(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  OAI221_X1 g338(.A(new_n758), .B1(new_n474), .B2(new_n759), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT96), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n757), .B1(new_n766), .B2(G29), .ZN(new_n767));
  AOI211_X1 g342(.A(new_n742), .B(new_n754), .C1(new_n755), .C2(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n717), .A2(G27), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G164), .B2(new_n717), .ZN(new_n770));
  INV_X1    g345(.A(G2078), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT24), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n773), .A2(G34), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n773), .A2(G34), .ZN(new_n775));
  NOR3_X1   g350(.A1(new_n717), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G160), .B2(G29), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n772), .B1(new_n777), .B2(G2084), .ZN(new_n778));
  NAND2_X1  g353(.A1(G162), .A2(new_n717), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G35), .B2(new_n717), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT29), .B(G2090), .Z(new_n781));
  OR2_X1    g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  NOR2_X1   g358(.A1(G4), .A2(G16), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n617), .B2(G16), .ZN(new_n785));
  INV_X1    g360(.A(G1348), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n695), .A2(G5), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G171), .B2(new_n695), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n789), .A2(G1961), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n782), .A2(new_n783), .A3(new_n787), .A4(new_n790), .ZN(new_n791));
  AOI211_X1 g366(.A(new_n778), .B(new_n791), .C1(G2084), .C2(new_n777), .ZN(new_n792));
  INV_X1    g367(.A(G32), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n793), .A2(G29), .ZN(new_n794));
  NAND3_X1  g369(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT26), .Z(new_n796));
  INV_X1    g371(.A(G105), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n477), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n494), .B2(G129), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT98), .ZN(new_n800));
  AND3_X1   g375(.A1(new_n482), .A2(new_n800), .A3(G141), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n800), .B1(new_n482), .B2(G141), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n799), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n803), .A2(KEYINPUT99), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(KEYINPUT99), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n794), .B1(new_n806), .B2(G29), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT27), .B(G1996), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n768), .B(new_n792), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n767), .A2(new_n755), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT97), .Z(new_n811));
  NAND2_X1  g386(.A1(new_n807), .A2(new_n808), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n789), .A2(G1961), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT101), .Z(new_n814));
  NAND2_X1  g389(.A1(new_n695), .A2(G21), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G168), .B2(new_n695), .ZN(new_n816));
  INV_X1    g391(.A(G1966), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n636), .A2(new_n718), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT31), .B(G11), .Z(new_n820));
  XOR2_X1   g395(.A(KEYINPUT100), .B(G28), .Z(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(KEYINPUT30), .ZN(new_n822));
  AOI21_X1  g397(.A(G29), .B1(new_n821), .B2(KEYINPUT30), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n820), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n814), .A2(new_n818), .A3(new_n819), .A4(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT102), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n811), .A2(new_n812), .A3(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n809), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n734), .A2(new_n828), .ZN(G150));
  INV_X1    g404(.A(G150), .ZN(G311));
  NOR2_X1   g405(.A1(new_n608), .A2(new_n618), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n518), .A2(G55), .A3(G543), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  AND3_X1   g410(.A1(new_n514), .A2(new_n518), .A3(G93), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT104), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  AOI22_X1  g414(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n840), .A2(new_n516), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n554), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n837), .A2(new_n838), .ZN(new_n843));
  NOR3_X1   g418(.A1(new_n835), .A2(new_n836), .A3(KEYINPUT104), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n841), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n845), .A2(new_n622), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n833), .B(new_n847), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n848), .A2(KEYINPUT39), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n848), .A2(KEYINPUT39), .ZN(new_n850));
  NOR3_X1   g425(.A1(new_n849), .A2(new_n850), .A3(G860), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n845), .A2(G860), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT37), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n851), .A2(new_n853), .ZN(G145));
  NAND2_X1  g429(.A1(new_n494), .A2(G130), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n474), .A2(G118), .ZN(new_n856));
  OAI21_X1  g431(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n858), .B1(G142), .B2(new_n482), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(new_n629), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n724), .ZN(new_n861));
  INV_X1    g436(.A(new_n512), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT105), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n863), .B1(new_n864), .B2(new_n501), .ZN(new_n865));
  AOI211_X1 g440(.A(KEYINPUT105), .B(new_n502), .C1(new_n506), .C2(KEYINPUT4), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n862), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n804), .A2(new_n805), .A3(new_n751), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n751), .B1(new_n804), .B2(new_n805), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n867), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n870), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n500), .B1(new_n482), .B2(G138), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT105), .B1(new_n873), .B2(new_n502), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n864), .A2(new_n863), .A3(new_n501), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n512), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n872), .A2(new_n876), .A3(new_n868), .ZN(new_n877));
  AND3_X1   g452(.A1(new_n871), .A2(new_n877), .A3(new_n764), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n766), .B1(new_n871), .B2(new_n877), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n861), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n871), .A2(new_n877), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(new_n765), .ZN(new_n882));
  INV_X1    g457(.A(new_n861), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n871), .A2(new_n877), .A3(new_n764), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n880), .A2(new_n885), .ZN(new_n886));
  XOR2_X1   g461(.A(G160), .B(new_n636), .Z(new_n887));
  XOR2_X1   g462(.A(new_n887), .B(G162), .Z(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(G37), .ZN(new_n890));
  INV_X1    g465(.A(new_n888), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n880), .A2(new_n885), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n889), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT106), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(G37), .B1(new_n886), .B2(new_n888), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n896), .A2(KEYINPUT106), .A3(new_n892), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n895), .A2(new_n897), .A3(KEYINPUT40), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT40), .B1(new_n895), .B2(new_n897), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(G395));
  NAND2_X1  g475(.A1(new_n845), .A2(new_n609), .ZN(new_n901));
  XOR2_X1   g476(.A(G288), .B(KEYINPUT108), .Z(new_n902));
  OR2_X1    g477(.A1(new_n902), .A2(new_n706), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n706), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(G303), .A2(new_n595), .ZN(new_n906));
  NAND2_X1  g481(.A1(G166), .A2(G290), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n903), .A2(new_n906), .A3(new_n907), .A4(new_n904), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n911), .A2(KEYINPUT109), .ZN(new_n912));
  XOR2_X1   g487(.A(KEYINPUT110), .B(KEYINPUT42), .Z(new_n913));
  XNOR2_X1  g488(.A(new_n912), .B(new_n913), .ZN(new_n914));
  XOR2_X1   g489(.A(new_n847), .B(new_n624), .Z(new_n915));
  NAND2_X1  g490(.A1(G299), .A2(new_n617), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n565), .A2(new_n608), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT107), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT107), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n919), .B1(G299), .B2(new_n617), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n915), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n916), .A2(new_n917), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n923), .A2(KEYINPUT41), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n918), .A2(new_n920), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n924), .B1(new_n925), .B2(KEYINPUT41), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n922), .B1(new_n915), .B2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n914), .B(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n901), .B1(new_n928), .B2(new_n609), .ZN(G295));
  OAI21_X1  g504(.A(new_n901), .B1(new_n928), .B2(new_n609), .ZN(G331));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n839), .A2(new_n554), .A3(new_n841), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n845), .A2(new_n622), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n932), .A2(new_n933), .A3(G301), .ZN(new_n934));
  AOI21_X1  g509(.A(G301), .B1(new_n932), .B2(new_n933), .ZN(new_n935));
  NOR3_X1   g510(.A1(new_n934), .A2(new_n935), .A3(G286), .ZN(new_n936));
  OAI21_X1  g511(.A(G171), .B1(new_n842), .B2(new_n846), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n932), .A2(new_n933), .A3(G301), .ZN(new_n938));
  AOI21_X1  g513(.A(G168), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT111), .B1(new_n940), .B2(new_n921), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n925), .A2(KEYINPUT41), .ZN(new_n942));
  INV_X1    g517(.A(new_n924), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n937), .A2(G168), .A3(new_n938), .ZN(new_n944));
  OAI21_X1  g519(.A(G286), .B1(new_n934), .B2(new_n935), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n942), .A2(new_n943), .A3(new_n944), .A4(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n921), .B1(new_n945), .B2(new_n944), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT111), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n941), .A2(new_n911), .A3(new_n946), .A4(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT113), .ZN(new_n951));
  AOI22_X1  g526(.A1(new_n926), .A2(new_n940), .B1(new_n947), .B2(new_n948), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT113), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n952), .A2(new_n953), .A3(new_n911), .A4(new_n941), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n940), .A2(KEYINPUT41), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n956), .A2(new_n925), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n911), .B1(new_n956), .B2(new_n923), .ZN(new_n958));
  AOI21_X1  g533(.A(G37), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n955), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(KEYINPUT43), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT43), .B1(new_n951), .B2(new_n954), .ZN(new_n962));
  INV_X1    g537(.A(new_n911), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n946), .A2(new_n949), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n947), .A2(new_n948), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT112), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n966), .A2(new_n967), .A3(new_n890), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n967), .B1(new_n966), .B2(new_n890), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n962), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n931), .B1(new_n961), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n955), .B1(new_n968), .B2(new_n969), .ZN(new_n972));
  AOI22_X1  g547(.A1(new_n972), .A2(KEYINPUT43), .B1(new_n959), .B2(new_n962), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n971), .B1(new_n931), .B2(new_n973), .ZN(G397));
  INV_X1    g549(.A(G1384), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT45), .B1(new_n867), .B2(new_n975), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n492), .A2(G40), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n481), .A2(new_n485), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n980), .A2(G1996), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n981), .A2(new_n805), .A3(new_n804), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT114), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n980), .B(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n751), .B(new_n753), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n987), .B1(new_n806), .B2(G1996), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n982), .B1(new_n985), .B2(new_n988), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n989), .B(KEYINPUT115), .ZN(new_n990));
  INV_X1    g565(.A(new_n726), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n724), .A2(new_n991), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n724), .A2(new_n991), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n984), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n990), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n980), .ZN(new_n996));
  XOR2_X1   g571(.A(new_n595), .B(G1986), .Z(new_n997));
  AOI21_X1  g572(.A(new_n995), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT116), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n1000), .A2(G1384), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n999), .B1(new_n876), .B2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n867), .A2(KEYINPUT116), .A3(new_n1001), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n975), .B1(new_n507), .B2(new_n512), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n1000), .ZN(new_n1007));
  XNOR2_X1  g582(.A(KEYINPUT56), .B(G2072), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1005), .A2(new_n1007), .A3(new_n979), .A4(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G1956), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n874), .A2(new_n875), .ZN(new_n1011));
  AOI21_X1  g586(.A(G1384), .B1(new_n1011), .B2(new_n862), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT50), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n979), .B1(KEYINPUT50), .B2(new_n1006), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1010), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1009), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n565), .B(KEYINPUT57), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n867), .A2(new_n979), .A3(new_n975), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT120), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1012), .A2(KEYINPUT120), .A3(new_n979), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n867), .A2(new_n1013), .A3(new_n975), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT117), .B1(new_n1006), .B2(KEYINPUT50), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n1006), .A2(KEYINPUT117), .A3(KEYINPUT50), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1026), .B(new_n979), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n1025), .A2(new_n753), .B1(new_n1029), .B2(new_n786), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n1030), .A2(new_n608), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1009), .A2(new_n1018), .A3(new_n1016), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1020), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1018), .B1(new_n1009), .B2(new_n1016), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT122), .ZN(new_n1035));
  NOR3_X1   g610(.A1(new_n1032), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1017), .A2(new_n1035), .A3(new_n1019), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT61), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1009), .A2(new_n1018), .A3(new_n1016), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1020), .A2(KEYINPUT61), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1029), .A2(new_n786), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT120), .B1(new_n1012), .B2(new_n979), .ZN(new_n1044));
  NOR4_X1   g619(.A1(new_n876), .A2(new_n978), .A3(new_n1022), .A4(G1384), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n753), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT60), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT123), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1047), .B1(new_n617), .B2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1043), .A2(new_n1046), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n608), .A2(KEYINPUT123), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1050), .B(new_n1051), .C1(new_n1030), .C2(KEYINPUT60), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1030), .A2(KEYINPUT123), .A3(KEYINPUT60), .A4(new_n608), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1042), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1040), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n978), .A2(G1996), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1005), .A2(new_n1007), .A3(new_n1056), .ZN(new_n1057));
  XOR2_X1   g632(.A(KEYINPUT58), .B(G1341), .Z(new_n1058));
  NAND3_X1  g633(.A1(new_n1023), .A2(new_n1024), .A3(new_n1058), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1057), .A2(new_n1059), .A3(KEYINPUT121), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT121), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n554), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g637(.A(new_n1062), .B(KEYINPUT59), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1033), .B1(new_n1055), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n979), .B1(G164), .B2(new_n1002), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n817), .B1(new_n976), .B2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n978), .A2(G2084), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1026), .B(new_n1067), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(G286), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1066), .A2(new_n1068), .A3(G168), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1070), .A2(KEYINPUT51), .A3(G8), .A4(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT124), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1071), .A2(G8), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1072), .A2(new_n1073), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1073), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1005), .A2(new_n771), .A3(new_n1007), .A4(new_n979), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT53), .ZN(new_n1081));
  INV_X1    g656(.A(G1961), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n1080), .A2(new_n1081), .B1(new_n1082), .B2(new_n1029), .ZN(new_n1083));
  INV_X1    g658(.A(new_n481), .ZN(new_n1084));
  INV_X1    g659(.A(new_n485), .ZN(new_n1085));
  OR3_X1    g660(.A1(new_n1084), .A2(new_n1085), .A3(KEYINPUT125), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT125), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1086), .A2(new_n977), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT126), .ZN(new_n1089));
  NOR3_X1   g664(.A1(new_n976), .A2(new_n1081), .A3(G2078), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT126), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1086), .A2(new_n1091), .A3(new_n977), .A4(new_n1087), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1089), .A2(new_n1090), .A3(new_n1005), .A4(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1083), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(G171), .ZN(new_n1095));
  OR4_X1    g670(.A1(new_n1081), .A2(new_n976), .A3(new_n1065), .A4(G2078), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1083), .A2(G301), .A3(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1095), .A2(KEYINPUT54), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT54), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1094), .A2(G171), .ZN(new_n1100));
  AOI21_X1  g675(.A(G301), .B1(new_n1083), .B2(new_n1096), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1099), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(G8), .ZN(new_n1103));
  NOR2_X1   g678(.A1(G166), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT55), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1105), .A2(KEYINPUT118), .ZN(new_n1106));
  OR2_X1    g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1104), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1107), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1005), .A2(new_n1007), .A3(new_n979), .ZN(new_n1111));
  INV_X1    g686(.A(G1971), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1029), .A2(G2090), .ZN(new_n1114));
  OAI211_X1 g689(.A(G8), .B(new_n1110), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1110), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1012), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1015), .B1(new_n1117), .B2(KEYINPUT50), .ZN(new_n1118));
  INV_X1    g693(.A(G2090), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1111), .A2(new_n1112), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1116), .B1(new_n1120), .B2(new_n1103), .ZN(new_n1121));
  INV_X1    g696(.A(new_n586), .ZN(new_n1122));
  OAI21_X1  g697(.A(G1981), .B1(new_n584), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(G1981), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n588), .A2(new_n581), .A3(new_n1124), .A4(new_n583), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1123), .A2(new_n1125), .A3(KEYINPUT119), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT119), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1127), .B(G1981), .C1(new_n584), .C2(new_n1122), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT49), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1103), .B1(new_n1012), .B2(new_n979), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT49), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1126), .A2(new_n1132), .A3(new_n1128), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1130), .A2(new_n1131), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n697), .A2(G1976), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1131), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT52), .B1(G288), .B2(new_n700), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1134), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  AND2_X1   g714(.A1(new_n1136), .A2(KEYINPUT52), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AND3_X1   g716(.A1(new_n1115), .A2(new_n1121), .A3(new_n1141), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1079), .A2(new_n1098), .A3(new_n1102), .A4(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1064), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT62), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1145), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1072), .A2(new_n1076), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(KEYINPUT124), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1072), .A2(new_n1076), .A3(new_n1073), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1148), .A2(KEYINPUT62), .A3(new_n1149), .ZN(new_n1150));
  AND4_X1   g725(.A1(new_n1101), .A2(new_n1115), .A3(new_n1121), .A4(new_n1141), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1146), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n1134), .A2(new_n700), .A3(new_n697), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1125), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1131), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1141), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1155), .B1(new_n1156), .B2(new_n1115), .ZN(new_n1157));
  AOI211_X1 g732(.A(new_n1103), .B(G286), .C1(new_n1066), .C2(new_n1068), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1115), .A2(new_n1121), .A3(new_n1141), .A4(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT63), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(G8), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(new_n1116), .ZN(new_n1163));
  AND2_X1   g738(.A1(new_n1158), .A2(KEYINPUT63), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1163), .A2(new_n1115), .A3(new_n1164), .A4(new_n1141), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1157), .B1(new_n1161), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1152), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n998), .B1(new_n1144), .B2(new_n1167), .ZN(new_n1168));
  XOR2_X1   g743(.A(new_n981), .B(KEYINPUT46), .Z(new_n1169));
  OAI21_X1  g744(.A(new_n984), .B1(new_n806), .B2(new_n987), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(KEYINPUT47), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n980), .A2(G1986), .A3(G290), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1173), .B(KEYINPUT48), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1172), .B1(new_n995), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n990), .A2(new_n992), .ZN(new_n1176));
  OR2_X1    g751(.A1(new_n751), .A2(G2067), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n985), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1175), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1168), .A2(new_n1179), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g755(.A(G319), .B1(new_n654), .B2(new_n655), .ZN(new_n1182));
  NOR3_X1   g756(.A1(G229), .A2(G227), .A3(new_n1182), .ZN(new_n1183));
  INV_X1    g757(.A(new_n897), .ZN(new_n1184));
  AOI21_X1  g758(.A(KEYINPUT106), .B1(new_n896), .B2(new_n892), .ZN(new_n1185));
  OAI21_X1  g759(.A(new_n1183), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g760(.A1(new_n1186), .A2(new_n973), .ZN(G308));
  NAND2_X1  g761(.A1(new_n895), .A2(new_n897), .ZN(new_n1188));
  AND2_X1   g762(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n1189));
  AND2_X1   g763(.A1(new_n962), .A2(new_n959), .ZN(new_n1190));
  OAI211_X1 g764(.A(new_n1188), .B(new_n1183), .C1(new_n1189), .C2(new_n1190), .ZN(G225));
endmodule


