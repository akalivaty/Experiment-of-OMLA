//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 1 1 0 0 0 1 1 1 0 0 1 1 1 1 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 0 1 0 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314;
  NOR2_X1   g0000(.A1(G50), .A2(G58), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  INV_X1    g0003(.A(G77), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n202), .A2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NOR2_X1   g0007(.A1(G58), .A2(G68), .ZN(new_n208));
  OR2_X1    g0008(.A1(new_n208), .A2(KEYINPUT64), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(KEYINPUT64), .ZN(new_n210));
  NAND3_X1  g0010(.A1(new_n209), .A2(G50), .A3(new_n210), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT65), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT0), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G50), .ZN(new_n222));
  INV_X1    g0022(.A(G226), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(KEYINPUT66), .B(G244), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n224), .B1(G77), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(KEYINPUT67), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n229));
  NAND3_X1  g0029(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n226), .A2(KEYINPUT67), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n217), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT68), .Z(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n216), .B(new_n220), .C1(new_n234), .C2(KEYINPUT1), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n235), .B1(KEYINPUT1), .B2(new_n234), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  NAND2_X1  g0044(.A1(G68), .A2(G77), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n205), .A2(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n246), .B(KEYINPUT69), .Z(new_n247));
  XOR2_X1   g0047(.A(G50), .B(G58), .Z(new_n248));
  XOR2_X1   g0048(.A(new_n247), .B(new_n248), .Z(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT70), .ZN(new_n251));
  XOR2_X1   g0051(.A(G107), .B(G116), .Z(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n249), .B(new_n253), .ZN(G351));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n213), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G20), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  OAI22_X1  g0059(.A1(new_n259), .A2(new_n204), .B1(new_n214), .B2(G68), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n214), .A2(new_n257), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(new_n222), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n256), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g0063(.A(new_n263), .B(KEYINPUT11), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(G13), .A3(G20), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(KEYINPUT73), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT73), .ZN(new_n268));
  NAND4_X1  g0068(.A1(new_n268), .A2(new_n265), .A3(G13), .A4(G20), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n256), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n265), .A2(G20), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(G68), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n264), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n267), .A2(new_n269), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G68), .ZN(new_n275));
  XNOR2_X1  g0075(.A(new_n275), .B(KEYINPUT12), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT14), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT71), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G41), .A2(G45), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n280), .B1(new_n281), .B2(G1), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G33), .A2(G41), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(G1), .A3(G13), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n265), .B(KEYINPUT71), .C1(G41), .C2(G45), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n282), .A2(G238), .A3(new_n284), .A4(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n281), .A2(G1), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n287), .A2(new_n284), .A3(G274), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT77), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n286), .A2(KEYINPUT77), .A3(new_n288), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G232), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G1698), .ZN(new_n295));
  AND2_X1   g0095(.A1(KEYINPUT3), .A2(G33), .ZN(new_n296));
  NOR2_X1   g0096(.A1(KEYINPUT3), .A2(G33), .ZN(new_n297));
  OAI221_X1 g0097(.A(new_n295), .B1(G226), .B2(G1698), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(G33), .A2(G97), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT75), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT75), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n301), .A2(G33), .A3(G97), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT76), .ZN(new_n305));
  INV_X1    g0105(.A(new_n284), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT76), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n298), .A2(new_n307), .A3(new_n303), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n305), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT13), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n293), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n310), .B1(new_n293), .B2(new_n309), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n279), .B(G169), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n293), .A2(new_n309), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT13), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n316), .A2(G179), .A3(new_n311), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n311), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n279), .B1(new_n319), .B2(G169), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n278), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n316), .A2(G190), .A3(new_n311), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n277), .ZN(new_n323));
  INV_X1    g0123(.A(G200), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n324), .B1(new_n316), .B2(new_n311), .ZN(new_n325));
  OR2_X1    g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT78), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n321), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n327), .B1(new_n321), .B2(new_n326), .ZN(new_n330));
  INV_X1    g0130(.A(G1698), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT3), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n257), .ZN(new_n333));
  NAND2_X1  g0133(.A1(KEYINPUT3), .A2(G33), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n331), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G223), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n333), .A2(new_n334), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n337), .A2(G222), .A3(new_n331), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n296), .A2(new_n297), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(G77), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n336), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n306), .ZN(new_n342));
  INV_X1    g0142(.A(new_n288), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n282), .A2(new_n284), .A3(new_n285), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n343), .B1(new_n345), .B2(G226), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G179), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n274), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n222), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT74), .ZN(new_n353));
  INV_X1    g0153(.A(new_n271), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n353), .B1(new_n354), .B2(new_n222), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n271), .A2(KEYINPUT74), .A3(G50), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n270), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n352), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g0158(.A(KEYINPUT8), .B(G58), .ZN(new_n359));
  INV_X1    g0159(.A(G150), .ZN(new_n360));
  OAI22_X1  g0160(.A1(new_n359), .A2(new_n259), .B1(new_n360), .B2(new_n261), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n214), .B1(new_n201), .B2(new_n203), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n256), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT72), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI211_X1 g0165(.A(KEYINPUT72), .B(new_n256), .C1(new_n361), .C2(new_n362), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n358), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G169), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n347), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n350), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n366), .A2(new_n352), .A3(new_n357), .ZN(new_n372));
  INV_X1    g0172(.A(new_n362), .ZN(new_n373));
  OAI221_X1 g0173(.A(new_n373), .B1(new_n360), .B2(new_n261), .C1(new_n259), .C2(new_n359), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT72), .B1(new_n374), .B2(new_n256), .ZN(new_n375));
  OAI21_X1  g0175(.A(KEYINPUT9), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT9), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n358), .A2(new_n365), .A3(new_n377), .A4(new_n366), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n324), .B1(new_n342), .B2(new_n346), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n380), .B1(new_n348), .B2(G190), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT10), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT10), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n379), .A2(new_n381), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n371), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT16), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT7), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n337), .B2(G20), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n339), .A2(KEYINPUT7), .A3(new_n214), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n203), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(KEYINPUT79), .A2(G58), .A3(G68), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT79), .B1(G58), .B2(G68), .ZN(new_n394));
  NOR3_X1   g0194(.A1(new_n393), .A2(new_n394), .A3(new_n208), .ZN(new_n395));
  INV_X1    g0195(.A(G159), .ZN(new_n396));
  OAI22_X1  g0196(.A1(new_n395), .A2(new_n214), .B1(new_n396), .B2(new_n261), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n387), .B1(new_n391), .B2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT7), .B1(new_n339), .B2(new_n214), .ZN(new_n399));
  NOR4_X1   g0199(.A1(new_n296), .A2(new_n297), .A3(new_n388), .A4(G20), .ZN(new_n400));
  OAI21_X1  g0200(.A(G68), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n261), .A2(new_n396), .ZN(new_n402));
  INV_X1    g0202(.A(new_n394), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n403), .B(new_n392), .C1(G58), .C2(G68), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n402), .B1(new_n404), .B2(G20), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n401), .A2(new_n405), .A3(KEYINPUT16), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n398), .A2(new_n406), .A3(new_n256), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n359), .B1(new_n265), .B2(G20), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n351), .A2(new_n359), .B1(new_n408), .B2(new_n270), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  OAI211_X1 g0211(.A(G223), .B(new_n331), .C1(new_n296), .C2(new_n297), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT80), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n337), .A2(KEYINPUT80), .A3(G223), .A4(new_n331), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n335), .A2(G226), .B1(G33), .B2(G87), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n284), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n288), .B1(new_n344), .B2(new_n294), .ZN(new_n419));
  OAI21_X1  g0219(.A(G200), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n419), .ZN(new_n421));
  OAI211_X1 g0221(.A(G226), .B(G1698), .C1(new_n296), .C2(new_n297), .ZN(new_n422));
  INV_X1    g0222(.A(G87), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n422), .B1(new_n257), .B2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n424), .B1(new_n414), .B2(new_n415), .ZN(new_n425));
  OAI211_X1 g0225(.A(G190), .B(new_n421), .C1(new_n425), .C2(new_n284), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n420), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT81), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n411), .A2(new_n427), .A3(new_n428), .A4(KEYINPUT17), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT17), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n407), .A2(new_n420), .A3(new_n409), .A4(new_n426), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n430), .B1(new_n431), .B2(KEYINPUT81), .ZN(new_n432));
  AND2_X1   g0232(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(G169), .B1(new_n418), .B2(new_n419), .ZN(new_n434));
  OAI211_X1 g0234(.A(G179), .B(new_n421), .C1(new_n425), .C2(new_n284), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n410), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT18), .ZN(new_n438));
  XNOR2_X1  g0238(.A(new_n437), .B(new_n438), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n335), .A2(G238), .B1(new_n339), .B2(G107), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n337), .A2(G232), .A3(new_n331), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n306), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n343), .B1(new_n345), .B2(new_n225), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n368), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n270), .A2(G77), .A3(new_n271), .ZN(new_n447));
  NAND2_X1  g0247(.A1(G20), .A2(G77), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n448), .B1(new_n359), .B2(new_n261), .ZN(new_n449));
  XNOR2_X1  g0249(.A(KEYINPUT15), .B(G87), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n449), .B1(new_n258), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n256), .ZN(new_n453));
  OAI221_X1 g0253(.A(new_n447), .B1(G77), .B2(new_n274), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n446), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n445), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n349), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n454), .B1(G200), .B2(new_n445), .ZN(new_n459));
  INV_X1    g0259(.A(G190), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n459), .B1(new_n460), .B2(new_n445), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n386), .A2(new_n433), .A3(new_n439), .A4(new_n462), .ZN(new_n463));
  NOR3_X1   g0263(.A1(new_n329), .A2(new_n330), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G45), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(G1), .ZN(new_n466));
  AND2_X1   g0266(.A1(KEYINPUT5), .A2(G41), .ZN(new_n467));
  NOR2_X1   g0267(.A1(KEYINPUT5), .A2(G41), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AND2_X1   g0269(.A1(new_n469), .A2(new_n284), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G257), .ZN(new_n471));
  XNOR2_X1  g0271(.A(KEYINPUT5), .B(G41), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n472), .A2(G274), .A3(new_n284), .A4(new_n466), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(G244), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n475), .B1(new_n333), .B2(new_n334), .ZN(new_n476));
  AND2_X1   g0276(.A1(new_n331), .A2(KEYINPUT4), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n476), .A2(new_n477), .B1(G33), .B2(G283), .ZN(new_n478));
  OAI211_X1 g0278(.A(G244), .B(new_n331), .C1(new_n296), .C2(new_n297), .ZN(new_n479));
  XOR2_X1   g0279(.A(KEYINPUT82), .B(KEYINPUT4), .Z(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT83), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n482), .B1(new_n335), .B2(G250), .ZN(new_n483));
  OAI211_X1 g0283(.A(G250), .B(G1698), .C1(new_n296), .C2(new_n297), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(KEYINPUT83), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n478), .B(new_n481), .C1(new_n483), .C2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT84), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n284), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n484), .A2(KEYINPUT83), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n337), .A2(new_n482), .A3(G250), .A4(G1698), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n491), .A2(KEYINPUT84), .A3(new_n481), .A4(new_n478), .ZN(new_n492));
  AOI211_X1 g0292(.A(G179), .B(new_n474), .C1(new_n488), .C2(new_n492), .ZN(new_n493));
  AND2_X1   g0293(.A1(new_n489), .A2(new_n490), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G33), .A2(G283), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n337), .A2(G244), .A3(new_n477), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n481), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n487), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n498), .A2(new_n492), .A3(new_n306), .ZN(new_n499));
  INV_X1    g0299(.A(new_n474), .ZN(new_n500));
  AOI21_X1  g0300(.A(G169), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT6), .ZN(new_n502));
  INV_X1    g0302(.A(G97), .ZN(new_n503));
  NOR3_X1   g0303(.A1(new_n502), .A2(new_n503), .A3(G107), .ZN(new_n504));
  XNOR2_X1  g0304(.A(G97), .B(G107), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n504), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  OAI22_X1  g0306(.A1(new_n506), .A2(new_n214), .B1(new_n204), .B2(new_n261), .ZN(new_n507));
  INV_X1    g0307(.A(G107), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n508), .B1(new_n389), .B2(new_n390), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n256), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n351), .A2(new_n503), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n257), .A2(G1), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n270), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G97), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n510), .A2(new_n511), .A3(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NOR3_X1   g0318(.A1(new_n493), .A2(new_n501), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n474), .B1(new_n488), .B2(new_n492), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G190), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT85), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n324), .B1(new_n499), .B2(new_n500), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n499), .A2(KEYINPUT85), .A3(G190), .A4(new_n500), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n525), .A2(new_n518), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n519), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT21), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n274), .A2(new_n453), .A3(G116), .A4(new_n513), .ZN(new_n529));
  INV_X1    g0329(.A(G116), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n255), .A2(new_n213), .B1(G20), .B2(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n495), .B(new_n214), .C1(G33), .C2(new_n503), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT20), .ZN(new_n534));
  OR2_X1    g0334(.A1(new_n534), .A2(KEYINPUT88), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(KEYINPUT88), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n533), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n267), .A2(new_n530), .A3(new_n269), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n531), .A2(KEYINPUT88), .A3(new_n532), .A4(new_n534), .ZN(new_n539));
  AND4_X1   g0339(.A1(new_n529), .A2(new_n537), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n331), .A2(G264), .ZN(new_n541));
  NOR2_X1   g0341(.A1(G257), .A2(G1698), .ZN(new_n542));
  OAI22_X1  g0342(.A1(new_n541), .A2(new_n542), .B1(new_n296), .B2(new_n297), .ZN(new_n543));
  OR2_X1    g0343(.A1(KEYINPUT87), .A2(G303), .ZN(new_n544));
  NAND2_X1  g0344(.A1(KEYINPUT87), .A2(G303), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n544), .A2(new_n333), .A3(new_n334), .A4(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n543), .A2(new_n546), .A3(new_n306), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n469), .A2(G270), .A3(new_n284), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n547), .A2(new_n473), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G169), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n528), .B1(new_n540), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(G200), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n547), .A2(G190), .A3(new_n473), .A4(new_n548), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n540), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n547), .A2(G179), .A3(new_n473), .A4(new_n548), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n529), .A2(new_n537), .A3(new_n538), .A4(new_n539), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n557), .A2(KEYINPUT21), .A3(G169), .A4(new_n549), .ZN(new_n559));
  AND4_X1   g0359(.A1(new_n551), .A2(new_n554), .A3(new_n558), .A4(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(G244), .B(G1698), .C1(new_n296), .C2(new_n297), .ZN(new_n561));
  OAI211_X1 g0361(.A(G238), .B(new_n331), .C1(new_n296), .C2(new_n297), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G33), .A2(G116), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n306), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n284), .A2(G274), .A3(new_n466), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n265), .A2(G45), .ZN(new_n567));
  AND2_X1   g0367(.A1(G33), .A2(G41), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n567), .B(G250), .C1(new_n568), .C2(new_n213), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  AND4_X1   g0371(.A1(KEYINPUT86), .A2(new_n565), .A3(new_n571), .A4(new_n349), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n570), .B1(new_n564), .B2(new_n306), .ZN(new_n573));
  AOI21_X1  g0373(.A(KEYINPUT86), .B1(new_n573), .B2(new_n349), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(G169), .B1(new_n565), .B2(new_n571), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n274), .A2(new_n451), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n423), .A2(new_n503), .A3(new_n508), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT19), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n579), .B1(new_n300), .B2(new_n302), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n578), .B1(new_n580), .B2(G20), .ZN(new_n581));
  AOI21_X1  g0381(.A(G20), .B1(new_n333), .B2(new_n334), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n214), .A2(G33), .A3(G97), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n582), .A2(G68), .B1(new_n579), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n577), .B1(new_n585), .B2(new_n256), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n515), .A2(new_n451), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n576), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI211_X1 g0388(.A(new_n460), .B(new_n570), .C1(new_n306), .C2(new_n564), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n324), .B1(new_n565), .B2(new_n571), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n514), .A2(new_n423), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n453), .B1(new_n581), .B2(new_n584), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n592), .A2(new_n593), .A3(new_n577), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n575), .A2(new_n588), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT24), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n214), .B(G87), .C1(new_n296), .C2(new_n297), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(KEYINPUT22), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT22), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n337), .A2(new_n599), .A3(new_n214), .A4(G87), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT23), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(new_n214), .B2(G107), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n508), .A2(KEYINPUT23), .A3(G20), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n603), .A2(new_n604), .B1(new_n258), .B2(G116), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n596), .B1(new_n601), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n601), .A2(new_n596), .A3(new_n605), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n453), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n351), .A2(KEYINPUT25), .A3(new_n508), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT25), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(new_n274), .B2(G107), .ZN(new_n612));
  AOI22_X1  g0412(.A1(G107), .A2(new_n515), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n469), .A2(G264), .A3(new_n284), .ZN(new_n615));
  INV_X1    g0415(.A(G294), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n257), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(G250), .A2(G1698), .ZN(new_n618));
  INV_X1    g0418(.A(G257), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n618), .B1(new_n619), .B2(G1698), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n617), .B1(new_n620), .B2(new_n337), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n473), .B(new_n615), .C1(new_n621), .C2(new_n284), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n622), .A2(KEYINPUT89), .A3(G169), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n619), .A2(G1698), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n624), .B1(G250), .B2(G1698), .ZN(new_n625));
  OAI22_X1  g0425(.A1(new_n625), .A2(new_n339), .B1(new_n257), .B2(new_n616), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n306), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n627), .A2(G179), .A3(new_n473), .A4(new_n615), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT89), .B1(new_n622), .B2(G169), .ZN(new_n630));
  OAI22_X1  g0430(.A1(new_n609), .A2(new_n614), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n601), .A2(new_n596), .A3(new_n605), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n256), .B1(new_n632), .B2(new_n606), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n622), .A2(new_n324), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(G190), .B2(new_n622), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n633), .A2(new_n635), .A3(new_n613), .ZN(new_n636));
  AND4_X1   g0436(.A1(new_n560), .A2(new_n595), .A3(new_n631), .A4(new_n636), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n464), .A2(new_n527), .A3(new_n637), .ZN(G372));
  NAND2_X1  g0438(.A1(new_n383), .A2(new_n385), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n429), .A2(new_n432), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n323), .A2(new_n325), .ZN(new_n641));
  AOI211_X1 g0441(.A(new_n640), .B(new_n641), .C1(new_n321), .C2(new_n458), .ZN(new_n642));
  XNOR2_X1  g0442(.A(new_n437), .B(KEYINPUT18), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n639), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n370), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n464), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n573), .A2(new_n349), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n588), .A2(new_n648), .B1(new_n591), .B2(new_n594), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n623), .A2(new_n628), .ZN(new_n650));
  INV_X1    g0450(.A(new_n630), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n650), .A2(new_n651), .B1(new_n633), .B2(new_n613), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n551), .A2(new_n558), .A3(new_n559), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n649), .B(new_n636), .C1(new_n652), .C2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n524), .A2(new_n526), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n499), .A2(new_n349), .A3(new_n500), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n657), .B(new_n517), .C1(G169), .C2(new_n520), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n655), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n501), .A2(new_n518), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT26), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n660), .A2(new_n661), .A3(new_n657), .A4(new_n649), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n588), .A2(new_n648), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n575), .A2(new_n588), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n591), .A2(new_n594), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(KEYINPUT26), .B1(new_n658), .B2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n659), .A2(new_n664), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n646), .B1(new_n647), .B2(new_n670), .ZN(G369));
  NAND3_X1  g0471(.A1(new_n265), .A2(new_n214), .A3(G13), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G213), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g0475(.A(KEYINPUT90), .B(G343), .Z(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n557), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n560), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n653), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n679), .B1(new_n680), .B2(new_n678), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(G330), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n631), .A2(new_n636), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n677), .B1(new_n609), .B2(new_n614), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n677), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n686), .B1(new_n631), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n680), .A2(new_n677), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n684), .A2(new_n690), .ZN(new_n691));
  OAI211_X1 g0491(.A(new_n689), .B(new_n691), .C1(new_n631), .C2(new_n677), .ZN(G399));
  NAND2_X1  g0492(.A1(new_n525), .A2(new_n518), .ZN(new_n693));
  OAI21_X1  g0493(.A(KEYINPUT85), .B1(new_n520), .B2(new_n324), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n693), .B1(new_n521), .B2(new_n694), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n695), .A2(new_n654), .A3(new_n519), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n668), .A2(new_n663), .A3(new_n662), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n687), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT93), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT29), .ZN(new_n701));
  OAI211_X1 g0501(.A(KEYINPUT93), .B(new_n687), .C1(new_n696), .C2(new_n697), .ZN(new_n702));
  AND3_X1   g0502(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n663), .A2(new_n666), .ZN(new_n705));
  OAI21_X1  g0505(.A(KEYINPUT26), .B1(new_n658), .B2(new_n705), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n660), .A2(new_n661), .A3(new_n657), .A4(new_n595), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(new_n663), .A3(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT94), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n708), .A2(new_n709), .B1(new_n527), .B2(new_n655), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n706), .A2(new_n707), .A3(KEYINPUT94), .A4(new_n663), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n701), .B1(new_n712), .B2(new_n687), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT92), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n499), .A2(new_n500), .ZN(new_n716));
  INV_X1    g0516(.A(new_n573), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n717), .A2(new_n349), .A3(new_n549), .A4(new_n622), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(KEYINPUT30), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n565), .A2(new_n627), .A3(new_n571), .A4(new_n615), .ZN(new_n721));
  OAI21_X1  g0521(.A(KEYINPUT30), .B1(new_n721), .B2(new_n555), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT30), .ZN(new_n723));
  AOI22_X1  g0523(.A1(G264), .A2(new_n470), .B1(new_n626), .B2(new_n306), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n556), .A2(new_n723), .A3(new_n573), .A4(new_n724), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n722), .A2(new_n499), .A3(new_n725), .A4(new_n500), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n720), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n687), .B1(new_n727), .B2(KEYINPUT91), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT91), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n720), .A2(new_n729), .A3(new_n726), .ZN(new_n730));
  AOI21_X1  g0530(.A(KEYINPUT31), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n727), .A2(KEYINPUT31), .A3(new_n677), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n715), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  AND4_X1   g0534(.A1(new_n499), .A2(new_n722), .A3(new_n500), .A4(new_n725), .ZN(new_n735));
  AOI22_X1  g0535(.A1(new_n499), .A2(new_n500), .B1(new_n718), .B2(KEYINPUT30), .ZN(new_n736));
  OAI21_X1  g0536(.A(KEYINPUT91), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(new_n677), .A3(new_n730), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT31), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(KEYINPUT92), .A3(new_n732), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n637), .A2(new_n656), .A3(new_n658), .A4(new_n687), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n734), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G330), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n704), .A2(new_n714), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(new_n265), .ZN(new_n746));
  INV_X1    g0546(.A(new_n218), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G41), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n578), .A2(G116), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n749), .A2(G1), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(new_n211), .B2(new_n749), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT28), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n746), .A2(new_n753), .ZN(G364));
  NAND2_X1  g0554(.A1(new_n214), .A2(G13), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n265), .B1(new_n756), .B2(G45), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n748), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n683), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n760), .B1(G330), .B2(new_n681), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G13), .A2(G33), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n213), .B1(G20), .B2(new_n368), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n747), .A2(new_n337), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n769), .B1(new_n212), .B2(new_n465), .ZN(new_n770));
  INV_X1    g0570(.A(new_n249), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n770), .B1(new_n771), .B2(new_n465), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n747), .A2(new_n339), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n773), .A2(G355), .B1(new_n530), .B2(new_n747), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n767), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n765), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n214), .A2(new_n349), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n460), .A2(new_n324), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G326), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G190), .A2(G200), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G311), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n779), .A2(new_n780), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n460), .A2(G179), .A3(G200), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n214), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n784), .B1(G294), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT97), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n777), .A2(G190), .A3(new_n324), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n214), .A2(G179), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n778), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n791), .A2(G322), .B1(new_n794), .B2(G303), .ZN(new_n795));
  INV_X1    g0595(.A(G283), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n324), .A2(G190), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n792), .A2(new_n797), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n795), .B(new_n339), .C1(new_n796), .C2(new_n798), .ZN(new_n799));
  AND3_X1   g0599(.A1(new_n777), .A2(KEYINPUT96), .A3(new_n797), .ZN(new_n800));
  AOI21_X1  g0600(.A(KEYINPUT96), .B1(new_n777), .B2(new_n797), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(KEYINPUT33), .B(G317), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n799), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n792), .A2(new_n781), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n807), .A2(KEYINPUT98), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(KEYINPUT98), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G329), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n789), .A2(new_n805), .A3(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n786), .A2(new_n503), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n339), .B(new_n814), .C1(G87), .C2(new_n794), .ZN(new_n815));
  INV_X1    g0615(.A(G58), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n790), .A2(new_n816), .B1(new_n782), .B2(new_n204), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n779), .A2(new_n222), .B1(new_n798), .B2(new_n508), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n806), .A2(new_n396), .ZN(new_n820));
  XNOR2_X1  g0620(.A(KEYINPUT95), .B(KEYINPUT32), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n803), .A2(G68), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n815), .A2(new_n819), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n776), .B1(new_n813), .B2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n759), .ZN(new_n826));
  NOR3_X1   g0626(.A1(new_n775), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n764), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n827), .B1(new_n681), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n761), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(G396));
  NAND4_X1  g0631(.A1(new_n457), .A2(new_n454), .A3(new_n446), .A4(new_n677), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(KEYINPUT100), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT100), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n455), .A2(new_n834), .A3(new_n457), .A4(new_n677), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n454), .A2(new_n677), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n458), .A2(new_n461), .A3(new_n837), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(new_n700), .B2(new_n702), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT101), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n677), .B1(new_n836), .B2(new_n838), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n842), .B1(new_n669), .B2(new_n843), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n843), .B(new_n842), .C1(new_n696), .C2(new_n697), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  OR3_X1    g0647(.A1(new_n841), .A2(new_n847), .A3(new_n744), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n744), .B1(new_n841), .B2(new_n847), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n848), .A2(new_n826), .A3(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n765), .A2(new_n762), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n851), .B(KEYINPUT99), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n826), .B1(new_n853), .B2(new_n204), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n798), .A2(new_n203), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n337), .B1(new_n793), .B2(new_n222), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n855), .B(new_n856), .C1(G58), .C2(new_n787), .ZN(new_n857));
  INV_X1    g0657(.A(G132), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n857), .B1(new_n858), .B2(new_n810), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT34), .ZN(new_n860));
  INV_X1    g0660(.A(new_n779), .ZN(new_n861));
  INV_X1    g0661(.A(new_n782), .ZN(new_n862));
  AOI22_X1  g0662(.A1(G137), .A2(new_n861), .B1(new_n862), .B2(G159), .ZN(new_n863));
  INV_X1    g0663(.A(G143), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n863), .B1(new_n864), .B2(new_n790), .C1(new_n360), .C2(new_n802), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n859), .B1(new_n860), .B2(new_n865), .ZN(new_n866));
  OR2_X1    g0666(.A1(new_n865), .A2(new_n860), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n337), .B(new_n814), .C1(G303), .C2(new_n861), .ZN(new_n868));
  INV_X1    g0668(.A(new_n798), .ZN(new_n869));
  AOI22_X1  g0669(.A1(G116), .A2(new_n862), .B1(new_n869), .B2(G87), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n791), .A2(G294), .B1(new_n794), .B2(G107), .ZN(new_n871));
  AND3_X1   g0671(.A1(new_n868), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n811), .A2(G311), .B1(G283), .B2(new_n803), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n866), .A2(new_n867), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OAI221_X1 g0674(.A(new_n854), .B1(new_n776), .B2(new_n874), .C1(new_n840), .C2(new_n763), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n850), .A2(new_n875), .ZN(G384));
  OAI21_X1  g0676(.A(new_n464), .B1(new_n703), .B2(new_n713), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n646), .ZN(new_n878));
  XOR2_X1   g0678(.A(new_n878), .B(KEYINPUT104), .Z(new_n879));
  INV_X1    g0679(.A(KEYINPUT39), .ZN(new_n880));
  INV_X1    g0680(.A(new_n409), .ZN(new_n881));
  OR3_X1    g0681(.A1(new_n391), .A2(new_n397), .A3(KEYINPUT103), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT103), .B1(new_n391), .B2(new_n397), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n882), .A2(new_n387), .A3(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n391), .A2(new_n397), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n453), .B1(new_n885), .B2(KEYINPUT16), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n881), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n431), .B1(new_n887), .B2(new_n675), .ZN(new_n888));
  INV_X1    g0688(.A(new_n436), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(KEYINPUT37), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n675), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n410), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n437), .A2(new_n893), .A3(new_n431), .ZN(new_n894));
  OR2_X1    g0694(.A1(new_n894), .A2(KEYINPUT37), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n887), .A2(new_n675), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n643), .B2(new_n640), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n896), .A2(new_n898), .A3(KEYINPUT38), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n410), .B(new_n892), .C1(new_n643), .C2(new_n640), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n894), .B(KEYINPUT37), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT38), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n880), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n896), .A2(new_n898), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT38), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n907), .A2(KEYINPUT39), .A3(new_n899), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(G169), .B1(new_n312), .B2(new_n313), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(KEYINPUT14), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n911), .A2(new_n317), .A3(new_n314), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n912), .A2(new_n278), .A3(new_n687), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n909), .A2(new_n913), .B1(new_n439), .B2(new_n892), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n458), .A2(new_n677), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n843), .B1(new_n696), .B2(new_n697), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(KEYINPUT101), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n915), .B1(new_n917), .B2(new_n845), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n907), .A2(new_n899), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n278), .B(new_n677), .C1(new_n912), .C2(new_n641), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n278), .A2(new_n677), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n321), .A2(new_n326), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n918), .A2(new_n919), .A3(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n914), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n879), .B(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n900), .A2(new_n903), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n839), .B1(new_n920), .B2(new_n922), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n737), .A2(KEYINPUT31), .A3(new_n677), .A4(new_n730), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(KEYINPUT105), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT105), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n728), .A2(new_n933), .A3(KEYINPUT31), .A4(new_n730), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n932), .A2(new_n740), .A3(new_n934), .A4(new_n742), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n930), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(KEYINPUT40), .B1(new_n929), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT40), .B1(new_n907), .B2(new_n899), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n930), .A2(new_n935), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n464), .A2(new_n935), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n941), .A2(new_n942), .ZN(new_n944));
  INV_X1    g0744(.A(G330), .ZN(new_n945));
  NOR3_X1   g0745(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  OAI22_X1  g0746(.A1(new_n928), .A2(new_n946), .B1(new_n265), .B2(new_n756), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(new_n946), .B2(new_n928), .ZN(new_n948));
  INV_X1    g0748(.A(new_n506), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n949), .A2(KEYINPUT35), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(KEYINPUT35), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n950), .A2(G116), .A3(new_n215), .A4(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(KEYINPUT102), .B(KEYINPUT36), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n952), .B(new_n953), .ZN(new_n954));
  OR4_X1    g0754(.A1(new_n204), .A2(new_n211), .A3(new_n394), .A4(new_n393), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n222), .A2(G68), .ZN(new_n956));
  AOI211_X1 g0756(.A(new_n265), .B(G13), .C1(new_n955), .C2(new_n956), .ZN(new_n957));
  OR3_X1    g0757(.A1(new_n948), .A2(new_n954), .A3(new_n957), .ZN(G367));
  OAI211_X1 g0758(.A(new_n656), .B(new_n658), .C1(new_n518), .C2(new_n687), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n519), .A2(new_n677), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n961), .A2(new_n691), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n658), .B1(new_n959), .B2(new_n631), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n962), .A2(KEYINPUT42), .B1(new_n963), .B2(new_n687), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(KEYINPUT42), .B2(new_n962), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n649), .B1(new_n594), .B2(new_n687), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n594), .A2(new_n687), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n966), .B1(new_n663), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n965), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n971), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n961), .A2(new_n689), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n974), .A2(KEYINPUT106), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n972), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n974), .A2(KEYINPUT106), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n976), .B(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n691), .B1(new_n631), .B2(new_n677), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n961), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT45), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n961), .A2(new_n979), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT44), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n982), .B(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(new_n689), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n683), .A2(KEYINPUT107), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n691), .B1(new_n688), .B2(new_n690), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n987), .B(new_n988), .Z(new_n989));
  AOI21_X1  g0789(.A(new_n745), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n748), .B(KEYINPUT41), .Z(new_n991));
  OAI21_X1  g0791(.A(new_n757), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n978), .A2(new_n992), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n766), .B1(new_n218), .B2(new_n450), .C1(new_n243), .C2(new_n769), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n759), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT108), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n779), .A2(new_n864), .B1(new_n793), .B2(new_n816), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n339), .B(new_n997), .C1(G77), .C2(new_n869), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n786), .A2(new_n203), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n803), .A2(G159), .ZN(new_n1001));
  XOR2_X1   g0801(.A(KEYINPUT110), .B(G137), .Z(new_n1002));
  OAI22_X1  g0802(.A1(new_n790), .A2(new_n360), .B1(new_n1002), .B2(new_n806), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(G50), .B2(new_n862), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n998), .A2(new_n1000), .A3(new_n1001), .A4(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n544), .A2(new_n545), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n1006), .A2(new_n791), .B1(new_n861), .B2(G311), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT109), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n1007), .A2(new_n1008), .B1(new_n803), .B2(G294), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n794), .A2(G116), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT46), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1009), .B(new_n1011), .C1(new_n1008), .C2(new_n1007), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(G283), .A2(new_n862), .B1(new_n807), .B2(G317), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n337), .B1(new_n869), .B2(G97), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1013), .B(new_n1014), .C1(new_n508), .C2(new_n786), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1005), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT47), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n765), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n996), .B1(new_n1019), .B2(new_n1020), .C1(new_n968), .C2(new_n828), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n993), .A2(new_n1021), .ZN(G387));
  INV_X1    g0822(.A(new_n989), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n745), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n745), .A2(new_n1023), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1024), .A2(new_n748), .A3(new_n1025), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n790), .A2(new_n222), .B1(new_n793), .B2(new_n204), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n339), .B(new_n1027), .C1(G97), .C2(new_n869), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n786), .A2(new_n450), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n359), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n803), .A2(new_n1031), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n779), .A2(new_n396), .B1(new_n782), .B2(new_n203), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(G150), .B2(new_n807), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1028), .A2(new_n1030), .A3(new_n1032), .A4(new_n1034), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(G322), .A2(new_n861), .B1(new_n862), .B2(new_n1006), .ZN(new_n1036));
  INV_X1    g0836(.A(G317), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1036), .B1(new_n1037), .B2(new_n790), .C1(new_n802), .C2(new_n783), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT48), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n787), .A2(G283), .B1(new_n794), .B2(G294), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT111), .Z(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(KEYINPUT49), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n339), .B1(new_n806), .B2(new_n780), .C1(new_n530), .C2(new_n798), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT112), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1044), .A2(KEYINPUT49), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1035), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AND2_X1   g0850(.A1(new_n1050), .A2(new_n765), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n750), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n773), .A2(new_n1052), .B1(new_n508), .B2(new_n747), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n240), .A2(new_n465), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1031), .A2(new_n222), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT50), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n750), .A2(new_n465), .A3(new_n245), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n768), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1053), .B1(new_n1054), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n826), .B1(new_n1059), .B2(new_n766), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n688), .B2(new_n828), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1026), .B1(new_n757), .B2(new_n1023), .C1(new_n1051), .C2(new_n1061), .ZN(G393));
  NAND2_X1  g0862(.A1(new_n986), .A2(new_n758), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n961), .A2(new_n764), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n786), .A2(new_n204), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n339), .B(new_n1065), .C1(G87), .C2(new_n869), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n793), .A2(new_n203), .B1(new_n806), .B2(new_n864), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n1031), .B2(new_n862), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1066), .B(new_n1068), .C1(new_n222), .C2(new_n802), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n790), .A2(new_n396), .B1(new_n779), .B2(new_n360), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT51), .Z(new_n1071));
  OAI22_X1  g0871(.A1(new_n790), .A2(new_n783), .B1(new_n779), .B2(new_n1037), .ZN(new_n1072));
  XOR2_X1   g0872(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n1073));
  XNOR2_X1  g0873(.A(new_n1072), .B(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1006), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1074), .B1(new_n1075), .B2(new_n802), .ZN(new_n1076));
  INV_X1    g0876(.A(G322), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n782), .A2(new_n616), .B1(new_n806), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(G283), .B2(new_n794), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n337), .B1(new_n869), .B2(G107), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1079), .B(new_n1080), .C1(new_n530), .C2(new_n786), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n1069), .A2(new_n1071), .B1(new_n1076), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n765), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n253), .A2(new_n768), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n767), .B1(G97), .B2(new_n747), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n826), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1064), .A2(new_n1083), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1063), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n986), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1089), .A2(new_n1024), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1090), .A2(new_n749), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1089), .A2(new_n1024), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1088), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(G390));
  INV_X1    g0894(.A(KEYINPUT116), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n913), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n903), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1096), .B1(new_n1097), .B2(new_n899), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n677), .B1(new_n710), .B2(new_n711), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n915), .B1(new_n1099), .B2(new_n840), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1098), .B1(new_n1100), .B2(new_n924), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n743), .A2(G330), .A3(new_n923), .A4(new_n840), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n915), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n844), .B2(new_n846), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1096), .B1(new_n1104), .B2(new_n923), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n909), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1101), .B(new_n1102), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n913), .B1(new_n918), .B2(new_n924), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n677), .B(new_n839), .C1(new_n710), .C2(new_n711), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n923), .B1(new_n1109), .B2(new_n915), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1108), .A2(new_n909), .B1(new_n1110), .B2(new_n1098), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n930), .A2(new_n935), .A3(G330), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1107), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n330), .A2(new_n463), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n935), .A2(new_n1115), .A3(G330), .A4(new_n328), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT114), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n464), .A2(KEYINPUT114), .A3(G330), .A4(new_n935), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n877), .A2(new_n646), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n935), .A2(G330), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n839), .B1(new_n1122), .B2(KEYINPUT115), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT115), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n935), .A2(new_n1124), .A3(G330), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n923), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n733), .B1(new_n738), .B2(new_n739), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n742), .B1(new_n1128), .B2(KEYINPUT92), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n731), .A2(new_n715), .A3(new_n733), .ZN(new_n1130));
  OAI211_X1 g0930(.A(G330), .B(new_n840), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1112), .B1(new_n1131), .B2(new_n924), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n1126), .A2(new_n1127), .B1(new_n1132), .B2(new_n918), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1121), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1095), .B1(new_n1114), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n877), .A2(new_n646), .A3(new_n1120), .ZN(new_n1136));
  OR2_X1    g0936(.A1(new_n1132), .A2(new_n918), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1122), .A2(KEYINPUT115), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1138), .A2(new_n840), .A3(new_n1125), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n924), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1136), .B1(new_n1137), .B2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1101), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n1112), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1143), .A2(KEYINPUT116), .A3(new_n1107), .A4(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1135), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n749), .B1(new_n1114), .B2(new_n1134), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1114), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n909), .A2(new_n762), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n759), .B1(new_n852), .B2(new_n1031), .ZN(new_n1152));
  XOR2_X1   g0952(.A(new_n1152), .B(KEYINPUT117), .Z(new_n1153));
  NAND2_X1  g0953(.A1(new_n811), .A2(G125), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(KEYINPUT54), .B(G143), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n790), .A2(new_n858), .B1(new_n782), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(G50), .B2(new_n869), .ZN(new_n1157));
  INV_X1    g0957(.A(G128), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n337), .B1(new_n779), .B2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(G159), .B2(new_n787), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1002), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT53), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n793), .B2(new_n360), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n794), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n803), .A2(new_n1161), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1154), .A2(new_n1157), .A3(new_n1160), .A4(new_n1165), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n790), .A2(new_n530), .B1(new_n782), .B2(new_n503), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n855), .B(new_n1167), .C1(G283), .C2(new_n861), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n337), .B(new_n1065), .C1(G87), .C2(new_n794), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n810), .A2(new_n616), .B1(new_n508), .B2(new_n802), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1166), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1153), .B1(new_n1172), .B2(new_n765), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1150), .A2(new_n758), .B1(new_n1151), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1149), .A2(new_n1174), .ZN(G378));
  NAND2_X1  g0975(.A1(new_n367), .A2(new_n892), .ZN(new_n1176));
  XOR2_X1   g0976(.A(new_n386), .B(new_n1176), .Z(new_n1177));
  XNOR2_X1  g0977(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1177), .B(new_n1178), .Z(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1180), .A2(new_n941), .A3(G330), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1180), .B1(new_n941), .B2(G330), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n927), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n941), .A2(G330), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n1179), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1186), .A2(new_n926), .A3(new_n1181), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1184), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n758), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n759), .B1(new_n852), .B2(G50), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n1190), .B(KEYINPUT120), .Z(new_n1191));
  NOR2_X1   g0991(.A1(new_n337), .A2(G41), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n222), .B1(G33), .B2(G41), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n798), .A2(new_n816), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(G107), .B2(new_n791), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1196), .B1(new_n530), .B2(new_n779), .C1(new_n450), .C2(new_n782), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n810), .A2(new_n796), .B1(new_n503), .B2(new_n802), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1000), .B(new_n1192), .C1(new_n204), .C2(new_n793), .ZN(new_n1199));
  NOR3_X1   g0999(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1194), .B1(new_n1200), .B2(KEYINPUT58), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(KEYINPUT58), .B2(new_n1200), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n790), .A2(new_n1158), .B1(new_n793), .B2(new_n1155), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT118), .Z(new_n1204));
  NAND2_X1  g1004(.A1(new_n803), .A2(G132), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n787), .A2(G150), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(G125), .A2(new_n861), .B1(new_n862), .B2(G137), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  XOR2_X1   g1008(.A(new_n1208), .B(KEYINPUT59), .Z(new_n1209));
  OR2_X1    g1009(.A1(new_n1209), .A2(KEYINPUT119), .ZN(new_n1210));
  AOI211_X1 g1010(.A(G33), .B(G41), .C1(new_n869), .C2(G159), .ZN(new_n1211));
  INV_X1    g1011(.A(G124), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1211), .B1(new_n1212), .B2(new_n806), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n1209), .B2(KEYINPUT119), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1202), .B1(new_n1210), .B2(new_n1214), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n1191), .B1(new_n776), .B2(new_n1215), .C1(new_n1180), .C2(new_n763), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1189), .A2(KEYINPUT121), .A3(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT121), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n757), .B1(new_n1184), .B2(new_n1187), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1216), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1218), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1217), .A2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1147), .A2(new_n1121), .ZN(new_n1223));
  AOI21_X1  g1023(.A(KEYINPUT57), .B1(new_n1223), .B2(new_n1188), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1136), .B1(new_n1135), .B2(new_n1146), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1188), .A2(KEYINPUT57), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n748), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1222), .B1(new_n1224), .B2(new_n1227), .ZN(G375));
  NAND2_X1  g1028(.A1(new_n924), .A2(new_n762), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n337), .B1(new_n798), .B2(new_n816), .C1(new_n786), .C2(new_n222), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n779), .A2(new_n858), .B1(new_n793), .B2(new_n396), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n790), .A2(new_n1002), .B1(new_n782), .B2(new_n360), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1233), .B1(new_n1158), .B2(new_n810), .C1(new_n802), .C2(new_n1155), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n811), .A2(G303), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n779), .A2(new_n616), .B1(new_n793), .B2(new_n503), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n790), .A2(new_n796), .B1(new_n782), .B2(new_n508), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n337), .B(new_n1029), .C1(G77), .C2(new_n869), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n803), .A2(G116), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1235), .A2(new_n1238), .A3(new_n1239), .A4(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n776), .B1(new_n1234), .B2(new_n1241), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n826), .B(new_n1242), .C1(new_n203), .C2(new_n853), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n1133), .A2(new_n758), .B1(new_n1229), .B2(new_n1243), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n1143), .A2(new_n991), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1121), .A2(new_n1133), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1244), .B1(new_n1245), .B2(new_n1246), .ZN(G381));
  NOR3_X1   g1047(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1248));
  XOR2_X1   g1048(.A(new_n1248), .B(KEYINPUT122), .Z(new_n1249));
  NAND3_X1  g1049(.A1(new_n993), .A2(new_n1093), .A3(new_n1021), .ZN(new_n1250));
  NOR3_X1   g1050(.A1(new_n1249), .A2(G381), .A3(new_n1250), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(G375), .A2(G378), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(G407));
  NAND2_X1  g1053(.A1(new_n676), .A2(G213), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1252), .A2(new_n1255), .ZN(new_n1256));
  XOR2_X1   g1056(.A(new_n1256), .B(KEYINPUT123), .Z(new_n1257));
  NAND3_X1  g1057(.A1(new_n1257), .A2(G213), .A3(G407), .ZN(G409));
  INV_X1    g1058(.A(KEYINPUT61), .ZN(new_n1259));
  OAI211_X1 g1059(.A(G378), .B(new_n1222), .C1(new_n1224), .C2(new_n1227), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1149), .A2(new_n1174), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1188), .ZN(new_n1262));
  NOR3_X1   g1062(.A1(new_n1225), .A2(new_n991), .A3(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1189), .A2(new_n1216), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1261), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1255), .B1(new_n1260), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1246), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1134), .A2(KEYINPUT60), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1246), .A2(KEYINPUT60), .A3(new_n1134), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1269), .A2(new_n748), .A3(new_n1270), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(G384), .B(KEYINPUT124), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1271), .A2(new_n1244), .A3(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n1271), .A2(new_n1244), .B1(KEYINPUT124), .B2(G384), .ZN(new_n1275));
  OAI211_X1 g1075(.A(G2897), .B(new_n1255), .C1(new_n1274), .C2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1275), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1255), .A2(G2897), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1277), .A2(new_n1273), .A3(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1276), .A2(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1259), .B1(new_n1266), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(KEYINPUT126), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT126), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1283), .B(new_n1259), .C1(new_n1266), .C2(new_n1280), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1266), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(KEYINPUT62), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT62), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1266), .A2(new_n1288), .A3(new_n1285), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1282), .A2(new_n1284), .A3(new_n1287), .A4(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1093), .B1(new_n993), .B2(new_n1021), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(G393), .B(new_n830), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1292), .A2(new_n1250), .A3(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1250), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1293), .B1(new_n1296), .B2(new_n1291), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1290), .A2(new_n1298), .ZN(new_n1299));
  AND2_X1   g1099(.A1(new_n1266), .A2(new_n1285), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1298), .B1(new_n1300), .B2(KEYINPUT63), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1281), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT63), .ZN(new_n1303));
  AND3_X1   g1103(.A1(new_n1286), .A2(KEYINPUT125), .A3(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(KEYINPUT125), .B1(new_n1286), .B2(new_n1303), .ZN(new_n1305));
  OAI211_X1 g1105(.A(new_n1301), .B(new_n1302), .C1(new_n1304), .C2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1299), .A2(new_n1306), .ZN(G405));
  NAND2_X1  g1107(.A1(G375), .A2(new_n1261), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(new_n1260), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n1285), .ZN(new_n1310));
  OAI211_X1 g1110(.A(new_n1308), .B(new_n1260), .C1(new_n1274), .C2(new_n1275), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT127), .ZN(new_n1312));
  OAI211_X1 g1112(.A(new_n1310), .B(new_n1311), .C1(new_n1298), .C2(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(KEYINPUT127), .B1(new_n1295), .B2(new_n1297), .ZN(new_n1314));
  XNOR2_X1  g1114(.A(new_n1313), .B(new_n1314), .ZN(G402));
endmodule


