//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 0 1 0 1 1 0 1 0 0 0 1 1 1 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n561, new_n563, new_n564, new_n565,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n621, new_n622, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT64), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  AOI22_X1  g035(.A1(new_n460), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT65), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(new_n460), .A3(G137), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n467), .A2(new_n472), .ZN(G160));
  OAI221_X1 g048(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n466), .C2(G112), .ZN(new_n474));
  INV_X1    g049(.A(G136), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n460), .A2(new_n462), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  XNOR2_X1  g052(.A(KEYINPUT65), .B(G2105), .ZN(new_n478));
  AND3_X1   g053(.A1(new_n460), .A2(new_n478), .A3(KEYINPUT66), .ZN(new_n479));
  AOI21_X1  g054(.A(KEYINPUT66), .B1(new_n460), .B2(new_n478), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n477), .B1(new_n482), .B2(G124), .ZN(G162));
  OR2_X1    g058(.A1(G102), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G114), .C2(new_n462), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n486));
  AND2_X1   g061(.A1(G126), .A2(G2105), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(new_n460), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT3), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2104), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n489), .A2(new_n491), .A3(new_n487), .A4(new_n486), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n485), .B1(new_n488), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT68), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT69), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(KEYINPUT4), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n466), .A2(new_n460), .A3(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n501), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n466), .A2(new_n460), .A3(new_n503), .A4(new_n499), .ZN(new_n504));
  AND2_X1   g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n489), .A2(new_n491), .A3(new_n487), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT67), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(new_n492), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT68), .A3(new_n485), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n496), .A2(new_n505), .A3(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G164));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  OAI21_X1  g089(.A(KEYINPUT5), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n516), .A2(KEYINPUT70), .A3(G543), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G62), .ZN(new_n519));
  NAND2_X1  g094(.A1(G75), .A2(G543), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n512), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n524), .A2(new_n514), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G50), .ZN(new_n526));
  OAI211_X1 g101(.A(new_n515), .B(new_n517), .C1(new_n523), .C2(new_n522), .ZN(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT71), .B(G88), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n521), .A2(new_n529), .ZN(G166));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  INV_X1    g107(.A(G89), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n527), .B2(new_n533), .ZN(new_n534));
  XOR2_X1   g109(.A(new_n534), .B(KEYINPUT72), .Z(new_n535));
  NAND3_X1  g110(.A1(new_n518), .A2(G63), .A3(G651), .ZN(new_n536));
  INV_X1    g111(.A(G51), .ZN(new_n537));
  INV_X1    g112(.A(new_n525), .ZN(new_n538));
  OAI211_X1 g113(.A(new_n535), .B(new_n536), .C1(new_n537), .C2(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n515), .A2(new_n517), .ZN(new_n542));
  INV_X1    g117(.A(G64), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(KEYINPUT73), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(KEYINPUT73), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n545), .A2(G651), .A3(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n527), .ZN(new_n548));
  XOR2_X1   g123(.A(KEYINPUT74), .B(G52), .Z(new_n549));
  AOI22_X1  g124(.A1(new_n548), .A2(G90), .B1(new_n525), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(G171));
  NAND2_X1  g127(.A1(new_n518), .A2(G56), .ZN(new_n553));
  NAND2_X1  g128(.A1(G68), .A2(G543), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n512), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n525), .A2(G43), .ZN(new_n556));
  INV_X1    g131(.A(G81), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n557), .B2(new_n527), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  AND3_X1   g135(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G36), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT75), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n561), .A2(new_n565), .ZN(G188));
  NAND2_X1  g141(.A1(new_n525), .A2(G53), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT9), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n548), .A2(KEYINPUT76), .A3(G91), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT76), .ZN(new_n570));
  INV_X1    g145(.A(G91), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n527), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n518), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n574));
  OR2_X1    g149(.A1(new_n574), .A2(new_n512), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n568), .A2(new_n573), .A3(new_n575), .ZN(G299));
  INV_X1    g151(.A(KEYINPUT77), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n551), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n551), .A2(new_n577), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G301));
  INV_X1    g157(.A(G166), .ZN(G303));
  NAND2_X1  g158(.A1(new_n548), .A2(G87), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n585));
  INV_X1    g160(.A(G49), .ZN(new_n586));
  OAI211_X1 g161(.A(new_n584), .B(new_n585), .C1(new_n586), .C2(new_n538), .ZN(G288));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n542), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(G651), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n548), .A2(G86), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n525), .A2(G48), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT78), .ZN(G305));
  NAND2_X1  g170(.A1(new_n518), .A2(G60), .ZN(new_n596));
  NAND2_X1  g171(.A1(G72), .A2(G543), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n512), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n525), .A2(G47), .ZN(new_n599));
  INV_X1    g174(.A(G85), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n600), .B2(new_n527), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(new_n548), .A2(G92), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT10), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n604), .B(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT79), .ZN(new_n608));
  INV_X1    g183(.A(G66), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n542), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G651), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n525), .A2(G54), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n606), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(new_n581), .B2(new_n614), .ZN(G284));
  OAI21_X1  g191(.A(new_n615), .B1(new_n581), .B2(new_n614), .ZN(G321));
  NAND2_X1  g192(.A1(G299), .A2(new_n614), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(G168), .B2(new_n614), .ZN(G297));
  OAI21_X1  g194(.A(new_n618), .B1(G168), .B2(new_n614), .ZN(G280));
  AND3_X1   g195(.A1(new_n606), .A2(new_n611), .A3(new_n612), .ZN(new_n621));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(G860), .ZN(G148));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G868), .B2(new_n559), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n460), .A2(new_n470), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2100), .ZN(new_n631));
  OAI221_X1 g206(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n466), .C2(G111), .ZN(new_n632));
  INV_X1    g207(.A(G135), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(new_n633), .B2(new_n476), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n634), .B1(new_n482), .B2(G123), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2096), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n631), .A2(new_n636), .ZN(G156));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2438), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2427), .B(G2430), .Z(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT14), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n644), .A2(KEYINPUT81), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(KEYINPUT81), .ZN(new_n646));
  NAND4_X1  g221(.A1(new_n642), .A2(new_n643), .A3(new_n645), .A4(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2443), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2446), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n649), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n653), .B(new_n654), .Z(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(G14), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G401));
  XNOR2_X1  g232(.A(G2072), .B(G2078), .ZN(new_n658));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT82), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT18), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n658), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT83), .ZN(new_n666));
  XOR2_X1   g241(.A(G2096), .B(G2100), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n662), .A2(KEYINPUT17), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n660), .A2(new_n661), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n664), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n668), .B(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(G227));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n680));
  INV_X1    g255(.A(new_n675), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n676), .A2(new_n677), .ZN(new_n682));
  AOI22_X1  g257(.A1(new_n679), .A2(new_n680), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n682), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n684), .A2(new_n675), .A3(new_n678), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n683), .B(new_n685), .C1(new_n679), .C2(new_n680), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT86), .ZN(new_n687));
  INV_X1    g262(.A(G1996), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT85), .B(G1986), .Z(new_n690));
  XNOR2_X1  g265(.A(G1981), .B(G1991), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n689), .B(new_n694), .Z(G229));
  XNOR2_X1  g270(.A(KEYINPUT89), .B(G16), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G24), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(new_n602), .B2(new_n697), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(G1986), .ZN(new_n700));
  MUX2_X1   g275(.A(G6), .B(G305), .S(G16), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT32), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n702), .A2(G1981), .ZN(new_n703));
  INV_X1    g278(.A(G22), .ZN(new_n704));
  OAI21_X1  g279(.A(KEYINPUT92), .B1(new_n696), .B2(new_n704), .ZN(new_n705));
  OR3_X1    g280(.A1(new_n696), .A2(KEYINPUT92), .A3(new_n704), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n705), .B(new_n706), .C1(G166), .C2(new_n697), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n707), .A2(G1971), .ZN(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G23), .ZN(new_n710));
  INV_X1    g285(.A(G288), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(new_n709), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT90), .B(KEYINPUT91), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n712), .B(new_n713), .Z(new_n714));
  XOR2_X1   g289(.A(KEYINPUT33), .B(G1976), .Z(new_n715));
  AND2_X1   g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n714), .A2(new_n715), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n707), .A2(G1971), .ZN(new_n718));
  NOR3_X1   g293(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n702), .A2(G1981), .ZN(new_n720));
  NAND4_X1  g295(.A1(new_n703), .A2(new_n708), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  AOI211_X1 g296(.A(KEYINPUT93), .B(new_n700), .C1(new_n721), .C2(KEYINPUT34), .ZN(new_n722));
  INV_X1    g297(.A(new_n476), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n482), .A2(G119), .B1(G131), .B2(new_n723), .ZN(new_n724));
  OAI221_X1 g299(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n466), .C2(G107), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT87), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  MUX2_X1   g302(.A(G25), .B(new_n727), .S(G29), .Z(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT35), .B(G1991), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT88), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n728), .B(new_n730), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n722), .B(new_n731), .C1(KEYINPUT34), .C2(new_n721), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT36), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n723), .A2(G141), .B1(G105), .B2(new_n470), .ZN(new_n735));
  NAND3_X1  g310(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT26), .Z(new_n737));
  INV_X1    g312(.A(G129), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n735), .B(new_n737), .C1(new_n481), .C2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT97), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT98), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  MUX2_X1   g318(.A(G32), .B(new_n743), .S(G29), .Z(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT27), .B(G1996), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n732), .A2(new_n733), .ZN(new_n747));
  INV_X1    g322(.A(G29), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G26), .ZN(new_n749));
  OAI221_X1 g324(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n466), .C2(G116), .ZN(new_n750));
  INV_X1    g325(.A(G140), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n750), .B1(new_n751), .B2(new_n476), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n482), .B2(G128), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT96), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n749), .B1(new_n756), .B2(new_n748), .ZN(new_n757));
  MUX2_X1   g332(.A(new_n749), .B(new_n757), .S(KEYINPUT28), .Z(new_n758));
  INV_X1    g333(.A(G2067), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(KEYINPUT99), .B1(G5), .B2(G16), .ZN(new_n761));
  OR3_X1    g336(.A1(KEYINPUT99), .A2(G5), .A3(G16), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n761), .B(new_n762), .C1(new_n551), .C2(new_n709), .ZN(new_n763));
  INV_X1    g338(.A(G1961), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n748), .A2(G27), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G164), .B2(new_n748), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(G2078), .Z(new_n768));
  NAND3_X1  g343(.A1(new_n760), .A2(new_n765), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n709), .A2(G21), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G168), .B2(new_n709), .ZN(new_n771));
  INV_X1    g346(.A(G1966), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT30), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n748), .B1(new_n774), .B2(G28), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n774), .B2(G28), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n763), .A2(new_n764), .ZN(new_n777));
  AOI211_X1 g352(.A(new_n776), .B(new_n777), .C1(G29), .C2(new_n635), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT31), .B(G11), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n773), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT100), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n621), .A2(new_n709), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G4), .B2(new_n709), .ZN(new_n783));
  INV_X1    g358(.A(G1348), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n748), .A2(G33), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT25), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n723), .A2(G139), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n787), .B(new_n788), .C1(new_n466), .C2(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n785), .B1(new_n790), .B2(G29), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n783), .A2(new_n784), .B1(new_n792), .B2(G2072), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G2072), .B2(new_n792), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n559), .A2(new_n697), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT94), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n697), .A2(G19), .ZN(new_n797));
  NOR3_X1   g372(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n796), .B2(new_n797), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT95), .B(G1341), .Z(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n794), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n697), .A2(KEYINPUT23), .A3(G20), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT23), .ZN(new_n804));
  INV_X1    g379(.A(G20), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n696), .B2(new_n805), .ZN(new_n806));
  AND3_X1   g381(.A1(new_n568), .A2(new_n573), .A3(new_n575), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n803), .B(new_n806), .C1(new_n807), .C2(new_n709), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT101), .B(G1956), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n783), .A2(new_n784), .ZN(new_n811));
  OR2_X1    g386(.A1(KEYINPUT24), .A2(G34), .ZN(new_n812));
  NAND2_X1  g387(.A1(KEYINPUT24), .A2(G34), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n812), .A2(new_n748), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(G160), .B2(new_n748), .ZN(new_n815));
  AOI211_X1 g390(.A(new_n810), .B(new_n811), .C1(G2084), .C2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n748), .A2(G35), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G162), .B2(new_n748), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT29), .B(G2090), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n802), .A2(new_n816), .A3(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n815), .A2(G2084), .ZN(new_n822));
  NOR4_X1   g397(.A1(new_n769), .A2(new_n781), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n734), .A2(new_n746), .A3(new_n747), .A4(new_n823), .ZN(G150));
  INV_X1    g399(.A(G150), .ZN(G311));
  NAND2_X1  g400(.A1(new_n525), .A2(G55), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT102), .B(G93), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n518), .A2(G67), .ZN(new_n828));
  NAND2_X1  g403(.A1(G80), .A2(G543), .ZN(new_n829));
  AND2_X1   g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OAI221_X1 g405(.A(new_n826), .B1(new_n527), .B2(new_n827), .C1(new_n830), .C2(new_n512), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(G860), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT37), .Z(new_n833));
  OR2_X1    g408(.A1(new_n831), .A2(new_n559), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n831), .A2(new_n559), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT39), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n621), .A2(G559), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT38), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n837), .B(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n833), .B1(new_n840), .B2(G860), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT103), .ZN(G145));
  XNOR2_X1  g417(.A(new_n755), .B(new_n741), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n502), .A2(new_n508), .A3(new_n504), .A4(new_n485), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n843), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT105), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n790), .B2(KEYINPUT98), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n790), .A2(new_n847), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n850), .A2(new_n848), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n849), .B1(new_n846), .B2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n727), .B(new_n629), .ZN(new_n853));
  OAI221_X1 g428(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n466), .C2(G118), .ZN(new_n854));
  INV_X1    g429(.A(G142), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n854), .B1(new_n855), .B2(new_n476), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(new_n482), .B2(G130), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n853), .B(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n852), .B(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(G162), .B(KEYINPUT104), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(G160), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(new_n635), .Z(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(G37), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n859), .A2(new_n863), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(KEYINPUT40), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT40), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n864), .A2(new_n869), .A3(new_n865), .A4(new_n866), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(G395));
  NAND2_X1  g446(.A1(new_n831), .A2(new_n614), .ZN(new_n872));
  OR3_X1    g447(.A1(new_n613), .A2(new_n807), .A3(KEYINPUT106), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT106), .B1(new_n613), .B2(new_n807), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT107), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(new_n621), .B2(G299), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n613), .A2(new_n807), .A3(KEYINPUT107), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n836), .B(new_n624), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT41), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n875), .A2(KEYINPUT41), .A3(new_n879), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n883), .B1(new_n887), .B2(new_n882), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT42), .ZN(new_n889));
  XNOR2_X1  g464(.A(G166), .B(G288), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(G305), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(new_n602), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n892), .A2(KEYINPUT108), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n889), .B(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n872), .B1(new_n894), .B2(new_n614), .ZN(G295));
  OAI21_X1  g470(.A(new_n872), .B1(new_n894), .B2(new_n614), .ZN(G331));
  INV_X1    g471(.A(new_n580), .ZN(new_n897));
  AOI21_X1  g472(.A(G286), .B1(new_n897), .B2(new_n578), .ZN(new_n898));
  NAND2_X1  g473(.A1(G286), .A2(G171), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n835), .B(new_n834), .C1(new_n898), .C2(new_n900), .ZN(new_n901));
  OAI211_X1 g476(.A(new_n836), .B(new_n899), .C1(new_n581), .C2(G286), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n885), .A2(new_n886), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n902), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n881), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n892), .ZN(new_n907));
  INV_X1    g482(.A(new_n892), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n903), .A2(new_n908), .A3(new_n905), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n907), .A2(new_n865), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(KEYINPUT43), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n907), .A2(new_n912), .A3(new_n865), .A4(new_n909), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT109), .ZN(new_n915));
  OAI21_X1  g490(.A(KEYINPUT110), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n917), .B1(new_n914), .B2(new_n915), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT110), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n911), .A2(KEYINPUT109), .A3(new_n919), .A4(new_n913), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n916), .A2(new_n918), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n918), .B1(new_n916), .B2(new_n920), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(G397));
  INV_X1    g498(.A(G1384), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n502), .A2(new_n504), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n924), .B1(new_n925), .B2(new_n494), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT45), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(G160), .A2(G40), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n743), .A2(G1996), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n755), .B(G2067), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n741), .A2(G1996), .A3(new_n930), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(KEYINPUT111), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT112), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n936), .B(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n930), .ZN(new_n939));
  INV_X1    g514(.A(new_n729), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n727), .B(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n939), .B1(new_n942), .B2(KEYINPUT113), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n943), .B1(KEYINPUT113), .B2(new_n942), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n602), .B(G1986), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n938), .B(new_n944), .C1(new_n939), .C2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT114), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n946), .B(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G8), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n929), .A2(new_n926), .ZN(new_n950));
  AOI211_X1 g525(.A(new_n949), .B(new_n950), .C1(G1976), .C2(new_n711), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT52), .ZN(new_n952));
  OR2_X1    g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n951), .B(new_n952), .C1(G1976), .C2(new_n711), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n594), .B(KEYINPUT49), .ZN(new_n955));
  INV_X1    g530(.A(G1981), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n956), .B1(new_n591), .B2(KEYINPUT117), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n955), .B(new_n957), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n950), .A2(new_n949), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AND3_X1   g535(.A1(new_n953), .A2(new_n954), .A3(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(KEYINPUT118), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n510), .A2(new_n924), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n927), .ZN(new_n964));
  INV_X1    g539(.A(G40), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n467), .A2(new_n472), .A3(new_n965), .ZN(new_n966));
  OAI211_X1 g541(.A(KEYINPUT45), .B(new_n924), .C1(new_n925), .C2(new_n494), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT115), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n844), .A2(KEYINPUT115), .A3(KEYINPUT45), .A4(new_n924), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n964), .A2(new_n966), .A3(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n973), .A2(G1971), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n963), .A2(KEYINPUT50), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT50), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n844), .A2(new_n976), .A3(new_n924), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n975), .A2(new_n966), .A3(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n978), .A2(G2090), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n974), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n980), .A2(new_n949), .ZN(new_n981));
  NOR2_X1   g556(.A1(G166), .A2(new_n949), .ZN(new_n982));
  XOR2_X1   g557(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT55), .ZN(new_n985));
  OAI22_X1  g560(.A1(G166), .A2(new_n949), .B1(KEYINPUT116), .B2(new_n985), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n981), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n510), .A2(new_n976), .A3(new_n924), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n926), .A2(KEYINPUT50), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n990), .A2(new_n966), .A3(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n992), .A2(G2090), .ZN(new_n993));
  OAI21_X1  g568(.A(G8), .B1(new_n974), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n987), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n962), .A2(new_n989), .A3(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n996), .B(KEYINPUT125), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT122), .ZN(new_n998));
  INV_X1    g573(.A(G1956), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n992), .A2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g575(.A(KEYINPUT56), .B(G2072), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n964), .A2(new_n971), .A3(new_n966), .A4(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT57), .ZN(new_n1003));
  XNOR2_X1  g578(.A(G299), .B(new_n1003), .ZN(new_n1004));
  AND3_X1   g579(.A1(new_n1000), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1004), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT61), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1004), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT61), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1000), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1007), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT121), .ZN(new_n1015));
  XOR2_X1   g590(.A(KEYINPUT58), .B(G1341), .Z(new_n1016));
  OAI21_X1  g591(.A(new_n1016), .B1(new_n929), .B2(new_n926), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1017), .B1(new_n972), .B2(G1996), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n559), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT59), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT59), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1018), .A2(new_n1021), .A3(new_n559), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n1014), .A2(new_n1015), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1015), .B1(new_n1014), .B2(new_n1023), .ZN(new_n1025));
  AOI22_X1  g600(.A1(new_n978), .A2(new_n784), .B1(new_n759), .B2(new_n950), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1026), .B1(KEYINPUT60), .B2(new_n621), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n621), .A2(KEYINPUT60), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n1027), .B(new_n1029), .ZN(new_n1030));
  NOR3_X1   g605(.A1(new_n1024), .A2(new_n1025), .A3(new_n1030), .ZN(new_n1031));
  OR3_X1    g606(.A1(new_n1005), .A2(new_n613), .A3(new_n1026), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n1010), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n998), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1035), .B1(new_n972), .B2(G2078), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n978), .A2(new_n764), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT119), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n928), .A2(new_n1039), .A3(new_n966), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT45), .B1(new_n844), .B2(new_n924), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT119), .B1(new_n1041), .B2(new_n929), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n510), .A2(KEYINPUT45), .A3(new_n924), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1040), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  OR3_X1    g619(.A1(new_n1044), .A2(new_n1035), .A3(G2078), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1038), .A2(G301), .A3(new_n1045), .ZN(new_n1046));
  NOR3_X1   g621(.A1(new_n1041), .A2(new_n1035), .A3(G2078), .ZN(new_n1047));
  INV_X1    g622(.A(new_n467), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n468), .A2(KEYINPUT124), .A3(new_n471), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT124), .B1(new_n468), .B2(new_n471), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n1049), .A2(new_n1050), .A3(new_n965), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1047), .A2(new_n971), .A3(new_n1048), .A4(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1036), .A2(new_n1037), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(G171), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n1046), .A2(KEYINPUT54), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1038), .A2(new_n1045), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n581), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1038), .A2(G301), .A3(new_n1052), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT54), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT51), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1044), .A2(new_n772), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT120), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(G2084), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n975), .A2(new_n1064), .A3(new_n966), .A4(new_n977), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1044), .A2(KEYINPUT120), .A3(new_n772), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1063), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1060), .B1(new_n1067), .B2(G286), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1063), .A2(G168), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(G8), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1060), .B1(new_n1069), .B2(G8), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT123), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1070), .A2(KEYINPUT51), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT123), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1074), .B(new_n1075), .C1(new_n1070), .C2(new_n1068), .ZN(new_n1076));
  AOI211_X1 g651(.A(new_n1055), .B(new_n1059), .C1(new_n1073), .C2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1033), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1014), .A2(new_n1023), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT121), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1014), .A2(new_n1015), .A3(new_n1023), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(KEYINPUT122), .B(new_n1078), .C1(new_n1082), .C2(new_n1030), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1034), .A2(new_n1077), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT62), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT62), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1073), .A2(new_n1087), .A3(new_n1076), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1086), .A2(new_n581), .A3(new_n1056), .A4(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n997), .B1(new_n1084), .B2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n981), .A2(new_n961), .A3(new_n988), .ZN(new_n1091));
  AOI211_X1 g666(.A(G1976), .B(G288), .C1(new_n958), .C2(new_n959), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n594), .A2(G1981), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n959), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n996), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1067), .ZN(new_n1096));
  NOR3_X1   g671(.A1(new_n1096), .A2(new_n949), .A3(G286), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT63), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n987), .B1(new_n980), .B2(new_n949), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n989), .A2(KEYINPUT63), .A3(new_n961), .A4(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1097), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1091), .B(new_n1094), .C1(new_n1098), .C2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n948), .B1(new_n1090), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n930), .B1(new_n932), .B2(new_n741), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n930), .A2(new_n688), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1106), .B(KEYINPUT46), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  XOR2_X1   g683(.A(new_n1108), .B(KEYINPUT47), .Z(new_n1109));
  NAND4_X1  g684(.A1(new_n938), .A2(new_n726), .A3(new_n724), .A4(new_n940), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n756), .A2(new_n759), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n939), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n938), .A2(new_n944), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n939), .A2(G1986), .A3(G290), .ZN(new_n1114));
  XOR2_X1   g689(.A(new_n1114), .B(KEYINPUT126), .Z(new_n1115));
  XNOR2_X1  g690(.A(new_n1115), .B(KEYINPUT48), .ZN(new_n1116));
  AOI211_X1 g691(.A(new_n1109), .B(new_n1112), .C1(new_n1113), .C2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1104), .A2(new_n1117), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g693(.A(G229), .ZN(new_n1120));
  NAND3_X1  g694(.A1(new_n656), .A2(G319), .A3(new_n672), .ZN(new_n1121));
  INV_X1    g695(.A(KEYINPUT127), .ZN(new_n1122));
  OAI21_X1  g696(.A(new_n1120), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g697(.A(new_n1123), .B1(new_n1122), .B2(new_n1121), .ZN(new_n1124));
  NAND3_X1  g698(.A1(new_n867), .A2(new_n914), .A3(new_n1124), .ZN(G225));
  INV_X1    g699(.A(G225), .ZN(G308));
endmodule


