//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 0 0 1 0 0 1 0 0 1 0 0 1 0 1 0 1 0 0 0 1 0 0 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 0 1 1 0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1037, new_n1038, new_n1039, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083, new_n1084, new_n1085,
    new_n1086, new_n1087, new_n1088, new_n1089, new_n1090, new_n1091;
  INV_X1    g000(.A(KEYINPUT95), .ZN(new_n187));
  OAI21_X1  g001(.A(G214), .B1(G237), .B2(G902), .ZN(new_n188));
  NAND2_X1  g002(.A1(G234), .A2(G237), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(G952), .A3(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  XOR2_X1   g006(.A(KEYINPUT21), .B(G898), .Z(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n189), .A2(G902), .A3(G953), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n192), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G104), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT3), .B1(new_n199), .B2(G107), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n201));
  INV_X1    g015(.A(G107), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G104), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n199), .A2(G107), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n200), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G101), .ZN(new_n206));
  INV_X1    g020(.A(G101), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n200), .A2(new_n203), .A3(new_n207), .A4(new_n204), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n206), .A2(KEYINPUT4), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT4), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n205), .A2(new_n210), .A3(G101), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G116), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(G119), .ZN(new_n214));
  INV_X1    g028(.A(G119), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT64), .B1(new_n215), .B2(G116), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT64), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(new_n213), .A3(G119), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n214), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT2), .B(G113), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n219), .B(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT79), .B1(new_n212), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n220), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n219), .B(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT79), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n224), .A2(new_n225), .A3(new_n209), .A4(new_n211), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n222), .A2(new_n226), .ZN(new_n227));
  XOR2_X1   g041(.A(G110), .B(G122), .Z(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(G104), .B(G107), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT75), .B1(new_n230), .B2(new_n207), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT75), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n202), .A2(G104), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n199), .A2(G107), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n232), .B(G101), .C1(new_n233), .C2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n231), .A2(new_n208), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT76), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT76), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n231), .A2(new_n238), .A3(new_n235), .A4(new_n208), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT80), .B(KEYINPUT5), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n219), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G113), .ZN(new_n243));
  XOR2_X1   g057(.A(KEYINPUT80), .B(KEYINPUT5), .Z(new_n244));
  AOI21_X1  g058(.A(new_n243), .B1(new_n244), .B2(new_n214), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n242), .A2(new_n245), .B1(new_n219), .B2(new_n223), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n240), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n227), .A2(KEYINPUT82), .A3(new_n229), .A4(new_n247), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n247), .A2(new_n222), .A3(new_n229), .A4(new_n226), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT82), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G146), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G143), .ZN(new_n254));
  INV_X1    g068(.A(G143), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G146), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(KEYINPUT0), .A2(G128), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n257), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n254), .A2(new_n256), .A3(new_n258), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(G125), .A3(new_n262), .ZN(new_n263));
  OR2_X1    g077(.A1(new_n263), .A2(KEYINPUT83), .ZN(new_n264));
  INV_X1    g078(.A(G128), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(KEYINPUT1), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(new_n254), .A3(new_n256), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n265), .A2(new_n253), .A3(G143), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n255), .B(G146), .C1(new_n265), .C2(KEYINPUT1), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n263), .B(KEYINPUT83), .C1(G125), .C2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G224), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n272), .A2(G953), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n264), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n264), .A2(new_n271), .ZN(new_n275));
  INV_X1    g089(.A(new_n273), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n275), .A2(KEYINPUT7), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n214), .ZN(new_n278));
  OAI21_X1  g092(.A(G113), .B1(new_n241), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n279), .B1(KEYINPUT5), .B2(new_n219), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n219), .A2(new_n223), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NOR3_X1   g096(.A1(new_n280), .A2(new_n282), .A3(new_n236), .ZN(new_n283));
  INV_X1    g097(.A(new_n236), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT85), .B1(new_n246), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT85), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n279), .B1(new_n219), .B2(new_n241), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n286), .B(new_n236), .C1(new_n287), .C2(new_n282), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n283), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  XOR2_X1   g103(.A(KEYINPUT84), .B(KEYINPUT8), .Z(new_n290));
  XNOR2_X1  g104(.A(new_n228), .B(new_n290), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n274), .B(new_n277), .C1(new_n289), .C2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n275), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT7), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n252), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G902), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n275), .A2(new_n276), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n274), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n247), .A2(new_n222), .A3(new_n226), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT6), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n304), .A2(KEYINPUT81), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n303), .A2(new_n228), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n305), .B1(new_n303), .B2(new_n228), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n248), .A2(KEYINPUT6), .A3(new_n251), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n302), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(G210), .B1(G237), .B2(G902), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n299), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n248), .A2(KEYINPUT6), .A3(new_n251), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n303), .A2(new_n228), .ZN(new_n315));
  INV_X1    g129(.A(new_n305), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n303), .A2(new_n228), .A3(new_n305), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n301), .B1(new_n314), .B2(new_n319), .ZN(new_n320));
  AOI22_X1  g134(.A1(new_n248), .A2(new_n251), .B1(new_n295), .B2(new_n294), .ZN(new_n321));
  AOI21_X1  g135(.A(G902), .B1(new_n321), .B2(new_n293), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n311), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n188), .B(new_n198), .C1(new_n313), .C2(new_n323), .ZN(new_n324));
  NOR2_X1   g138(.A1(G237), .A2(G953), .ZN(new_n325));
  AND3_X1   g139(.A1(new_n325), .A2(G143), .A3(G214), .ZN(new_n326));
  AOI21_X1  g140(.A(G143), .B1(new_n325), .B2(G214), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n326), .A2(new_n327), .A3(G131), .ZN(new_n328));
  INV_X1    g142(.A(G131), .ZN(new_n329));
  INV_X1    g143(.A(G237), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(new_n190), .A3(G214), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n255), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n325), .A2(G143), .A3(G214), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n329), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OR3_X1    g148(.A1(new_n328), .A2(new_n334), .A3(KEYINPUT17), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT16), .ZN(new_n336));
  INV_X1    g150(.A(G125), .ZN(new_n337));
  INV_X1    g151(.A(G140), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(G125), .A2(G140), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n336), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n336), .A2(new_n338), .A3(G125), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n253), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  AND2_X1   g158(.A1(G125), .A2(G140), .ZN(new_n345));
  NOR2_X1   g159(.A1(G125), .A2(G140), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT16), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(G146), .A3(new_n342), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n344), .A2(KEYINPUT71), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT71), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n350), .B(new_n253), .C1(new_n341), .C2(new_n343), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n334), .A2(KEYINPUT17), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n335), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(KEYINPUT18), .A2(G131), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n356), .B1(new_n326), .B2(new_n327), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(KEYINPUT86), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n332), .A2(new_n333), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT86), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n360), .A3(new_n356), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n332), .A2(new_n333), .A3(new_n355), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n253), .B1(new_n345), .B2(new_n346), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n339), .A2(G146), .A3(new_n340), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n358), .A2(new_n361), .A3(new_n362), .A4(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n354), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(G113), .B(G122), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n368), .B(new_n199), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n354), .A2(new_n369), .A3(new_n366), .ZN(new_n372));
  AOI21_X1  g186(.A(G902), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G475), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(G475), .A2(G902), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT87), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n360), .B1(new_n359), .B2(new_n356), .ZN(new_n378));
  AOI211_X1 g192(.A(KEYINPUT86), .B(new_n355), .C1(new_n332), .C2(new_n333), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n362), .A2(new_n365), .ZN(new_n380));
  NOR3_X1   g194(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT19), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n382), .B1(new_n345), .B2(new_n346), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n339), .A2(KEYINPUT19), .A3(new_n340), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(new_n253), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n348), .ZN(new_n386));
  INV_X1    g200(.A(new_n328), .ZN(new_n387));
  INV_X1    g201(.A(new_n334), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n377), .B1(new_n381), .B2(new_n389), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n348), .B(new_n385), .C1(new_n328), .C2(new_n334), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n366), .A2(KEYINPUT87), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(new_n370), .A3(new_n392), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n393), .A2(KEYINPUT88), .A3(new_n372), .ZN(new_n394));
  AOI21_X1  g208(.A(KEYINPUT88), .B1(new_n393), .B2(new_n372), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n376), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT20), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT89), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n393), .A2(new_n372), .ZN(new_n399));
  INV_X1    g213(.A(new_n376), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n400), .A2(KEYINPUT20), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n398), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n401), .ZN(new_n403));
  AOI211_X1 g217(.A(KEYINPUT89), .B(new_n403), .C1(new_n393), .C2(new_n372), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n375), .B1(new_n397), .B2(new_n405), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n266), .A2(new_n254), .A3(new_n256), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n269), .A2(new_n268), .ZN(new_n408));
  OAI21_X1  g222(.A(KEYINPUT65), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT65), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n267), .A2(new_n410), .A3(new_n268), .A4(new_n269), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n240), .A2(KEYINPUT10), .A3(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n212), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n261), .A2(new_n262), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n270), .A2(new_n231), .A3(new_n208), .A4(new_n235), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT10), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT11), .ZN(new_n420));
  INV_X1    g234(.A(G134), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n420), .B1(new_n421), .B2(G137), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(G137), .ZN(new_n423));
  INV_X1    g237(.A(G137), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(KEYINPUT11), .A3(G134), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n422), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(G131), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n422), .A2(new_n425), .A3(new_n329), .A4(new_n423), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT77), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n429), .B(new_n430), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n413), .A2(new_n416), .A3(new_n419), .A4(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(G110), .B(G140), .ZN(new_n433));
  INV_X1    g247(.A(G227), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n434), .A2(G953), .ZN(new_n435));
  XOR2_X1   g249(.A(new_n433), .B(new_n435), .Z(new_n436));
  AND2_X1   g250(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n413), .A2(new_n419), .A3(new_n416), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n429), .ZN(new_n439));
  INV_X1    g253(.A(new_n270), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n236), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n417), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n429), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT12), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n442), .A2(KEYINPUT12), .A3(new_n429), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n432), .ZN(new_n448));
  INV_X1    g262(.A(new_n436), .ZN(new_n449));
  AOI22_X1  g263(.A1(new_n437), .A2(new_n439), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(G469), .B1(new_n450), .B2(G902), .ZN(new_n451));
  INV_X1    g265(.A(G469), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT78), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n445), .A2(new_n453), .A3(new_n446), .ZN(new_n454));
  INV_X1    g268(.A(new_n429), .ZN(new_n455));
  AOI211_X1 g269(.A(new_n444), .B(new_n455), .C1(new_n441), .C2(new_n417), .ZN(new_n456));
  AOI21_X1  g270(.A(KEYINPUT12), .B1(new_n442), .B2(new_n429), .ZN(new_n457));
  OAI21_X1  g271(.A(KEYINPUT78), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n454), .A2(new_n458), .A3(new_n432), .A4(new_n436), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n436), .B1(new_n439), .B2(new_n432), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n452), .B(new_n298), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n451), .A2(new_n462), .ZN(new_n463));
  XOR2_X1   g277(.A(KEYINPUT9), .B(G234), .Z(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(G221), .B1(new_n465), .B2(G902), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(KEYINPUT74), .ZN(new_n467));
  INV_X1    g281(.A(G478), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT94), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n469), .A2(KEYINPUT15), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n469), .A2(KEYINPUT15), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n468), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(G128), .B(G143), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n475), .B(new_n421), .ZN(new_n476));
  INV_X1    g290(.A(G122), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(G116), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n213), .A2(G122), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n478), .A2(new_n479), .A3(new_n202), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n213), .A2(KEYINPUT14), .A3(G122), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n478), .A2(new_n479), .ZN(new_n482));
  OAI211_X1 g296(.A(G107), .B(new_n481), .C1(new_n482), .C2(KEYINPUT14), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n476), .A2(new_n480), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT90), .ZN(new_n485));
  AND3_X1   g299(.A1(new_n478), .A2(new_n479), .A3(new_n202), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n202), .B1(new_n478), .B2(new_n479), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n482), .A2(G107), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n489), .A2(KEYINPUT90), .A3(new_n480), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n255), .A2(G128), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n265), .A2(G143), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(new_n493), .A3(new_n421), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT92), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n475), .A2(KEYINPUT92), .A3(new_n421), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(KEYINPUT91), .B(KEYINPUT13), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n475), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n500), .B(G134), .C1(new_n492), .C2(new_n499), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n491), .A2(KEYINPUT93), .A3(new_n498), .A4(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  XOR2_X1   g317(.A(KEYINPUT91), .B(KEYINPUT13), .Z(new_n504));
  INV_X1    g318(.A(new_n492), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n421), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AOI22_X1  g320(.A1(new_n488), .A2(new_n490), .B1(new_n506), .B2(new_n500), .ZN(new_n507));
  AOI21_X1  g321(.A(KEYINPUT93), .B1(new_n507), .B2(new_n498), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n484), .B1(new_n503), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n464), .A2(G217), .A3(new_n190), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NOR3_X1   g325(.A1(new_n486), .A2(new_n487), .A3(new_n485), .ZN(new_n512));
  AOI21_X1  g326(.A(KEYINPUT90), .B1(new_n489), .B2(new_n480), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n498), .B(new_n501), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT93), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n502), .ZN(new_n517));
  INV_X1    g331(.A(new_n510), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n517), .A2(new_n484), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n511), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n474), .B1(new_n520), .B2(new_n298), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n518), .B1(new_n517), .B2(new_n484), .ZN(new_n522));
  INV_X1    g336(.A(new_n484), .ZN(new_n523));
  AOI211_X1 g337(.A(new_n523), .B(new_n510), .C1(new_n516), .C2(new_n502), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n298), .B(new_n474), .C1(new_n522), .C2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n406), .A2(new_n463), .A3(new_n467), .A4(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n187), .B1(new_n324), .B2(new_n528), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n237), .A2(new_n239), .B1(new_n409), .B2(new_n411), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n530), .A2(KEYINPUT10), .B1(new_n415), .B2(new_n414), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n455), .B1(new_n531), .B2(new_n419), .ZN(new_n532));
  INV_X1    g346(.A(new_n432), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n449), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AOI211_X1 g348(.A(G469), .B(G902), .C1(new_n534), .C2(new_n459), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n448), .A2(new_n449), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n439), .A2(new_n432), .A3(new_n436), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n452), .B1(new_n538), .B2(new_n298), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n467), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n375), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT20), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT88), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n366), .A2(KEYINPUT87), .A3(new_n391), .ZN(new_n544));
  AOI21_X1  g358(.A(KEYINPUT87), .B1(new_n366), .B2(new_n391), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n544), .A2(new_n545), .A3(new_n369), .ZN(new_n546));
  INV_X1    g360(.A(new_n372), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n543), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n393), .A2(KEYINPUT88), .A3(new_n372), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n542), .B1(new_n550), .B2(new_n376), .ZN(new_n551));
  INV_X1    g365(.A(new_n402), .ZN(new_n552));
  INV_X1    g366(.A(new_n404), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n527), .B(new_n541), .C1(new_n551), .C2(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n540), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n188), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n312), .B1(new_n299), .B2(new_n310), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n320), .A2(new_n322), .A3(new_n311), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n556), .A2(KEYINPUT95), .A3(new_n560), .A4(new_n198), .ZN(new_n561));
  AOI21_X1  g375(.A(G146), .B1(new_n339), .B2(new_n340), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n265), .A2(G119), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n265), .A2(G119), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT23), .ZN(new_n565));
  OAI211_X1 g379(.A(KEYINPUT69), .B(new_n563), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT69), .ZN(new_n567));
  OAI211_X1 g381(.A(G119), .B(new_n265), .C1(new_n567), .C2(KEYINPUT23), .ZN(new_n568));
  XNOR2_X1  g382(.A(KEYINPUT72), .B(G110), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n564), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n563), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT24), .B(G110), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n562), .B1(new_n570), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n348), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT73), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n575), .A2(KEYINPUT73), .A3(new_n348), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n352), .ZN(new_n581));
  OR2_X1    g395(.A1(new_n572), .A2(new_n573), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n566), .A2(new_n568), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(G110), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT70), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n583), .A2(KEYINPUT70), .A3(G110), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n581), .A2(new_n582), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n580), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(KEYINPUT22), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(G137), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n580), .A2(new_n588), .A3(new_n592), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n298), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(KEYINPUT25), .ZN(new_n597));
  INV_X1    g411(.A(G217), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n598), .B1(G234), .B2(new_n298), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT25), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n594), .A2(new_n600), .A3(new_n595), .A4(new_n298), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n597), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n594), .A2(new_n595), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n599), .A2(G902), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n424), .A2(G134), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n421), .A2(G137), .ZN(new_n609));
  OAI21_X1  g423(.A(G131), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n428), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n269), .A2(new_n268), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n410), .B1(new_n613), .B2(new_n267), .ZN(new_n614));
  INV_X1    g428(.A(new_n411), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n612), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AOI22_X1  g430(.A1(new_n427), .A2(new_n428), .B1(new_n261), .B2(new_n262), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n616), .A2(new_n618), .A3(KEYINPUT30), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT30), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n440), .A2(new_n611), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n620), .B1(new_n621), .B2(new_n617), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n619), .A2(new_n224), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n616), .A2(new_n618), .A3(new_n221), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G101), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n325), .A2(G210), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n623), .A2(new_n624), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(KEYINPUT31), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT31), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n623), .A2(new_n624), .A3(new_n631), .A4(new_n628), .ZN(new_n632));
  AOI21_X1  g446(.A(KEYINPUT66), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT66), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n634), .B1(new_n629), .B2(KEYINPUT31), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n624), .B(KEYINPUT28), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n224), .B1(new_n621), .B2(new_n617), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n628), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n633), .A2(new_n635), .A3(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(G472), .A2(G902), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  OAI21_X1  g455(.A(KEYINPUT32), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n630), .A2(new_n632), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n634), .ZN(new_n644));
  INV_X1    g458(.A(new_n635), .ZN(new_n645));
  INV_X1    g459(.A(new_n638), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT32), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n647), .A2(new_n648), .A3(new_n640), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n642), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n221), .B1(new_n616), .B2(new_n618), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n611), .B1(new_n409), .B2(new_n411), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n652), .A2(new_n224), .A3(new_n617), .ZN(new_n653));
  OAI21_X1  g467(.A(KEYINPUT28), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(KEYINPUT67), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT28), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n624), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT67), .ZN(new_n658));
  OAI211_X1 g472(.A(new_n658), .B(KEYINPUT28), .C1(new_n651), .C2(new_n653), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n655), .A2(KEYINPUT29), .A3(new_n657), .A4(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n628), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n298), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT68), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT29), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n661), .B1(new_n636), .B2(new_n637), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n623), .A2(new_n624), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n667), .A2(new_n628), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n665), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  OAI211_X1 g483(.A(KEYINPUT68), .B(new_n298), .C1(new_n660), .C2(new_n661), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n664), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(G472), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n607), .B1(new_n650), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n529), .A2(new_n561), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G101), .ZN(G3));
  INV_X1    g489(.A(new_n324), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n540), .A2(new_n607), .ZN(new_n677));
  OAI21_X1  g491(.A(G472), .B1(new_n639), .B2(G902), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n647), .A2(new_n640), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n676), .A2(new_n677), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g496(.A(KEYINPUT33), .B1(new_n522), .B2(new_n524), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT33), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n511), .A2(new_n684), .A3(new_n519), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n683), .A2(new_n685), .A3(G478), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n520), .A2(new_n468), .A3(new_n298), .ZN(new_n687));
  NAND2_X1  g501(.A1(G478), .A2(G902), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n400), .B1(new_n548), .B2(new_n549), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n405), .B1(new_n690), .B2(new_n542), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n689), .B1(new_n691), .B2(new_n541), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n682), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT34), .B(G104), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT96), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n694), .B(new_n696), .ZN(G6));
  XOR2_X1   g511(.A(new_n375), .B(KEYINPUT97), .Z(new_n698));
  INV_X1    g512(.A(new_n527), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n690), .A2(new_n542), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n397), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n698), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n682), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT35), .B(G107), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G9));
  OR2_X1    g519(.A1(new_n593), .A2(KEYINPUT36), .ZN(new_n706));
  OR2_X1    g520(.A1(new_n589), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n589), .A2(new_n706), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n707), .A2(new_n605), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(KEYINPUT98), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n602), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n529), .A2(new_n561), .A3(new_n681), .A4(new_n711), .ZN(new_n712));
  XOR2_X1   g526(.A(new_n712), .B(KEYINPUT37), .Z(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G110), .ZN(G12));
  INV_X1    g528(.A(new_n560), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n710), .A2(new_n602), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(G900), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n196), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n191), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n702), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n540), .B1(new_n650), .B2(new_n672), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n717), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G128), .ZN(G30));
  NAND2_X1  g539(.A1(new_n558), .A2(new_n559), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(KEYINPUT99), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT99), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n728), .B1(new_n558), .B2(new_n559), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(KEYINPUT38), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT38), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n732), .B1(new_n727), .B2(new_n729), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n734), .A2(new_n557), .ZN(new_n735));
  INV_X1    g549(.A(G472), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n667), .A2(new_n628), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n651), .A2(new_n653), .ZN(new_n738));
  AOI21_X1  g552(.A(G902), .B1(new_n738), .B2(new_n661), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n736), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n650), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n720), .B(KEYINPUT39), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n463), .A2(new_n467), .A3(new_n743), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n742), .B(new_n716), .C1(new_n744), .C2(KEYINPUT40), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n541), .B1(new_n551), .B2(new_n554), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n699), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n744), .A2(KEYINPUT40), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n735), .A2(new_n746), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G143), .ZN(G45));
  INV_X1    g566(.A(KEYINPUT100), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n753), .B1(new_n692), .B2(new_n720), .ZN(new_n754));
  NOR4_X1   g568(.A1(new_n406), .A2(KEYINPUT100), .A3(new_n689), .A4(new_n721), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(new_n717), .A3(new_n723), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G146), .ZN(G48));
  NOR2_X1   g572(.A1(new_n452), .A2(KEYINPUT101), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n534), .A2(new_n459), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n760), .B1(new_n761), .B2(new_n298), .ZN(new_n762));
  AOI211_X1 g576(.A(G902), .B(new_n759), .C1(new_n534), .C2(new_n459), .ZN(new_n763));
  INV_X1    g577(.A(new_n466), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n673), .A2(new_n676), .A3(new_n692), .A4(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(KEYINPUT41), .B(G113), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n766), .B(new_n767), .ZN(G15));
  INV_X1    g582(.A(new_n702), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n673), .A2(new_n676), .A3(new_n769), .A4(new_n765), .ZN(new_n770));
  XOR2_X1   g584(.A(KEYINPUT102), .B(G116), .Z(new_n771));
  XNOR2_X1  g585(.A(new_n770), .B(new_n771), .ZN(G18));
  AND2_X1   g586(.A1(new_n560), .A2(new_n765), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n197), .B1(new_n650), .B2(new_n672), .ZN(new_n774));
  INV_X1    g588(.A(new_n555), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n773), .A2(new_n774), .A3(new_n775), .A4(new_n711), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G119), .ZN(G21));
  INV_X1    g591(.A(KEYINPUT103), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n607), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n602), .A2(KEYINPUT103), .A3(new_n606), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n655), .A2(new_n659), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n628), .B1(new_n782), .B2(new_n657), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n640), .B1(new_n783), .B2(new_n643), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n678), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n786), .A2(new_n773), .A3(new_n198), .A4(new_n749), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G122), .ZN(G24));
  INV_X1    g602(.A(KEYINPUT104), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n789), .B1(new_n754), .B2(new_n755), .ZN(new_n790));
  INV_X1    g604(.A(new_n689), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n747), .A2(new_n791), .A3(new_n720), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(KEYINPUT100), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n692), .A2(new_n753), .A3(new_n720), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n793), .A2(new_n794), .A3(KEYINPUT104), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n785), .A2(new_n716), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n790), .A2(new_n795), .A3(new_n773), .A4(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G125), .ZN(G27));
  AOI22_X1  g612(.A1(new_n642), .A2(new_n649), .B1(new_n671), .B2(G472), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n764), .B1(new_n451), .B2(new_n462), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n800), .A2(new_n188), .A3(new_n558), .A4(new_n559), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n799), .A2(new_n801), .A3(new_n607), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n802), .A2(new_n790), .A3(new_n795), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT105), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT42), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n802), .A2(new_n790), .A3(KEYINPUT105), .A4(new_n795), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n799), .A2(new_n781), .A3(new_n806), .ZN(new_n809));
  INV_X1    g623(.A(new_n801), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n809), .A2(new_n790), .A3(new_n795), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G131), .ZN(G33));
  NAND2_X1  g627(.A1(new_n802), .A2(new_n722), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G134), .ZN(G36));
  NAND3_X1  g629(.A1(new_n558), .A2(new_n559), .A3(new_n188), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n747), .A2(new_n689), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n817), .A2(KEYINPUT43), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n406), .A2(KEYINPUT43), .A3(new_n791), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n680), .B(new_n711), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT44), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n816), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n818), .A2(new_n819), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n823), .A2(KEYINPUT44), .A3(new_n680), .A4(new_n711), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n450), .A2(KEYINPUT45), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT45), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n538), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n825), .A2(new_n827), .A3(G469), .ZN(new_n828));
  NAND2_X1  g642(.A1(G469), .A2(G902), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT46), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(new_n535), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n828), .A2(KEYINPUT46), .A3(new_n829), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n833), .A2(new_n466), .A3(new_n743), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n822), .A2(new_n824), .A3(new_n834), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(G137), .ZN(G39));
  AOI21_X1  g650(.A(new_n764), .B1(new_n831), .B2(new_n832), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(KEYINPUT47), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n754), .A2(new_n755), .A3(new_n816), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT106), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n799), .A2(new_n607), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n840), .B1(new_n839), .B2(new_n841), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n838), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT107), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n838), .B(KEYINPUT107), .C1(new_n842), .C2(new_n843), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(G140), .ZN(G42));
  INV_X1    g663(.A(KEYINPUT116), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT51), .ZN(new_n851));
  INV_X1    g665(.A(new_n816), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n786), .A2(new_n192), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n818), .A2(new_n819), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n762), .A2(new_n763), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n857), .A2(new_n467), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n852), .B(new_n855), .C1(new_n838), .C2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n852), .A2(new_n192), .A3(new_n765), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n854), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n796), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n188), .B1(new_n731), .B2(new_n733), .ZN(new_n863));
  INV_X1    g677(.A(new_n765), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n853), .A2(new_n854), .A3(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n863), .A2(new_n865), .A3(KEYINPUT50), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT50), .B1(new_n863), .B2(new_n865), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n859), .B(new_n862), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  OR3_X1    g683(.A1(new_n860), .A2(new_n607), .A3(new_n742), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n870), .A2(new_n747), .A3(new_n791), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n851), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n859), .A2(new_n862), .ZN(new_n873));
  INV_X1    g687(.A(new_n871), .ZN(new_n874));
  INV_X1    g688(.A(new_n868), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n866), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n873), .A2(KEYINPUT51), .A3(new_n874), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n855), .A2(new_n773), .ZN(new_n878));
  INV_X1    g692(.A(G952), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n799), .A2(new_n781), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n861), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(KEYINPUT115), .A2(KEYINPUT48), .ZN(new_n882));
  AOI211_X1 g696(.A(new_n879), .B(G953), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n872), .A2(new_n877), .A3(new_n878), .A4(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n870), .A2(new_n693), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT53), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT52), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n800), .A2(new_n720), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n742), .A2(new_n716), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n749), .A2(new_n560), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n891), .A2(KEYINPUT110), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT110), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n740), .B1(new_n642), .B2(new_n649), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n895), .A2(new_n711), .A3(new_n889), .ZN(new_n896));
  INV_X1    g710(.A(new_n892), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n894), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n723), .B(new_n717), .C1(new_n756), .C2(new_n722), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n797), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n888), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(KEYINPUT110), .B1(new_n891), .B2(new_n892), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n896), .A2(new_n897), .A3(new_n894), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n905), .A2(KEYINPUT52), .A3(new_n797), .A4(new_n900), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n902), .A2(KEYINPUT111), .A3(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n901), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT111), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n908), .A2(new_n909), .A3(KEYINPUT52), .A4(new_n905), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n787), .A2(new_n776), .A3(new_n766), .A4(new_n770), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(KEYINPUT108), .B1(new_n747), .B2(new_n527), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT108), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n406), .A2(new_n915), .A3(new_n699), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n914), .A2(new_n693), .A3(new_n916), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n917), .A2(new_n676), .A3(new_n677), .A4(new_n681), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n712), .A2(new_n674), .A3(new_n918), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n913), .A2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT109), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n698), .A2(new_n701), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n723), .A2(new_n922), .A3(new_n711), .A4(new_n852), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n699), .A2(new_n721), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n921), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NOR4_X1   g740(.A1(new_n799), .A2(new_n540), .A3(new_n716), .A4(new_n816), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n927), .A2(KEYINPUT109), .A3(new_n922), .A4(new_n924), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n790), .A2(new_n795), .A3(new_n796), .A4(new_n810), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n930), .A2(new_n814), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n920), .A2(new_n932), .A3(new_n812), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n887), .B1(new_n911), .B2(new_n933), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n808), .A2(new_n811), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n913), .A2(new_n929), .A3(new_n931), .A4(new_n919), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n902), .A2(new_n906), .ZN(new_n938));
  XOR2_X1   g752(.A(KEYINPUT112), .B(KEYINPUT53), .Z(new_n939));
  NAND3_X1  g753(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n934), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(KEYINPUT54), .ZN(new_n942));
  AND4_X1   g756(.A1(KEYINPUT53), .A2(new_n712), .A3(new_n674), .A4(new_n918), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n943), .A2(new_n929), .A3(new_n931), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n808), .B2(new_n811), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n912), .B(KEYINPUT113), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n945), .A2(new_n910), .A3(new_n907), .A4(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n939), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n902), .A2(new_n906), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n948), .B1(new_n933), .B2(new_n949), .ZN(new_n950));
  XOR2_X1   g764(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n947), .A2(new_n950), .A3(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n886), .A2(new_n942), .A3(new_n953), .ZN(new_n954));
  AND2_X1   g768(.A1(KEYINPUT115), .A2(KEYINPUT48), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n881), .A2(new_n882), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n850), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n879), .A2(new_n190), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n947), .A2(new_n950), .A3(new_n952), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT54), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n934), .B2(new_n940), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n956), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n962), .A2(KEYINPUT116), .A3(new_n963), .A4(new_n886), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n957), .A2(new_n958), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n781), .B1(KEYINPUT49), .B2(new_n857), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n966), .B(new_n467), .C1(KEYINPUT49), .C2(new_n857), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n967), .B1(new_n731), .B2(new_n733), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n968), .A2(new_n188), .A3(new_n895), .A4(new_n817), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n965), .A2(new_n969), .ZN(G75));
  INV_X1    g784(.A(G210), .ZN(new_n971));
  AOI211_X1 g785(.A(new_n971), .B(new_n298), .C1(new_n947), .C2(new_n950), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT56), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(KEYINPUT117), .ZN(new_n974));
  OAI21_X1  g788(.A(KEYINPUT55), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n314), .A2(new_n319), .A3(new_n301), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n976), .A2(new_n310), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n947), .A2(new_n950), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n978), .A2(G210), .A3(G902), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT55), .ZN(new_n980));
  INV_X1    g794(.A(new_n974), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  AND3_X1   g796(.A1(new_n975), .A2(new_n977), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n977), .B1(new_n975), .B2(new_n982), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n190), .A2(G952), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n983), .A2(new_n984), .A3(new_n985), .ZN(G51));
  XOR2_X1   g800(.A(new_n829), .B(KEYINPUT57), .Z(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n907), .A2(new_n910), .A3(new_n946), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n932), .A2(new_n812), .A3(new_n943), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n939), .B1(new_n937), .B2(new_n938), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n951), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n988), .B1(new_n993), .B2(new_n953), .ZN(new_n994));
  INV_X1    g808(.A(new_n761), .ZN(new_n995));
  OAI21_X1  g809(.A(KEYINPUT118), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n978), .A2(G902), .ZN(new_n997));
  OR2_X1    g811(.A1(new_n997), .A2(new_n828), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n952), .B1(new_n947), .B2(new_n950), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n987), .B1(new_n959), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT118), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n1000), .A2(new_n1001), .A3(new_n761), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n996), .A2(new_n998), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n879), .A2(G953), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n1003), .A2(new_n1004), .ZN(G54));
  INV_X1    g819(.A(new_n550), .ZN(new_n1006));
  NAND2_X1  g820(.A1(KEYINPUT58), .A2(G475), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1007), .B(KEYINPUT119), .ZN(new_n1008));
  OR3_X1    g822(.A1(new_n997), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1006), .B1(new_n997), .B2(new_n1008), .ZN(new_n1010));
  AND3_X1   g824(.A1(new_n1009), .A2(new_n1004), .A3(new_n1010), .ZN(G60));
  NAND2_X1  g825(.A1(new_n683), .A2(new_n685), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n688), .B(KEYINPUT59), .Z(new_n1013));
  INV_X1    g827(.A(new_n1013), .ZN(new_n1014));
  OAI211_X1 g828(.A(new_n1012), .B(new_n1014), .C1(new_n959), .C2(new_n999), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1013), .B1(new_n942), .B2(new_n953), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n1004), .B(new_n1015), .C1(new_n1016), .C2(new_n1012), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1017), .A2(KEYINPUT120), .ZN(new_n1018));
  OAI211_X1 g832(.A(new_n683), .B(new_n685), .C1(new_n962), .C2(new_n1013), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT120), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n1019), .A2(new_n1020), .A3(new_n1004), .A4(new_n1015), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1018), .A2(new_n1021), .ZN(G63));
  NAND2_X1  g836(.A1(G217), .A2(G902), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n1023), .B(KEYINPUT60), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1024), .B1(new_n947), .B2(new_n950), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n1025), .A2(new_n707), .A3(new_n708), .ZN(new_n1026));
  AND2_X1   g840(.A1(new_n1026), .A2(new_n1004), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n1025), .A2(new_n604), .ZN(new_n1028));
  INV_X1    g842(.A(new_n1028), .ZN(new_n1029));
  INV_X1    g843(.A(KEYINPUT121), .ZN(new_n1030));
  INV_X1    g844(.A(KEYINPUT61), .ZN(new_n1031));
  OAI211_X1 g845(.A(new_n1027), .B(new_n1029), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n1026), .A2(new_n1030), .A3(new_n1004), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1026), .A2(new_n1004), .ZN(new_n1034));
  OAI211_X1 g848(.A(new_n1033), .B(KEYINPUT61), .C1(new_n1034), .C2(new_n1028), .ZN(new_n1035));
  AND2_X1   g849(.A1(new_n1032), .A2(new_n1035), .ZN(G66));
  OAI21_X1  g850(.A(G953), .B1(new_n194), .B2(new_n272), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n1037), .B1(new_n920), .B2(G953), .ZN(new_n1038));
  OAI211_X1 g852(.A(new_n308), .B(new_n309), .C1(G898), .C2(new_n190), .ZN(new_n1039));
  XNOR2_X1  g853(.A(new_n1038), .B(new_n1039), .ZN(G69));
  AOI22_X1  g854(.A1(new_n846), .A2(new_n847), .B1(new_n722), .B2(new_n802), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n835), .A2(new_n908), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n1042), .A2(KEYINPUT123), .ZN(new_n1043));
  INV_X1    g857(.A(KEYINPUT123), .ZN(new_n1044));
  NAND3_X1  g858(.A1(new_n835), .A2(new_n908), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g860(.A1(new_n834), .A2(new_n880), .A3(new_n897), .ZN(new_n1047));
  NAND4_X1  g861(.A1(new_n1041), .A2(new_n1046), .A3(new_n812), .A4(new_n1047), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n1048), .A2(new_n190), .ZN(new_n1049));
  NOR2_X1   g863(.A1(new_n190), .A2(G900), .ZN(new_n1050));
  INV_X1    g864(.A(new_n1050), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g866(.A1(new_n1052), .A2(KEYINPUT124), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n619), .A2(new_n622), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n383), .A2(new_n384), .ZN(new_n1055));
  XOR2_X1   g869(.A(new_n1054), .B(new_n1055), .Z(new_n1056));
  INV_X1    g870(.A(new_n1056), .ZN(new_n1057));
  INV_X1    g871(.A(KEYINPUT124), .ZN(new_n1058));
  NAND3_X1  g872(.A1(new_n1049), .A2(new_n1058), .A3(new_n1051), .ZN(new_n1059));
  NAND3_X1  g873(.A1(new_n1053), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n751), .A2(new_n908), .ZN(new_n1061));
  INV_X1    g875(.A(KEYINPUT62), .ZN(new_n1062));
  NAND2_X1  g876(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g877(.A1(new_n751), .A2(KEYINPUT62), .A3(new_n908), .ZN(new_n1064));
  NAND2_X1  g878(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OR2_X1    g879(.A1(new_n917), .A2(KEYINPUT122), .ZN(new_n1066));
  AOI21_X1  g880(.A(new_n744), .B1(new_n917), .B2(KEYINPUT122), .ZN(new_n1067));
  NAND4_X1  g881(.A1(new_n1066), .A2(new_n1067), .A3(new_n673), .A4(new_n852), .ZN(new_n1068));
  NAND4_X1  g882(.A1(new_n1065), .A2(new_n835), .A3(new_n848), .A4(new_n1068), .ZN(new_n1069));
  NAND2_X1  g883(.A1(new_n1069), .A2(new_n190), .ZN(new_n1070));
  NAND2_X1  g884(.A1(new_n1070), .A2(new_n1056), .ZN(new_n1071));
  OAI21_X1  g885(.A(G953), .B1(new_n434), .B2(new_n718), .ZN(new_n1072));
  INV_X1    g886(.A(new_n1072), .ZN(new_n1073));
  AND3_X1   g887(.A1(new_n1060), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g888(.A(new_n1073), .B1(new_n1060), .B2(new_n1071), .ZN(new_n1075));
  NOR2_X1   g889(.A1(new_n1074), .A2(new_n1075), .ZN(G72));
  NAND2_X1  g890(.A1(G472), .A2(G902), .ZN(new_n1077));
  XOR2_X1   g891(.A(new_n1077), .B(KEYINPUT63), .Z(new_n1078));
  XNOR2_X1  g892(.A(new_n1078), .B(KEYINPUT125), .ZN(new_n1079));
  INV_X1    g893(.A(new_n920), .ZN(new_n1080));
  OAI21_X1  g894(.A(new_n1079), .B1(new_n1048), .B2(new_n1080), .ZN(new_n1081));
  XOR2_X1   g895(.A(new_n1081), .B(KEYINPUT127), .Z(new_n1082));
  INV_X1    g896(.A(new_n668), .ZN(new_n1083));
  NOR2_X1   g897(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g898(.A1(new_n941), .A2(new_n1083), .A3(new_n737), .A4(new_n1078), .ZN(new_n1085));
  OAI21_X1  g899(.A(new_n1079), .B1(new_n1069), .B2(new_n1080), .ZN(new_n1086));
  INV_X1    g900(.A(KEYINPUT126), .ZN(new_n1087));
  NAND2_X1  g901(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  OAI211_X1 g902(.A(KEYINPUT126), .B(new_n1079), .C1(new_n1069), .C2(new_n1080), .ZN(new_n1089));
  NAND2_X1  g903(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g904(.A(new_n1004), .B(new_n1085), .C1(new_n1090), .C2(new_n737), .ZN(new_n1091));
  NOR2_X1   g905(.A1(new_n1084), .A2(new_n1091), .ZN(G57));
endmodule


