//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 1 1 0 0 0 0 0 0 0 0 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 1 0 0 0 1 0 0 1 1 0 1 1 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n764, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n857, new_n858, new_n859, new_n860, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n970, new_n971;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(G134gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G127gat), .ZN(new_n205));
  INV_X1    g004(.A(G127gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G134gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G113gat), .B(G120gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n208), .B1(new_n209), .B2(KEYINPUT1), .ZN(new_n210));
  INV_X1    g009(.A(G120gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G113gat), .ZN(new_n212));
  INV_X1    g011(.A(G113gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G120gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G127gat), .B(G134gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT1), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n210), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G148gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT79), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT79), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G148gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n223), .A3(G141gat), .ZN(new_n224));
  INV_X1    g023(.A(G141gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G148gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(G155gat), .A2(G162gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT2), .ZN(new_n228));
  INV_X1    g027(.A(G155gat), .ZN(new_n229));
  INV_X1    g028(.A(G162gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  AOI22_X1  g030(.A1(new_n224), .A2(new_n226), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n229), .A2(new_n230), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(new_n227), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n220), .A2(G141gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n226), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n234), .B1(new_n228), .B2(new_n236), .ZN(new_n237));
  NOR3_X1   g036(.A1(new_n219), .A2(new_n232), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n224), .A2(new_n226), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n231), .A2(new_n227), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G141gat), .B(G148gat), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n227), .B(new_n233), .C1(new_n242), .C2(KEYINPUT2), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n241), .A2(new_n243), .B1(new_n218), .B2(new_n210), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n203), .B1(new_n238), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT80), .ZN(new_n246));
  OAI21_X1  g045(.A(KEYINPUT3), .B1(new_n232), .B2(new_n237), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n248));
  INV_X1    g047(.A(new_n226), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT79), .B(G148gat), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n249), .B1(new_n250), .B2(G141gat), .ZN(new_n251));
  INV_X1    g050(.A(new_n240), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n243), .B(new_n248), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n247), .A2(new_n253), .A3(new_n219), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT4), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n243), .B1(new_n251), .B2(new_n252), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n255), .B1(new_n256), .B2(new_n219), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n232), .A2(new_n237), .ZN(new_n258));
  AND2_X1   g057(.A1(new_n210), .A2(new_n218), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(new_n259), .A3(KEYINPUT4), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n254), .A2(new_n257), .A3(new_n260), .A4(new_n202), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT80), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n262), .B(new_n203), .C1(new_n238), .C2(new_n244), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n246), .A2(KEYINPUT5), .A3(new_n261), .A4(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT81), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT5), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n267), .B1(new_n245), .B2(KEYINPUT80), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n268), .A2(KEYINPUT81), .A3(new_n261), .A4(new_n263), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n261), .A2(KEYINPUT5), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  XOR2_X1   g072(.A(G1gat), .B(G29gat), .Z(new_n274));
  XNOR2_X1  g073(.A(new_n274), .B(KEYINPUT0), .ZN(new_n275));
  XNOR2_X1  g074(.A(G57gat), .B(G85gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n273), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n271), .B1(new_n266), .B2(new_n269), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT6), .B1(new_n280), .B2(new_n277), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n273), .A2(KEYINPUT6), .A3(new_n278), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AND2_X1   g083(.A1(G226gat), .A2(G233gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n285), .A2(KEYINPUT29), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT25), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT66), .B(G190gat), .ZN(new_n289));
  INV_X1    g088(.A(G183gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT24), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT24), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n294), .A2(G183gat), .A3(G190gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n288), .B1(new_n291), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n298), .A2(KEYINPUT23), .ZN(new_n299));
  AND2_X1   g098(.A1(G169gat), .A2(G176gat), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n300), .B1(KEYINPUT23), .B2(new_n298), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n297), .A2(new_n303), .ZN(new_n304));
  XOR2_X1   g103(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n305));
  INV_X1    g104(.A(G190gat), .ZN(new_n306));
  AOI22_X1  g105(.A1(new_n293), .A2(new_n295), .B1(new_n290), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n305), .B1(new_n302), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(G169gat), .A2(G176gat), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT26), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT68), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT68), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n313), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n300), .B1(new_n311), .B2(new_n310), .ZN(new_n316));
  AOI22_X1  g115(.A1(new_n315), .A2(new_n316), .B1(G183gat), .B2(G190gat), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT27), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G183gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT67), .ZN(new_n320));
  AND2_X1   g119(.A1(new_n289), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n290), .A2(KEYINPUT27), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT67), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT28), .B1(new_n321), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n306), .A2(KEYINPUT66), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT66), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(G190gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n327), .A2(new_n329), .A3(KEYINPUT28), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n330), .A2(new_n323), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n317), .B1(new_n326), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n287), .B1(new_n309), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n307), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n334), .A2(new_n299), .A3(new_n301), .ZN(new_n335));
  AOI22_X1  g134(.A1(new_n335), .A2(new_n305), .B1(new_n297), .B2(new_n303), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT69), .ZN(new_n337));
  XNOR2_X1  g136(.A(KEYINPUT27), .B(G183gat), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n289), .B(new_n320), .C1(new_n338), .C2(KEYINPUT67), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT28), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n331), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n315), .A2(new_n316), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(new_n292), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n337), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  OAI211_X1 g143(.A(KEYINPUT69), .B(new_n317), .C1(new_n326), .C2(new_n331), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n336), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n333), .B1(new_n346), .B2(new_n285), .ZN(new_n347));
  XNOR2_X1  g146(.A(G197gat), .B(G204gat), .ZN(new_n348));
  INV_X1    g147(.A(G218gat), .ZN(new_n349));
  INV_X1    g148(.A(G211gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT73), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT73), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(G211gat), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n349), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n348), .B1(new_n354), .B2(KEYINPUT22), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT74), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT74), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n357), .B(new_n348), .C1(new_n354), .C2(KEYINPUT22), .ZN(new_n358));
  XNOR2_X1  g157(.A(G211gat), .B(G218gat), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n356), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n348), .B(new_n359), .C1(new_n354), .C2(KEYINPUT22), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT75), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n359), .B1(new_n355), .B2(KEYINPUT74), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT75), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n366), .A2(new_n367), .A3(new_n358), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n347), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n309), .A2(new_n332), .A3(new_n285), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n369), .B(new_n371), .C1(new_n346), .C2(new_n287), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G8gat), .B(G36gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(G64gat), .B(G92gat), .ZN(new_n376));
  XOR2_X1   g175(.A(new_n375), .B(new_n376), .Z(new_n377));
  XOR2_X1   g176(.A(new_n377), .B(KEYINPUT76), .Z(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n372), .B(new_n377), .C1(new_n347), .C2(new_n369), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT30), .ZN(new_n381));
  OAI22_X1  g180(.A1(new_n374), .A2(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT77), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI221_X1 g183(.A(KEYINPUT77), .B1(new_n380), .B2(new_n381), .C1(new_n374), .C2(new_n379), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AND3_X1   g185(.A1(new_n380), .A2(KEYINPUT78), .A3(new_n381), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT78), .B1(new_n380), .B2(new_n381), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  AND4_X1   g189(.A1(KEYINPUT82), .A2(new_n284), .A3(new_n386), .A4(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n389), .B1(new_n282), .B2(new_n283), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT82), .B1(new_n392), .B2(new_n386), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n355), .A2(new_n360), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n362), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT29), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n258), .B1(new_n397), .B2(new_n248), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n253), .A2(new_n396), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n398), .B1(new_n369), .B2(new_n399), .ZN(new_n400));
  AND2_X1   g199(.A1(G228gat), .A2(G233gat), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  AND4_X1   g202(.A1(new_n367), .A2(new_n356), .A3(new_n358), .A4(new_n360), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n363), .B1(new_n366), .B2(new_n358), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n399), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n401), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n365), .A2(new_n396), .A3(new_n368), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n258), .B1(new_n408), .B2(new_n248), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT83), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n407), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n404), .A2(new_n405), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT3), .B1(new_n412), .B2(new_n396), .ZN(new_n413));
  OAI21_X1  g212(.A(KEYINPUT83), .B1(new_n413), .B2(new_n258), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n411), .A2(new_n414), .A3(KEYINPUT84), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT84), .B1(new_n411), .B2(new_n414), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n403), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(G22gat), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT84), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n408), .A2(new_n248), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n420), .A2(new_n410), .A3(new_n256), .ZN(new_n421));
  INV_X1    g220(.A(new_n407), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n409), .A2(new_n410), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n419), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n411), .A2(new_n414), .A3(KEYINPUT84), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n402), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(G22gat), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT85), .ZN(new_n430));
  XNOR2_X1  g229(.A(G78gat), .B(G106gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(KEYINPUT31), .B(G50gat), .ZN(new_n432));
  XOR2_X1   g231(.A(new_n431), .B(new_n432), .Z(new_n433));
  NAND4_X1  g232(.A1(new_n418), .A2(new_n429), .A3(new_n430), .A4(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT85), .B1(new_n427), .B2(new_n428), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n436), .A2(new_n433), .B1(new_n418), .B2(new_n429), .ZN(new_n437));
  OAI22_X1  g236(.A1(new_n391), .A2(new_n393), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n344), .A2(new_n345), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n219), .B1(new_n439), .B2(new_n336), .ZN(new_n440));
  NAND2_X1  g239(.A1(G227gat), .A2(G233gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n346), .A2(new_n259), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n441), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT34), .B1(new_n444), .B2(KEYINPUT71), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n440), .A2(new_n441), .A3(new_n442), .A4(new_n445), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g248(.A(G71gat), .B(G99gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n450), .B(KEYINPUT70), .ZN(new_n451));
  INV_X1    g250(.A(G15gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n451), .B(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(G43gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n453), .B(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n346), .A2(new_n259), .ZN(new_n457));
  AOI211_X1 g256(.A(new_n219), .B(new_n336), .C1(new_n344), .C2(new_n345), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n444), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT33), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n456), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n449), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n441), .B1(new_n440), .B2(new_n442), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n455), .B1(new_n463), .B2(KEYINPUT33), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n464), .A2(new_n448), .A3(new_n447), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n459), .A2(KEYINPUT32), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n462), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n467), .B1(new_n462), .B2(new_n465), .ZN(new_n470));
  AND2_X1   g269(.A1(KEYINPUT72), .A2(KEYINPUT36), .ZN(new_n471));
  NOR2_X1   g270(.A1(KEYINPUT72), .A2(KEYINPUT36), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NOR3_X1   g272(.A1(new_n469), .A2(new_n470), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n462), .A2(new_n465), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n466), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n471), .B1(new_n476), .B2(new_n468), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n377), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT37), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n480), .B1(new_n374), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT87), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI211_X1 g283(.A(KEYINPUT87), .B(new_n480), .C1(new_n374), .C2(new_n481), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n372), .B(new_n481), .C1(new_n347), .C2(new_n369), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT38), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n412), .B(new_n371), .C1(new_n346), .C2(new_n287), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n489), .B(KEYINPUT37), .C1(new_n347), .C2(new_n412), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n379), .A2(KEYINPUT38), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n486), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n492), .A2(new_n380), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n282), .A2(new_n283), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n488), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT86), .ZN(new_n496));
  OR2_X1    g295(.A1(new_n238), .A2(new_n244), .ZN(new_n497));
  OAI21_X1  g296(.A(KEYINPUT39), .B1(new_n497), .B2(new_n203), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n254), .A2(new_n257), .A3(new_n260), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n498), .B1(new_n203), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n203), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n277), .B1(new_n501), .B2(KEYINPUT39), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n496), .B1(new_n503), .B2(KEYINPUT40), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT40), .ZN(new_n505));
  OAI211_X1 g304(.A(KEYINPUT86), .B(new_n505), .C1(new_n500), .C2(new_n502), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n503), .A2(KEYINPUT40), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n507), .A2(new_n279), .A3(new_n508), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n389), .A2(new_n382), .ZN(new_n510));
  OR2_X1    g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n430), .B1(new_n417), .B2(G22gat), .ZN(new_n512));
  INV_X1    g311(.A(new_n433), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n427), .A2(new_n428), .ZN(new_n514));
  AOI211_X1 g313(.A(G22gat), .B(new_n402), .C1(new_n425), .C2(new_n426), .ZN(new_n515));
  OAI22_X1  g314(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n495), .A2(new_n511), .A3(new_n516), .A4(new_n434), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n438), .A2(new_n479), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT35), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n469), .A2(new_n470), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n516), .A2(new_n434), .A3(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n391), .A2(new_n393), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n519), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n382), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n284), .A2(new_n524), .A3(new_n390), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT88), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT88), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n392), .A2(new_n527), .A3(new_n524), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n526), .A2(new_n519), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n516), .A2(new_n434), .A3(new_n520), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n518), .B1(new_n523), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(G230gat), .A2(G233gat), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT103), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT7), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(KEYINPUT103), .A2(KEYINPUT7), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n537), .A2(G85gat), .A3(G92gat), .A4(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(G99gat), .ZN(new_n540));
  INV_X1    g339(.A(G106gat), .ZN(new_n541));
  OAI21_X1  g340(.A(KEYINPUT8), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(G85gat), .ZN(new_n543));
  INV_X1    g342(.A(G92gat), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n535), .B(new_n536), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n544), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n539), .A2(new_n542), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(G99gat), .B(G106gat), .Z(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT104), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OR2_X1    g350(.A1(new_n547), .A2(new_n548), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  NOR3_X1   g352(.A1(KEYINPUT100), .A2(G71gat), .A3(G78gat), .ZN(new_n554));
  OAI21_X1  g353(.A(KEYINPUT100), .B1(G71gat), .B2(G78gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(G71gat), .A2(G78gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(G57gat), .B(G64gat), .Z(new_n558));
  AOI211_X1 g357(.A(new_n554), .B(new_n557), .C1(new_n558), .C2(KEYINPUT9), .ZN(new_n559));
  INV_X1    g358(.A(G57gat), .ZN(new_n560));
  OR3_X1    g359(.A1(new_n560), .A2(KEYINPUT101), .A3(G64gat), .ZN(new_n561));
  OAI21_X1  g360(.A(G64gat), .B1(new_n560), .B2(KEYINPUT101), .ZN(new_n562));
  INV_X1    g361(.A(G71gat), .ZN(new_n563));
  INV_X1    g362(.A(G78gat), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT9), .ZN(new_n565));
  AOI22_X1  g364(.A1(new_n561), .A2(new_n562), .B1(new_n556), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n559), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT10), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n567), .A2(new_n552), .A3(new_n549), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  OR3_X1    g371(.A1(new_n553), .A2(new_n570), .A3(new_n568), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT105), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n534), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n576), .B1(new_n575), .B2(new_n574), .ZN(new_n577));
  XOR2_X1   g376(.A(G120gat), .B(G148gat), .Z(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT106), .ZN(new_n579));
  XNOR2_X1  g378(.A(G176gat), .B(G204gat), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n579), .B(new_n580), .Z(new_n581));
  NAND2_X1  g380(.A1(new_n569), .A2(new_n571), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n581), .B1(new_n582), .B2(new_n534), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n577), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n581), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n574), .A2(new_n533), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n582), .A2(new_n534), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OR2_X1    g388(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(KEYINPUT15), .B1(new_n454), .B2(G50gat), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n592), .B1(new_n454), .B2(G50gat), .ZN(new_n593));
  OR3_X1    g392(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(KEYINPUT90), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n594), .A2(KEYINPUT90), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(G29gat), .ZN(new_n600));
  INV_X1    g399(.A(G36gat), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n593), .B1(new_n599), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n593), .A2(new_n602), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n594), .A2(new_n596), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT92), .ZN(new_n606));
  INV_X1    g405(.A(G50gat), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n606), .B1(new_n607), .B2(G43gat), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT91), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n609), .B1(new_n454), .B2(G50gat), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n454), .A2(KEYINPUT92), .A3(G50gat), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n607), .A2(KEYINPUT91), .A3(G43gat), .ZN(new_n612));
  AND4_X1   g411(.A1(new_n608), .A2(new_n610), .A3(new_n611), .A4(new_n612), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n604), .B(new_n605), .C1(KEYINPUT15), .C2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n603), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT17), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n615), .B1(KEYINPUT93), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(KEYINPUT93), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n617), .B(new_n618), .Z(new_n619));
  XNOR2_X1  g418(.A(G15gat), .B(G22gat), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n620), .A2(KEYINPUT94), .ZN(new_n621));
  INV_X1    g420(.A(G1gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(KEYINPUT94), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT96), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n620), .B(KEYINPUT94), .Z(new_n626));
  OAI21_X1  g425(.A(KEYINPUT16), .B1(KEYINPUT95), .B2(G1gat), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n627), .B1(KEYINPUT95), .B2(G1gat), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n624), .B(new_n625), .C1(new_n626), .C2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(G8gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT97), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n619), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n615), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G229gat), .A2(G233gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT98), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n634), .A2(KEYINPUT18), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n630), .B(new_n615), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n636), .B(KEYINPUT13), .Z(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n632), .A2(new_n636), .A3(new_n633), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT18), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n637), .A2(new_n640), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G113gat), .B(G141gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(KEYINPUT89), .B(G197gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g446(.A(KEYINPUT11), .B(G169gat), .Z(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT12), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n644), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n637), .A2(new_n640), .A3(new_n643), .A4(new_n650), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n652), .A2(KEYINPUT99), .A3(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT99), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n644), .A2(new_n655), .A3(new_n651), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n619), .A2(new_n553), .ZN(new_n659));
  NAND2_X1  g458(.A1(G232gat), .A2(G233gat), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(KEYINPUT41), .ZN(new_n662));
  INV_X1    g461(.A(new_n615), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n662), .B1(new_n553), .B2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g465(.A(G190gat), .B(G218gat), .Z(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n661), .A2(KEYINPUT41), .ZN(new_n669));
  XNOR2_X1  g468(.A(G134gat), .B(G162gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n667), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n659), .A2(new_n672), .A3(new_n665), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n668), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n671), .B1(new_n668), .B2(new_n673), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n630), .B1(KEYINPUT21), .B2(new_n567), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n567), .A2(KEYINPUT21), .ZN(new_n678));
  XOR2_X1   g477(.A(G127gat), .B(G155gat), .Z(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n677), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(G231gat), .A2(G233gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT102), .ZN(new_n683));
  XOR2_X1   g482(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(G183gat), .B(G211gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n681), .B(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n676), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n532), .A2(new_n591), .A3(new_n658), .A4(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n690), .A2(new_n284), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(new_n622), .ZN(G1324gat));
  NOR2_X1   g491(.A1(new_n690), .A2(new_n510), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n694), .A2(G8gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(KEYINPUT16), .B(G8gat), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(KEYINPUT42), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n698), .B1(KEYINPUT42), .B2(new_n697), .ZN(G1325gat));
  OAI21_X1  g498(.A(G15gat), .B1(new_n690), .B2(new_n479), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n520), .A2(new_n452), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n700), .B1(new_n690), .B2(new_n701), .ZN(G1326gat));
  NOR2_X1   g501(.A1(new_n435), .A2(new_n437), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n690), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g503(.A(KEYINPUT43), .B(G22gat), .Z(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1327gat));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n392), .A2(new_n386), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT82), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n392), .A2(KEYINPUT82), .A3(new_n386), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT35), .B1(new_n712), .B2(new_n530), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n528), .A2(new_n519), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n521), .A2(new_n526), .A3(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n509), .A2(new_n510), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n716), .B1(new_n488), .B2(new_n494), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n478), .B1(new_n703), .B2(new_n717), .ZN(new_n718));
  AOI22_X1  g517(.A1(new_n713), .A2(new_n715), .B1(new_n718), .B2(new_n438), .ZN(new_n719));
  INV_X1    g518(.A(new_n676), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n707), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n532), .A2(KEYINPUT44), .A3(new_n676), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g522(.A(new_n688), .B(KEYINPUT107), .Z(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n657), .A2(new_n725), .A3(new_n590), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(G29gat), .B1(new_n727), .B2(new_n284), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n591), .A2(new_n688), .A3(new_n676), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n719), .A2(new_n657), .A3(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n284), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n730), .A2(new_n600), .A3(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT45), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n728), .A2(new_n733), .ZN(G1328gat));
  OAI21_X1  g533(.A(G36gat), .B1(new_n727), .B2(new_n510), .ZN(new_n735));
  INV_X1    g534(.A(new_n510), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n730), .A2(new_n601), .A3(new_n736), .ZN(new_n737));
  XOR2_X1   g536(.A(KEYINPUT108), .B(KEYINPUT46), .Z(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n735), .A2(new_n739), .ZN(G1329gat));
  OAI21_X1  g539(.A(G43gat), .B1(new_n727), .B2(new_n479), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT47), .B1(new_n741), .B2(KEYINPUT109), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n730), .A2(new_n454), .A3(new_n520), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n742), .B(new_n744), .ZN(G1330gat));
  OAI21_X1  g544(.A(G50gat), .B1(new_n727), .B2(new_n703), .ZN(new_n746));
  INV_X1    g545(.A(new_n703), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n730), .A2(new_n607), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(KEYINPUT48), .B1(new_n748), .B2(KEYINPUT110), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n749), .B(new_n750), .ZN(G1331gat));
  NAND4_X1  g550(.A1(new_n532), .A2(new_n590), .A3(new_n657), .A4(new_n689), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(new_n284), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(new_n560), .ZN(G1332gat));
  NOR2_X1   g553(.A1(new_n752), .A2(new_n510), .ZN(new_n755));
  NOR2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  AND2_X1   g555(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(new_n755), .B2(new_n756), .ZN(G1333gat));
  OAI21_X1  g558(.A(G71gat), .B1(new_n752), .B2(new_n479), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n520), .A2(new_n563), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n760), .B1(new_n752), .B2(new_n761), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n762), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g562(.A1(new_n752), .A2(new_n703), .ZN(new_n764));
  XNOR2_X1  g563(.A(KEYINPUT111), .B(G78gat), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n764), .B(new_n765), .ZN(G1335gat));
  NAND2_X1  g565(.A1(new_n657), .A2(new_n688), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n767), .A2(new_n591), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n723), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(G85gat), .B1(new_n769), .B2(new_n284), .ZN(new_n770));
  INV_X1    g569(.A(new_n767), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n532), .A2(new_n676), .A3(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n532), .A2(KEYINPUT51), .A3(new_n676), .A4(new_n771), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n590), .A2(new_n543), .A3(new_n731), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(KEYINPUT112), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n770), .B1(new_n777), .B2(new_n779), .ZN(G1336gat));
  INV_X1    g579(.A(KEYINPUT115), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n721), .A2(new_n736), .A3(new_n722), .A4(new_n768), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(G92gat), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n591), .A2(G92gat), .A3(new_n510), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n713), .A2(new_n715), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n720), .B1(new_n785), .B2(new_n518), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT51), .B1(new_n786), .B2(new_n771), .ZN(new_n787));
  INV_X1    g586(.A(new_n775), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n784), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  XOR2_X1   g588(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  AND4_X1   g590(.A1(new_n781), .A2(new_n783), .A3(new_n789), .A4(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n790), .B1(new_n776), .B2(new_n784), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n781), .B1(new_n793), .B2(new_n783), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796));
  AOI22_X1  g595(.A1(new_n789), .A2(KEYINPUT113), .B1(G92gat), .B2(new_n782), .ZN(new_n797));
  INV_X1    g596(.A(new_n784), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n798), .B1(new_n774), .B2(new_n775), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT113), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n796), .B1(new_n797), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(KEYINPUT116), .B1(new_n795), .B2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n801), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n783), .B1(new_n800), .B2(new_n799), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT52), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n806), .B(new_n807), .C1(new_n794), .C2(new_n792), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n803), .A2(new_n808), .ZN(G1337gat));
  OAI21_X1  g608(.A(G99gat), .B1(new_n769), .B2(new_n479), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n776), .A2(new_n540), .A3(new_n520), .A4(new_n590), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XOR2_X1   g611(.A(new_n812), .B(KEYINPUT117), .Z(G1338gat));
  OAI21_X1  g612(.A(G106gat), .B1(new_n769), .B2(new_n703), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n747), .A2(new_n541), .A3(new_n590), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n814), .B1(new_n777), .B2(new_n815), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g616(.A1(new_n657), .A2(new_n591), .A3(new_n689), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n634), .A2(new_n636), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n638), .A2(new_n639), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n649), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n590), .A2(new_n653), .A3(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n574), .A2(new_n823), .A3(new_n533), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n581), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT118), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n824), .A2(KEYINPUT118), .A3(new_n581), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n574), .A2(new_n533), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n829), .A2(new_n823), .ZN(new_n830));
  AOI22_X1  g629(.A1(new_n827), .A2(new_n828), .B1(new_n577), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT55), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n584), .B1(new_n831), .B2(KEYINPUT55), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT119), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n827), .A2(new_n828), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n577), .A2(new_n830), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n839), .A2(new_n840), .A3(new_n584), .A4(new_n832), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n835), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n822), .B1(new_n842), .B2(new_n657), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n676), .A2(new_n653), .A3(new_n821), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n835), .A2(new_n844), .A3(new_n841), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT120), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n835), .A2(new_n844), .A3(KEYINPUT120), .A4(new_n841), .ZN(new_n848));
  AOI22_X1  g647(.A1(new_n720), .A2(new_n843), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n818), .B1(new_n849), .B2(new_n725), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n736), .A2(new_n284), .ZN(new_n851));
  AND3_X1   g650(.A1(new_n850), .A2(new_n521), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n658), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n853), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n590), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(G120gat), .ZN(G1341gat));
  INV_X1    g655(.A(new_n688), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n852), .A2(new_n206), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n852), .A2(new_n725), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n858), .B1(new_n860), .B2(new_n206), .ZN(G1342gat));
  INV_X1    g660(.A(KEYINPUT56), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n852), .B(new_n676), .C1(new_n862), .C2(new_n204), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n204), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n863), .B(new_n864), .ZN(G1343gat));
  NAND2_X1  g664(.A1(new_n479), .A2(new_n851), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n843), .A2(new_n720), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n847), .A2(new_n848), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n725), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n818), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n747), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  XNOR2_X1  g670(.A(KEYINPUT121), .B(KEYINPUT57), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n839), .A2(new_n584), .A3(new_n832), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n822), .B1(new_n657), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n720), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n857), .B1(new_n868), .B2(new_n876), .ZN(new_n877));
  OAI211_X1 g676(.A(KEYINPUT57), .B(new_n747), .C1(new_n877), .C2(new_n870), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n866), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n657), .A2(new_n225), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n703), .A2(new_n478), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n850), .A2(new_n851), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n225), .B1(new_n883), .B2(new_n657), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT58), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n881), .A2(KEYINPUT58), .A3(new_n884), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(G1344gat));
  OAI21_X1  g688(.A(KEYINPUT59), .B1(new_n883), .B2(new_n591), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n250), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n866), .A2(new_n591), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n893), .A2(KEYINPUT59), .ZN(new_n894));
  INV_X1    g693(.A(new_n872), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n895), .B1(new_n850), .B2(new_n747), .ZN(new_n896));
  INV_X1    g695(.A(new_n878), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n894), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n850), .A2(new_n747), .A3(new_n895), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n844), .A2(new_n584), .A3(new_n832), .A4(new_n839), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n876), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n870), .B1(new_n902), .B2(new_n688), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n900), .B1(new_n903), .B2(new_n703), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n893), .B1(new_n899), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n891), .B(new_n898), .C1(new_n905), .C2(new_n906), .ZN(G1345gat));
  NOR3_X1   g706(.A1(new_n883), .A2(KEYINPUT122), .A3(new_n688), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n908), .A2(G155gat), .ZN(new_n909));
  OAI21_X1  g708(.A(KEYINPUT122), .B1(new_n883), .B2(new_n688), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n724), .A2(new_n229), .ZN(new_n911));
  AOI22_X1  g710(.A1(new_n909), .A2(new_n910), .B1(new_n879), .B2(new_n911), .ZN(G1346gat));
  AOI21_X1  g711(.A(new_n230), .B1(new_n879), .B2(new_n676), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n720), .A2(G162gat), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n850), .A2(new_n851), .A3(new_n882), .A4(new_n914), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT123), .ZN(new_n916));
  OAI21_X1  g715(.A(KEYINPUT124), .B1(new_n913), .B2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(new_n866), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n918), .B1(new_n896), .B2(new_n897), .ZN(new_n919));
  OAI21_X1  g718(.A(G162gat), .B1(new_n919), .B2(new_n720), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT123), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n915), .B(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT124), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n920), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n917), .A2(new_n924), .ZN(G1347gat));
  NOR3_X1   g724(.A1(new_n530), .A2(new_n731), .A3(new_n510), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n850), .A2(new_n658), .A3(new_n926), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(G169gat), .ZN(G1348gat));
  NAND3_X1  g727(.A1(new_n850), .A2(new_n590), .A3(new_n926), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g729(.A1(new_n850), .A2(new_n926), .ZN(new_n931));
  OAI21_X1  g730(.A(G183gat), .B1(new_n931), .B2(new_n724), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n857), .A2(new_n338), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g734(.A1(new_n850), .A2(new_n676), .A3(new_n926), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n937), .A2(KEYINPUT125), .A3(new_n306), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT125), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n939), .B1(new_n936), .B2(G190gat), .ZN(new_n940));
  XNOR2_X1  g739(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n941));
  OR3_X1    g740(.A1(new_n938), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NOR2_X1   g741(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n943), .B1(new_n938), .B2(new_n940), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n937), .A2(new_n289), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n942), .A2(new_n944), .A3(new_n945), .ZN(G1351gat));
  AND2_X1   g745(.A1(new_n850), .A2(new_n882), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n731), .A2(new_n510), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(G197gat), .B1(new_n950), .B2(new_n658), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n479), .A2(new_n948), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n952), .B1(new_n899), .B2(new_n904), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n658), .A2(G197gat), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n951), .B1(new_n953), .B2(new_n954), .ZN(G1352gat));
  OR2_X1    g754(.A1(new_n591), .A2(G204gat), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n949), .A2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT62), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n957), .B1(KEYINPUT127), .B2(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(new_n953), .ZN(new_n960));
  OAI21_X1  g759(.A(G204gat), .B1(new_n960), .B2(new_n591), .ZN(new_n961));
  XNOR2_X1  g760(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n962));
  OAI211_X1 g761(.A(new_n959), .B(new_n961), .C1(new_n957), .C2(new_n962), .ZN(G1353gat));
  NAND4_X1  g762(.A1(new_n950), .A2(new_n351), .A3(new_n353), .A4(new_n857), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n953), .A2(new_n857), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT63), .B1(new_n965), .B2(G211gat), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT63), .ZN(new_n967));
  AOI211_X1 g766(.A(new_n967), .B(new_n350), .C1(new_n953), .C2(new_n857), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n964), .B1(new_n966), .B2(new_n968), .ZN(G1354gat));
  OAI21_X1  g768(.A(G218gat), .B1(new_n960), .B2(new_n720), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n950), .A2(new_n349), .A3(new_n676), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(G1355gat));
endmodule


