//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 1 1 0 1 0 0 1 0 1 0 1 1 0 0 0 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1308, new_n1309,
    new_n1310, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1381, new_n1382, new_n1383;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI211_X1 g0005(.A(G50), .B(G77), .C1(new_n203), .C2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n209));
  INV_X1    g0009(.A(G238), .ZN(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  OAI221_X1 g0012(.A(new_n209), .B1(new_n202), .B2(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n214));
  INV_X1    g0014(.A(G77), .ZN(new_n215));
  INV_X1    g0015(.A(G244), .ZN(new_n216));
  INV_X1    g0016(.A(G107), .ZN(new_n217));
  INV_X1    g0017(.A(G264), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n208), .B1(new_n213), .B2(new_n219), .ZN(new_n220));
  OR2_X1    g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n208), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G257), .ZN(new_n224));
  AOI211_X1 g0024(.A(new_n212), .B(new_n223), .C1(new_n224), .C2(new_n218), .ZN(new_n225));
  OR2_X1    g0025(.A1(new_n225), .A2(KEYINPUT0), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n203), .A2(new_n205), .ZN(new_n227));
  INV_X1    g0027(.A(G50), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n229), .A2(G20), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n225), .A2(KEYINPUT0), .ZN(new_n233));
  NAND4_X1  g0033(.A1(new_n221), .A2(new_n226), .A3(new_n232), .A4(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n220), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(KEYINPUT65), .Z(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  INV_X1    g0037(.A(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G358));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n246), .B(new_n247), .Z(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XOR2_X1   g0049(.A(G107), .B(G116), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT66), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT66), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G33), .A3(G41), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n254), .A2(new_n256), .A3(new_n231), .ZN(new_n257));
  INV_X1    g0057(.A(G1), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n258), .B1(G41), .B2(G45), .ZN(new_n259));
  INV_X1    g0059(.A(G274), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n257), .A2(G232), .A3(new_n259), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G223), .A2(G1698), .ZN(new_n264));
  INV_X1    g0064(.A(G226), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n264), .B1(new_n265), .B2(G1698), .ZN(new_n266));
  OR2_X1    g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n266), .A2(new_n269), .B1(G33), .B2(G87), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n230), .B1(G33), .B2(G41), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  OAI211_X1 g0072(.A(new_n262), .B(new_n263), .C1(new_n270), .C2(new_n272), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n273), .A2(G169), .ZN(new_n274));
  INV_X1    g0074(.A(G179), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G20), .ZN(new_n278));
  INV_X1    g0078(.A(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G159), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G58), .A2(G68), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n203), .A2(new_n205), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n282), .B1(new_n284), .B2(G20), .ZN(new_n285));
  AND2_X1   g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NOR2_X1   g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  NOR3_X1   g0087(.A1(new_n286), .A2(new_n287), .A3(G20), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT7), .ZN(new_n289));
  OAI21_X1  g0089(.A(G68), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n267), .A2(new_n278), .A3(new_n268), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(KEYINPUT76), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT76), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT7), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g0096(.A(KEYINPUT16), .B(new_n285), .C1(new_n290), .C2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT77), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n202), .B1(new_n291), .B2(KEYINPUT7), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n299), .B1(new_n291), .B2(new_n295), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT77), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n300), .A2(new_n301), .A3(KEYINPUT16), .A4(new_n285), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT68), .ZN(new_n305));
  AND3_X1   g0105(.A1(new_n304), .A2(new_n305), .A3(new_n230), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n305), .B1(new_n304), .B2(new_n230), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n267), .A2(KEYINPUT7), .A3(new_n278), .A4(new_n268), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n309), .B1(new_n288), .B2(new_n295), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G68), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n285), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT16), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n303), .A2(new_n308), .A3(new_n314), .ZN(new_n315));
  XNOR2_X1  g0115(.A(KEYINPUT8), .B(G58), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT69), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n201), .A2(KEYINPUT69), .A3(KEYINPUT8), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n320), .B1(new_n258), .B2(G20), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n258), .A2(G13), .A3(G20), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n308), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n320), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n325), .B1(new_n326), .B2(new_n322), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n277), .B1(new_n315), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT18), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n304), .A2(new_n230), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT68), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n304), .A2(new_n305), .A3(new_n230), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n335), .B1(new_n298), .B2(new_n302), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n327), .B1(new_n336), .B2(new_n314), .ZN(new_n337));
  OAI21_X1  g0137(.A(KEYINPUT18), .B1(new_n337), .B2(new_n277), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n331), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G200), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n273), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(G190), .B2(new_n273), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n315), .A2(new_n342), .A3(new_n328), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT17), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n337), .A2(KEYINPUT17), .A3(new_n342), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n339), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(G20), .A2(G33), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n349), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n278), .A2(G33), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n350), .B1(new_n215), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n308), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT75), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n353), .A2(new_n354), .ZN(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT11), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n357), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT11), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n359), .A2(new_n360), .A3(new_n355), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n202), .B1(new_n258), .B2(G20), .ZN(new_n362));
  OAI21_X1  g0162(.A(KEYINPUT12), .B1(new_n322), .B2(G68), .ZN(new_n363));
  OR3_X1    g0163(.A1(new_n322), .A2(KEYINPUT12), .A3(G68), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n324), .A2(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n358), .A2(new_n361), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT14), .ZN(new_n367));
  XOR2_X1   g0167(.A(KEYINPUT74), .B(KEYINPUT13), .Z(new_n368));
  INV_X1    g0168(.A(new_n259), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n230), .B1(KEYINPUT66), .B2(new_n253), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n369), .B1(new_n370), .B2(new_n256), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n371), .A2(G238), .B1(new_n257), .B2(new_n261), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n238), .A2(G1698), .ZN(new_n373));
  OAI221_X1 g0173(.A(new_n373), .B1(G226), .B2(G1698), .C1(new_n286), .C2(new_n287), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G33), .A2(G97), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n374), .A2(KEYINPUT73), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n271), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT73), .B1(new_n374), .B2(new_n375), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n368), .B(new_n372), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n374), .A2(new_n375), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT73), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n383), .A2(new_n271), .A3(new_n376), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n368), .B1(new_n384), .B2(new_n372), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n367), .B(G169), .C1(new_n380), .C2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n372), .B1(new_n377), .B2(new_n378), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT13), .ZN(new_n389));
  OAI211_X1 g0189(.A(G179), .B(new_n379), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n368), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n387), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n379), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n367), .B1(new_n394), .B2(G169), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n366), .B1(new_n391), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n366), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n394), .A2(G200), .ZN(new_n398));
  OAI211_X1 g0198(.A(G190), .B(new_n379), .C1(new_n388), .C2(new_n389), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n269), .A2(G1698), .ZN(new_n401));
  OAI22_X1  g0201(.A1(new_n401), .A2(new_n210), .B1(new_n217), .B2(new_n269), .ZN(new_n402));
  INV_X1    g0202(.A(G1698), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n269), .A2(G232), .A3(new_n403), .ZN(new_n404));
  OR2_X1    g0204(.A1(new_n404), .A2(KEYINPUT70), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(KEYINPUT70), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n402), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n407), .A2(new_n272), .ZN(new_n408));
  INV_X1    g0208(.A(new_n371), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n262), .B1(new_n409), .B2(new_n216), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(G169), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G20), .A2(G77), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n211), .A2(KEYINPUT15), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT15), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(G87), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  OAI221_X1 g0220(.A(new_n415), .B1(new_n316), .B2(new_n280), .C1(new_n420), .C2(new_n351), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n421), .A2(new_n308), .B1(new_n215), .B2(new_n323), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n324), .B(G77), .C1(G1), .C2(new_n278), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n411), .A2(new_n275), .ZN(new_n425));
  AND3_X1   g0225(.A1(new_n414), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n412), .A2(G200), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n424), .B1(new_n411), .B2(G190), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AND4_X1   g0229(.A1(new_n348), .A2(new_n396), .A3(new_n400), .A4(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n262), .B1(new_n409), .B2(new_n265), .ZN(new_n431));
  INV_X1    g0231(.A(G223), .ZN(new_n432));
  OAI22_X1  g0232(.A1(new_n401), .A2(new_n432), .B1(new_n215), .B2(new_n269), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n269), .A2(G222), .A3(new_n403), .ZN(new_n434));
  OR2_X1    g0234(.A1(new_n434), .A2(KEYINPUT67), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(KEYINPUT67), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n433), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n431), .B1(new_n438), .B2(new_n271), .ZN(new_n439));
  OR2_X1    g0239(.A1(new_n439), .A2(G169), .ZN(new_n440));
  INV_X1    g0240(.A(G150), .ZN(new_n441));
  OAI22_X1  g0241(.A1(new_n320), .A2(new_n351), .B1(new_n441), .B2(new_n280), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n278), .B1(new_n227), .B2(new_n228), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n308), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n228), .B1(new_n258), .B2(G20), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n324), .A2(new_n445), .B1(new_n228), .B2(new_n323), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n439), .A2(new_n275), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n440), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  XNOR2_X1  g0249(.A(new_n447), .B(KEYINPUT71), .ZN(new_n450));
  OAI21_X1  g0250(.A(KEYINPUT72), .B1(new_n450), .B2(KEYINPUT9), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT71), .ZN(new_n452));
  XNOR2_X1  g0252(.A(new_n447), .B(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT72), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT9), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n451), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n439), .A2(G190), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n458), .B1(new_n340), .B2(new_n439), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n459), .B1(KEYINPUT9), .B2(new_n450), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT10), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT10), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n457), .A2(new_n463), .A3(new_n460), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n449), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n430), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT84), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n258), .A2(G33), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n335), .A2(new_n322), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n419), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT83), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT19), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n278), .B1(new_n375), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(G97), .A2(G107), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n211), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n278), .B(G68), .C1(new_n286), .C2(new_n287), .ZN(new_n478));
  INV_X1    g0278(.A(G97), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n473), .B1(new_n351), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n477), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n308), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n419), .A2(new_n322), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n472), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  AOI211_X1 g0285(.A(KEYINPUT83), .B(new_n483), .C1(new_n481), .C2(new_n308), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n471), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OR2_X1    g0287(.A1(KEYINPUT82), .A2(G116), .ZN(new_n488));
  NAND2_X1  g0288(.A1(KEYINPUT82), .A2(G116), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G33), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n210), .A2(new_n403), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n216), .A2(G1698), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n492), .B(new_n493), .C1(new_n286), .C2(new_n287), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n271), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n258), .A2(G45), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n212), .ZN(new_n498));
  INV_X1    g0298(.A(G45), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n499), .A2(G1), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n260), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n257), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n496), .A2(new_n275), .A3(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n502), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n272), .B1(new_n491), .B2(new_n494), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n413), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n487), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n470), .A2(G87), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n485), .B2(new_n486), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n496), .A2(G190), .A3(new_n502), .ZN(new_n511));
  OAI21_X1  g0311(.A(G200), .B1(new_n504), .B2(new_n505), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n467), .B1(new_n508), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n482), .A2(new_n484), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT83), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n482), .A2(new_n472), .A3(new_n484), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AND2_X1   g0319(.A1(new_n511), .A2(new_n512), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n519), .A2(new_n520), .A3(new_n509), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n487), .A2(new_n507), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT84), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n515), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n217), .A2(KEYINPUT6), .A3(G97), .ZN(new_n525));
  XOR2_X1   g0325(.A(G97), .B(G107), .Z(new_n526));
  OAI21_X1  g0326(.A(new_n525), .B1(new_n526), .B2(KEYINPUT6), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n527), .A2(G20), .B1(G77), .B2(new_n349), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n310), .A2(G107), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n335), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n322), .A2(G97), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(new_n469), .B2(new_n479), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n403), .A2(G244), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(new_n267), .B2(new_n268), .ZN(new_n536));
  OR2_X1    g0336(.A1(KEYINPUT78), .A2(KEYINPUT4), .ZN(new_n537));
  AOI21_X1  g0337(.A(KEYINPUT79), .B1(G33), .B2(G283), .ZN(new_n538));
  NAND3_X1  g0338(.A1(KEYINPUT79), .A2(G33), .A3(G283), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  OAI22_X1  g0340(.A1(new_n536), .A2(new_n537), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n216), .A2(G1698), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n542), .B(new_n537), .C1(new_n287), .C2(new_n286), .ZN(new_n543));
  OAI211_X1 g0343(.A(G250), .B(G1698), .C1(new_n286), .C2(new_n287), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n271), .B1(new_n541), .B2(new_n545), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n254), .A2(new_n256), .A3(new_n231), .ZN(new_n547));
  NOR2_X1   g0347(.A1(KEYINPUT5), .A2(G41), .ZN(new_n548));
  AND2_X1   g0348(.A1(KEYINPUT5), .A2(G41), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n500), .B(G274), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(KEYINPUT80), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n548), .ZN(new_n552));
  NAND2_X1  g0352(.A1(KEYINPUT5), .A2(G41), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n497), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT80), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n554), .A2(new_n257), .A3(new_n555), .A4(G274), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n547), .A2(new_n554), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(G257), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n546), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(G169), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n551), .A2(new_n556), .B1(new_n558), .B2(G257), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n562), .A2(G179), .A3(new_n546), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n534), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  OR2_X1    g0364(.A1(new_n530), .A2(new_n533), .ZN(new_n565));
  INV_X1    g0365(.A(new_n560), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n565), .B1(G190), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT81), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(new_n566), .B2(new_n340), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n560), .A2(KEYINPUT81), .A3(G200), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n564), .B1(new_n567), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT20), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n488), .A2(G20), .A3(new_n489), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n332), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n278), .B1(new_n479), .B2(G33), .ZN(new_n576));
  INV_X1    g0376(.A(new_n538), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n576), .B1(new_n577), .B2(new_n539), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n573), .B1(new_n575), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(G20), .B1(new_n279), .B2(G97), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(new_n540), .B2(new_n538), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n581), .A2(KEYINPUT20), .A3(new_n332), .A4(new_n574), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n335), .A2(G116), .A3(new_n322), .A4(new_n468), .ZN(new_n584));
  INV_X1    g0384(.A(new_n490), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n323), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(G303), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n267), .A2(new_n588), .A3(new_n268), .ZN(new_n589));
  NOR2_X1   g0389(.A1(G257), .A2(G1698), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n590), .B1(new_n218), .B2(G1698), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n286), .A2(new_n287), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n271), .B(new_n589), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n500), .B1(new_n549), .B2(new_n548), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n257), .A2(new_n594), .A3(G270), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n557), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n587), .A2(G169), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(KEYINPUT21), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT21), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n587), .A2(new_n600), .A3(G169), .A4(new_n597), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n596), .A2(new_n557), .A3(G179), .ZN(new_n604));
  OAI21_X1  g0404(.A(KEYINPUT85), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n604), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT85), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n606), .A2(new_n607), .A3(new_n587), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(G250), .A2(G1698), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n610), .B1(new_n224), .B2(G1698), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n269), .ZN(new_n612));
  NAND2_X1  g0412(.A1(G33), .A2(G294), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n272), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n257), .A2(new_n594), .A3(G264), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n617), .A2(new_n275), .A3(new_n557), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n557), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n413), .ZN(new_n620));
  AND2_X1   g0420(.A1(KEYINPUT82), .A2(G116), .ZN(new_n621));
  NOR2_X1   g0421(.A1(KEYINPUT82), .A2(G116), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n278), .B(G33), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  OR2_X1    g0423(.A1(new_n623), .A2(KEYINPUT86), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT23), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n625), .B1(new_n278), .B2(G107), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n217), .A2(KEYINPUT23), .A3(G20), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n623), .A2(KEYINPUT86), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n278), .B(G87), .C1(new_n286), .C2(new_n287), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT22), .ZN(new_n631));
  XNOR2_X1  g0431(.A(new_n630), .B(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(KEYINPUT24), .B1(new_n629), .B2(new_n632), .ZN(new_n633));
  XNOR2_X1  g0433(.A(new_n630), .B(KEYINPUT22), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT24), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n634), .A2(new_n635), .A3(new_n624), .A4(new_n628), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n335), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n322), .A2(G107), .ZN(new_n638));
  XNOR2_X1  g0438(.A(new_n638), .B(KEYINPUT25), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(new_n469), .B2(new_n217), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n618), .B(new_n620), .C1(new_n637), .C2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n602), .A2(new_n609), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(G190), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n617), .A2(new_n643), .A3(new_n557), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(KEYINPUT87), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT87), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n617), .A2(new_n557), .A3(new_n646), .A4(new_n643), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n619), .A2(new_n340), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n645), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n633), .A2(new_n636), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n640), .B1(new_n650), .B2(new_n308), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n587), .B1(G200), .B2(new_n597), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n653), .B1(new_n643), .B2(new_n597), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n642), .A2(new_n655), .ZN(new_n656));
  AND4_X1   g0456(.A1(new_n466), .A2(new_n524), .A3(new_n572), .A4(new_n656), .ZN(G372));
  INV_X1    g0457(.A(KEYINPUT89), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT26), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n659), .B1(new_n524), .B2(new_n564), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n561), .A2(new_n563), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n534), .B1(new_n661), .B2(KEYINPUT88), .ZN(new_n662));
  INV_X1    g0462(.A(new_n510), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n663), .A2(new_n520), .B1(new_n487), .B2(new_n507), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT88), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n561), .A2(new_n665), .A3(new_n563), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n662), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n522), .B1(new_n667), .B2(KEYINPUT26), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n658), .B1(new_n660), .B2(new_n668), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT84), .ZN(new_n670));
  AOI21_X1  g0470(.A(KEYINPUT84), .B1(new_n521), .B2(new_n522), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n564), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(KEYINPUT26), .ZN(new_n673));
  AND4_X1   g0473(.A1(G179), .A2(new_n546), .A3(new_n557), .A4(new_n559), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n413), .B1(new_n562), .B2(new_n546), .ZN(new_n675));
  OAI21_X1  g0475(.A(KEYINPUT88), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n676), .A2(new_n666), .A3(new_n565), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n521), .A2(new_n522), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n508), .B1(new_n679), .B2(new_n659), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n673), .A2(new_n680), .A3(KEYINPUT89), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n678), .B1(new_n651), .B2(new_n649), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n682), .A2(new_n572), .A3(new_n642), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n669), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n466), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n449), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n462), .A2(new_n464), .ZN(new_n687));
  INV_X1    g0487(.A(new_n400), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n347), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n414), .A2(new_n424), .A3(new_n425), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n396), .A2(new_n690), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n687), .B1(new_n339), .B2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n685), .A2(new_n686), .A3(new_n693), .ZN(G369));
  NAND2_X1  g0494(.A1(new_n602), .A2(new_n609), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n258), .A2(new_n278), .A3(G13), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G213), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(G343), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n603), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n695), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n654), .ZN(new_n705));
  INV_X1    g0505(.A(G330), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n701), .B1(new_n637), .B2(new_n640), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n652), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n641), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n641), .A2(new_n701), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n707), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n701), .B1(new_n602), .B2(new_n609), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n712), .B1(new_n710), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n714), .A2(new_n716), .ZN(G399));
  NOR2_X1   g0517(.A1(new_n223), .A2(G41), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n476), .A2(G116), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n719), .A2(G1), .A3(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n229), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n721), .B1(new_n722), .B2(new_n719), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT28), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT91), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n725), .B1(new_n684), .B2(new_n702), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n726), .A2(KEYINPUT29), .ZN(new_n727));
  AOI21_X1  g0527(.A(KEYINPUT91), .B1(new_n684), .B2(new_n702), .ZN(new_n728));
  OAI21_X1  g0528(.A(KEYINPUT92), .B1(new_n667), .B2(new_n659), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n729), .B1(new_n659), .B2(new_n672), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT92), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n679), .A2(new_n731), .A3(KEYINPUT26), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n683), .A2(new_n732), .A3(new_n522), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n702), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(KEYINPUT29), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n728), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n656), .A2(new_n524), .A3(new_n572), .A4(new_n702), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT31), .ZN(new_n738));
  AOI21_X1  g0538(.A(G179), .B1(new_n496), .B2(new_n502), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n619), .A2(new_n560), .A3(new_n597), .A4(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n492), .A2(new_n493), .ZN(new_n742));
  AOI22_X1  g0542(.A1(new_n742), .A2(new_n269), .B1(new_n490), .B2(G33), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n502), .B1(new_n743), .B2(new_n272), .ZN(new_n744));
  AOI22_X1  g0544(.A1(new_n611), .A2(new_n269), .B1(G33), .B2(G294), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n615), .B1(new_n745), .B2(new_n272), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n593), .A2(new_n595), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n748), .B1(new_n556), .B2(new_n551), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n747), .A2(new_n749), .A3(G179), .ZN(new_n750));
  OAI21_X1  g0550(.A(KEYINPUT30), .B1(new_n750), .B2(new_n560), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT30), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n566), .A2(new_n606), .A3(new_n752), .A4(new_n747), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n741), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT90), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n701), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AOI211_X1 g0556(.A(KEYINPUT90), .B(new_n741), .C1(new_n751), .C2(new_n753), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n738), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n751), .A2(new_n753), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n740), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n760), .A2(KEYINPUT31), .A3(new_n701), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n737), .A2(new_n758), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G330), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n727), .A2(new_n736), .A3(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n724), .B1(new_n765), .B2(G1), .ZN(G364));
  AND2_X1   g0566(.A1(new_n278), .A2(G13), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n258), .B1(new_n767), .B2(G45), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n718), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n707), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(G330), .B1(new_n704), .B2(new_n654), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G13), .A2(G33), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(G20), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n705), .A2(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n231), .B1(new_n278), .B2(G169), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n778), .A2(KEYINPUT93), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(KEYINPUT93), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n278), .A2(G179), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G190), .A2(G200), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G159), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n783), .A2(new_n643), .A3(G200), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n787), .A2(KEYINPUT32), .B1(G107), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(G20), .A2(G179), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G200), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n643), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n275), .A2(new_n340), .A3(G190), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G20), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n790), .B1(new_n228), .B2(new_n795), .C1(new_n479), .C2(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n783), .A2(G190), .A3(G200), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n211), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n793), .A2(G190), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n802), .B1(new_n787), .B2(KEYINPUT32), .C1(new_n202), .C2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n792), .A2(new_n784), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n791), .A2(new_n643), .A3(G200), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n269), .B1(new_n806), .B2(new_n215), .C1(new_n808), .C2(new_n201), .ZN(new_n809));
  OR3_X1    g0609(.A1(new_n799), .A2(new_n805), .A3(new_n809), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n786), .A2(G329), .B1(new_n807), .B2(G322), .ZN(new_n811));
  INV_X1    g0611(.A(new_n806), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n269), .B1(new_n812), .B2(G311), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n794), .A2(G326), .ZN(new_n815));
  XNOR2_X1  g0615(.A(KEYINPUT33), .B(G317), .ZN(new_n816));
  INV_X1    g0616(.A(new_n800), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n803), .A2(new_n816), .B1(new_n817), .B2(G303), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n789), .A2(G283), .B1(new_n797), .B2(G294), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n814), .A2(new_n815), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n782), .B1(new_n810), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n781), .A2(new_n776), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n822), .B(KEYINPUT94), .Z(new_n823));
  NAND2_X1  g0623(.A1(new_n269), .A2(new_n222), .ZN(new_n824));
  INV_X1    g0624(.A(G355), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n824), .A2(new_n825), .B1(G116), .B2(new_n222), .ZN(new_n826));
  OR2_X1    g0626(.A1(new_n248), .A2(new_n499), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n223), .A2(new_n269), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(new_n229), .B2(new_n499), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n826), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n770), .B1(new_n823), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n821), .A2(new_n832), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n771), .A2(new_n773), .B1(new_n777), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(G396));
  NOR2_X1   g0635(.A1(new_n781), .A2(new_n774), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n770), .B1(new_n837), .B2(G77), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n414), .A2(new_n424), .A3(new_n425), .A4(new_n702), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n427), .A2(new_n428), .B1(new_n424), .B2(new_n701), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n839), .B1(new_n426), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n842), .A2(new_n775), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n803), .A2(G283), .B1(new_n812), .B2(new_n490), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT95), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n798), .A2(new_n479), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n211), .A2(new_n788), .B1(new_n800), .B2(new_n217), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n846), .B(new_n847), .C1(G303), .C2(new_n794), .ZN(new_n848));
  INV_X1    g0648(.A(G294), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n592), .B1(new_n808), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(G311), .B2(new_n786), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n845), .A2(new_n848), .A3(new_n851), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n812), .A2(G159), .B1(G143), .B2(new_n807), .ZN(new_n853));
  INV_X1    g0653(.A(G137), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n853), .B1(new_n804), .B2(new_n441), .C1(new_n854), .C2(new_n795), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT34), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(G132), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n269), .B1(new_n785), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(G58), .B2(new_n797), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n817), .A2(G50), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n789), .A2(G68), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n857), .A2(new_n860), .A3(new_n861), .A4(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n855), .A2(new_n856), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n852), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n838), .B(new_n843), .C1(new_n781), .C2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n429), .A2(new_n702), .ZN(new_n867));
  INV_X1    g0667(.A(new_n683), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n673), .A2(new_n680), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n868), .B1(new_n869), .B2(new_n658), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n867), .B1(new_n870), .B2(new_n681), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n701), .B1(new_n870), .B2(new_n681), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n872), .B1(new_n873), .B2(new_n842), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n874), .A2(new_n763), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n874), .A2(new_n763), .ZN(new_n876));
  AOI211_X1 g0676(.A(new_n770), .B(new_n875), .C1(KEYINPUT96), .C2(new_n876), .ZN(new_n877));
  OR2_X1    g0677(.A1(new_n876), .A2(KEYINPUT96), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n866), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(G384));
  INV_X1    g0680(.A(G116), .ZN(new_n881));
  NOR3_X1   g0681(.A1(new_n230), .A2(new_n278), .A3(new_n881), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n527), .B(KEYINPUT97), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT35), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n886), .B1(new_n885), .B2(new_n884), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n887), .B(KEYINPUT36), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n229), .A2(G77), .A3(new_n283), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n228), .A2(G68), .ZN(new_n890));
  AOI211_X1 g0690(.A(new_n258), .B(G13), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n315), .A2(new_n342), .A3(new_n328), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n893), .A2(new_n329), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT37), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n699), .B(KEYINPUT99), .ZN(new_n896));
  AOI221_X4 g0696(.A(new_n335), .B1(new_n312), .B2(new_n313), .C1(new_n298), .C2(new_n302), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n896), .B1(new_n897), .B2(new_n327), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n894), .A2(new_n895), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n285), .B1(new_n290), .B2(new_n296), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT16), .B1(new_n900), .B2(KEYINPUT98), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(KEYINPUT98), .B2(new_n900), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n327), .B1(new_n902), .B2(new_n336), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n343), .B1(new_n903), .B2(new_n699), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n903), .A2(new_n277), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT37), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n899), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n903), .A2(new_n699), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n339), .B2(new_n347), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n907), .A2(new_n909), .A3(KEYINPUT38), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT102), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT101), .ZN(new_n912));
  AND4_X1   g0712(.A1(KEYINPUT17), .A2(new_n315), .A3(new_n342), .A4(new_n328), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT17), .B1(new_n337), .B2(new_n342), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n315), .A2(new_n328), .ZN(new_n916));
  INV_X1    g0716(.A(new_n277), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n330), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI211_X1 g0718(.A(KEYINPUT18), .B(new_n277), .C1(new_n315), .C2(new_n328), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n345), .A2(KEYINPUT101), .A3(new_n346), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n915), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n896), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(new_n315), .B2(new_n328), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT100), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n337), .B2(new_n923), .ZN(new_n927));
  AOI22_X1  g0727(.A1(new_n894), .A2(new_n898), .B1(KEYINPUT37), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n916), .A2(new_n917), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n929), .A2(new_n898), .A3(new_n343), .ZN(new_n930));
  OAI21_X1  g0730(.A(KEYINPUT37), .B1(new_n924), .B2(KEYINPUT100), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n925), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT38), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n911), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AOI211_X1 g0736(.A(KEYINPUT102), .B(KEYINPUT38), .C1(new_n925), .C2(new_n933), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n910), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n395), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n939), .A2(new_n390), .A3(new_n386), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n366), .B(new_n701), .C1(new_n940), .C2(new_n688), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n366), .A2(new_n701), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n396), .A2(new_n400), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n841), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n760), .A2(KEYINPUT90), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n754), .A2(new_n755), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n945), .A2(KEYINPUT31), .A3(new_n701), .A4(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n737), .A2(new_n947), .A3(new_n758), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n944), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(KEYINPUT104), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT104), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n944), .A2(new_n948), .A3(new_n951), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n952), .A2(KEYINPUT40), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n938), .A2(new_n950), .A3(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT40), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n907), .A2(new_n909), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n935), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n957), .A2(new_n910), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n955), .B1(new_n958), .B2(new_n949), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n954), .A2(new_n959), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT105), .Z(new_n961));
  NAND2_X1  g0761(.A1(new_n466), .A2(new_n948), .ZN(new_n962));
  OAI21_X1  g0762(.A(G330), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(new_n962), .B2(new_n961), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n940), .A2(new_n366), .A3(new_n702), .ZN(new_n965));
  INV_X1    g0765(.A(new_n910), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n966), .A2(KEYINPUT39), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n936), .B2(new_n937), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n957), .A2(new_n910), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(KEYINPUT39), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n965), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n941), .A2(new_n943), .ZN(new_n972));
  INV_X1    g0772(.A(new_n839), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n969), .B(new_n972), .C1(new_n871), .C2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n920), .A2(new_n896), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(KEYINPUT103), .B1(new_n971), .B2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n867), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n973), .B1(new_n684), .B2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n972), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n975), .B1(new_n982), .B2(new_n969), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT103), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n894), .A2(KEYINPUT100), .A3(KEYINPUT37), .A4(new_n898), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n930), .A2(new_n931), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(new_n924), .B2(new_n922), .ZN(new_n988));
  OAI21_X1  g0788(.A(KEYINPUT102), .B1(new_n988), .B2(KEYINPUT38), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n934), .A2(new_n911), .A3(new_n935), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n991), .A2(new_n967), .B1(KEYINPUT39), .B2(new_n969), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n983), .B(new_n984), .C1(new_n992), .C2(new_n965), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n978), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n693), .A2(new_n686), .ZN(new_n995));
  OAI22_X1  g0795(.A1(KEYINPUT29), .A2(new_n726), .B1(new_n728), .B2(new_n735), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n995), .B1(new_n996), .B2(new_n466), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n994), .B(new_n997), .Z(new_n998));
  OAI22_X1  g0798(.A1(new_n964), .A2(new_n998), .B1(new_n258), .B2(new_n767), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n964), .A2(new_n998), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n892), .B1(new_n999), .B2(new_n1000), .ZN(G367));
  OAI21_X1  g0801(.A(new_n822), .B1(new_n222), .B2(new_n420), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n244), .A2(new_n829), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n770), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT108), .Z(new_n1005));
  NOR2_X1   g0805(.A1(new_n663), .A2(new_n702), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n508), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n678), .B2(new_n1006), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n776), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n817), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1010));
  INV_X1    g0810(.A(G311), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1010), .B1(new_n217), .B2(new_n798), .C1(new_n1011), .C2(new_n795), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n269), .B1(new_n786), .B2(G317), .ZN(new_n1013));
  INV_X1    g0813(.A(G283), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1013), .B1(new_n1014), .B2(new_n806), .C1(new_n588), .C2(new_n808), .ZN(new_n1015));
  AOI21_X1  g0815(.A(KEYINPUT46), .B1(new_n817), .B2(new_n490), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n804), .A2(new_n849), .B1(new_n788), .B2(new_n479), .ZN(new_n1017));
  NOR4_X1   g0817(.A1(new_n1012), .A2(new_n1015), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n803), .A2(G159), .B1(new_n812), .B2(G50), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT109), .Z(new_n1020));
  INV_X1    g0820(.A(G143), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n795), .A2(new_n1021), .B1(new_n202), .B2(new_n798), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n269), .B1(new_n785), .B2(new_n854), .C1(new_n808), .C2(new_n441), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n201), .A2(new_n800), .B1(new_n788), .B2(new_n215), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1018), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1026), .A2(KEYINPUT47), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(KEYINPUT47), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n781), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1005), .B1(new_n1008), .B2(new_n1009), .C1(new_n1027), .C2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT45), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n716), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n565), .A2(new_n701), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n572), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n662), .A2(new_n666), .A3(new_n701), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1031), .B1(new_n1032), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n716), .A2(new_n1036), .A3(KEYINPUT45), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1032), .A2(new_n1037), .A3(KEYINPUT44), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT44), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n716), .B2(new_n1036), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1040), .A2(new_n714), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT107), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1040), .A2(new_n1044), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n714), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1047), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1048), .A2(new_n1046), .A3(new_n1049), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n713), .B(new_n715), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(new_n707), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n765), .B1(new_n1053), .B2(new_n1056), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n718), .B(KEYINPUT41), .Z(new_n1058));
  INV_X1    g0858(.A(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n769), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1008), .A2(KEYINPUT43), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1036), .B(KEYINPUT106), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n641), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n564), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n701), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n713), .A2(new_n715), .A3(new_n1036), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT42), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1061), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1008), .A2(KEYINPUT43), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1070), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1072), .B(new_n1061), .C1(new_n1066), .C2(new_n1068), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1062), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1075), .A2(new_n714), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1074), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1071), .A2(new_n1076), .A3(new_n1073), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1030), .B1(new_n1060), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT110), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  OAI211_X1 g0883(.A(KEYINPUT110), .B(new_n1030), .C1(new_n1060), .C2(new_n1080), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1083), .A2(new_n1084), .ZN(G387));
  NAND2_X1  g0885(.A1(new_n764), .A2(new_n1056), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1055), .A2(new_n727), .A3(new_n736), .A4(new_n763), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1086), .A2(new_n718), .A3(new_n1087), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n824), .A2(new_n720), .B1(G107), .B2(new_n222), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n829), .B1(new_n241), .B2(G45), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n316), .A2(G50), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT50), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n499), .B1(new_n202), .B2(new_n215), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n720), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1093), .B1(new_n1094), .B2(KEYINPUT111), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1092), .B(new_n1095), .C1(KEYINPUT111), .C2(new_n1094), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1089), .B1(new_n1090), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n770), .B1(new_n1097), .B2(new_n823), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n808), .A2(new_n228), .B1(new_n806), .B2(new_n202), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n592), .B(new_n1099), .C1(G150), .C2(new_n786), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(G159), .A2(new_n794), .B1(new_n789), .B2(G97), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n800), .A2(new_n215), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n419), .B2(new_n797), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n326), .A2(new_n803), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1100), .A2(new_n1101), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n269), .B1(new_n786), .B2(G326), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n798), .A2(new_n1014), .B1(new_n800), .B2(new_n849), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n812), .A2(G303), .B1(G317), .B2(new_n807), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(KEYINPUT112), .B(G322), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n1108), .B1(new_n804), .B2(new_n1011), .C1(new_n795), .C2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT48), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1107), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n1111), .B2(new_n1110), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT49), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n1106), .B1(new_n585), .B2(new_n788), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  AND2_X1   g0915(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1105), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1098), .B1(new_n1117), .B2(new_n781), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n713), .B2(new_n1009), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT113), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n1055), .B2(new_n769), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1088), .A2(new_n1121), .ZN(G393));
  NOR2_X1   g0922(.A1(new_n1053), .A2(new_n1087), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1123), .A2(new_n719), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1050), .A2(new_n1045), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1087), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n822), .B1(new_n479), .B2(new_n222), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(new_n251), .B2(new_n828), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n770), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n794), .A2(G150), .B1(G159), .B2(new_n807), .ZN(new_n1132));
  XOR2_X1   g0932(.A(new_n1132), .B(KEYINPUT51), .Z(new_n1133));
  OAI22_X1  g0933(.A1(new_n804), .A2(new_n228), .B1(new_n788), .B2(new_n211), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n269), .B1(new_n785), .B2(new_n1021), .C1(new_n316), .C2(new_n806), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n798), .A2(new_n215), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n800), .A2(new_n202), .ZN(new_n1137));
  NOR4_X1   g0937(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .A4(new_n1137), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n794), .A2(G317), .B1(G311), .B2(new_n807), .ZN(new_n1139));
  XOR2_X1   g0939(.A(new_n1139), .B(KEYINPUT52), .Z(new_n1140));
  OAI22_X1  g0940(.A1(new_n804), .A2(new_n588), .B1(new_n585), .B2(new_n798), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n592), .B1(new_n806), .B2(new_n849), .C1(new_n785), .C2(new_n1109), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n217), .A2(new_n788), .B1(new_n800), .B2(new_n1014), .ZN(new_n1143));
  NOR3_X1   g0943(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1133), .A2(new_n1138), .B1(new_n1140), .B2(new_n1144), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n1131), .B1(new_n782), .B2(new_n1145), .C1(new_n1062), .C2(new_n1009), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n1125), .B2(new_n768), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1127), .A2(new_n1148), .ZN(G390));
  OAI21_X1  g0949(.A(new_n965), .B1(new_n980), .B2(new_n981), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1150), .A2(new_n968), .A3(new_n970), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n965), .B(KEYINPUT114), .ZN(new_n1152));
  OR2_X1    g0952(.A1(new_n426), .A2(new_n840), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n702), .B(new_n1153), .C1(new_n730), .C2(new_n733), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(new_n839), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT115), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n396), .A2(new_n400), .A3(new_n942), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n942), .B1(new_n396), .B2(new_n400), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1156), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n941), .A2(KEYINPUT115), .A3(new_n943), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1152), .B1(new_n1155), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n938), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n841), .A2(new_n706), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n762), .A2(new_n972), .A3(new_n1165), .ZN(new_n1166));
  AND3_X1   g0966(.A1(new_n1151), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n948), .A2(new_n1165), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1168), .A2(new_n981), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(new_n1151), .B2(new_n1164), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1167), .A2(new_n1171), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1166), .A2(new_n1154), .A3(new_n839), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n1168), .A2(new_n1161), .A3(KEYINPUT117), .ZN(new_n1174));
  AOI21_X1  g0974(.A(KEYINPUT117), .B1(new_n1168), .B2(new_n1161), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1173), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n972), .B1(new_n762), .B2(new_n1165), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n1169), .A2(new_n1177), .B1(new_n871), .B2(new_n973), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n430), .A2(new_n465), .A3(G330), .A4(new_n948), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1180), .B(KEYINPUT116), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n997), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1172), .A2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1182), .B1(new_n1167), .B2(new_n1171), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1184), .A2(new_n1185), .A3(new_n718), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n804), .A2(new_n217), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1136), .B(new_n1187), .C1(G283), .C2(new_n794), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n785), .A2(new_n849), .B1(new_n806), .B2(new_n479), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n269), .B(new_n1189), .C1(G116), .C2(new_n807), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1188), .A2(new_n1190), .A3(new_n802), .A4(new_n862), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT54), .B(G143), .ZN(new_n1192));
  INV_X1    g0992(.A(G125), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n806), .A2(new_n1192), .B1(new_n785), .B2(new_n1193), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n592), .B(new_n1194), .C1(G132), .C2(new_n807), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n800), .A2(new_n441), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1196), .B(new_n1197), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(G128), .A2(new_n794), .B1(new_n789), .B2(G50), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n803), .A2(G137), .B1(G159), .B2(new_n797), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1195), .A2(new_n1198), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n782), .B1(new_n1191), .B2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1130), .B1(new_n836), .B2(new_n320), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT118), .Z(new_n1204));
  AOI211_X1 g1004(.A(new_n1202), .B(new_n1204), .C1(new_n992), .C2(new_n774), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(new_n1172), .B2(new_n769), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1186), .A2(new_n1206), .ZN(G378));
  INV_X1    g1007(.A(KEYINPUT122), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n687), .A2(new_n686), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n450), .A2(new_n699), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1210), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n465), .A2(new_n1212), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1211), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1214), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n465), .A2(new_n1212), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n449), .B(new_n1210), .C1(new_n462), .C2(new_n464), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1216), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1215), .A2(new_n1219), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n954), .A2(new_n1220), .A3(G330), .A4(new_n959), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n966), .B1(new_n989), .B2(new_n990), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n950), .A2(KEYINPUT40), .A3(new_n952), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n959), .B(G330), .C1(new_n1222), .C2(new_n1223), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n1215), .A2(new_n1219), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  AND4_X1   g1026(.A1(new_n993), .A2(new_n978), .A3(new_n1221), .A4(new_n1226), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n993), .A2(new_n978), .B1(new_n1226), .B2(new_n1221), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1208), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n997), .A2(new_n1181), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1184), .A2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1226), .A2(new_n1221), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n994), .A2(new_n1233), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n978), .A2(new_n993), .A3(new_n1226), .A4(new_n1221), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1234), .A2(KEYINPUT122), .A3(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1229), .A2(new_n1232), .A3(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT57), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1238), .B1(new_n1184), .B2(new_n1231), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n719), .B1(new_n1240), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1239), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1229), .A2(new_n769), .A3(new_n1236), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1225), .A2(new_n774), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n770), .B1(new_n837), .B2(G50), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n804), .A2(new_n479), .B1(new_n788), .B2(new_n201), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n269), .A2(G41), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n1249), .B1(new_n1014), .B2(new_n785), .C1(new_n420), .C2(new_n806), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n1102), .B(new_n1250), .C1(G68), .C2(new_n797), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n807), .A2(G107), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n1252), .B(KEYINPUT121), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1251), .A2(new_n1253), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n1248), .B(new_n1254), .C1(G116), .C2(new_n794), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(KEYINPUT58), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1249), .A2(new_n1257), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(KEYINPUT120), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1256), .A2(new_n1259), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n812), .A2(G137), .B1(G128), .B2(new_n807), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1261), .B1(new_n800), .B2(new_n1192), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n1193), .A2(new_n795), .B1(new_n804), .B2(new_n858), .ZN(new_n1263));
  AOI211_X1 g1063(.A(new_n1262), .B(new_n1263), .C1(G150), .C2(new_n797), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1265), .A2(KEYINPUT59), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(KEYINPUT59), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n789), .A2(G159), .ZN(new_n1268));
  AOI211_X1 g1068(.A(G33), .B(G41), .C1(new_n786), .C2(G124), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1267), .A2(new_n1268), .A3(new_n1269), .ZN(new_n1270));
  OAI221_X1 g1070(.A(new_n1260), .B1(KEYINPUT58), .B2(new_n1255), .C1(new_n1266), .C2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1247), .B1(new_n1271), .B2(new_n781), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1246), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1245), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1244), .A2(new_n1275), .ZN(G375));
  NAND2_X1  g1076(.A1(new_n1179), .A2(new_n769), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1130), .B1(new_n836), .B2(new_n202), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n794), .A2(G132), .ZN(new_n1279));
  OAI221_X1 g1079(.A(new_n1279), .B1(new_n854), .B2(new_n808), .C1(new_n804), .C2(new_n1192), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1280), .A2(KEYINPUT124), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n592), .B1(new_n786), .B2(G128), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1282), .B1(new_n441), .B2(new_n806), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n798), .A2(new_n228), .ZN(new_n1284));
  OAI22_X1  g1084(.A1(new_n201), .A2(new_n788), .B1(new_n800), .B2(new_n281), .ZN(new_n1285));
  NOR4_X1   g1085(.A1(new_n1281), .A2(new_n1283), .A3(new_n1284), .A4(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1280), .A2(KEYINPUT124), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n592), .B1(new_n788), .B2(new_n215), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(new_n1288), .B(KEYINPUT123), .ZN(new_n1289));
  AOI22_X1  g1089(.A1(G303), .A2(new_n786), .B1(new_n812), .B2(G107), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1290), .B1(new_n1014), .B2(new_n808), .ZN(new_n1291));
  OAI22_X1  g1091(.A1(new_n804), .A2(new_n585), .B1(new_n420), .B2(new_n798), .ZN(new_n1292));
  OAI22_X1  g1092(.A1(new_n795), .A2(new_n849), .B1(new_n800), .B2(new_n479), .ZN(new_n1293));
  NOR3_X1   g1093(.A1(new_n1291), .A2(new_n1292), .A3(new_n1293), .ZN(new_n1294));
  AOI22_X1  g1094(.A1(new_n1286), .A2(new_n1287), .B1(new_n1289), .B2(new_n1294), .ZN(new_n1295));
  OAI221_X1 g1095(.A(new_n1278), .B1(new_n782), .B2(new_n1295), .C1(new_n1162), .C2(new_n775), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1277), .A2(new_n1296), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1183), .A2(new_n1058), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1179), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1230), .A2(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1297), .B1(new_n1298), .B2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(G381));
  NAND3_X1  g1102(.A1(new_n1088), .A2(new_n834), .A3(new_n1121), .ZN(new_n1303));
  NOR3_X1   g1103(.A1(G390), .A2(G384), .A3(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(G378), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1304), .A2(new_n1305), .A3(new_n1301), .ZN(new_n1306));
  OR3_X1    g1106(.A1(G375), .A2(G387), .A3(new_n1306), .ZN(G407));
  NAND2_X1  g1107(.A1(new_n700), .A2(G213), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1305), .A2(new_n1309), .ZN(new_n1310));
  OAI211_X1 g1110(.A(G407), .B(G213), .C1(G375), .C2(new_n1310), .ZN(G409));
  XNOR2_X1  g1111(.A(new_n1081), .B(G390), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT125), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1303), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n834), .B1(new_n1088), .B2(new_n1121), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1313), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(G393), .A2(G396), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1317), .A2(KEYINPUT125), .A3(new_n1303), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1316), .A2(new_n1318), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1312), .A2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT126), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1147), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1083), .A2(new_n1084), .A3(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n768), .ZN(new_n1325));
  AND2_X1   g1125(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1327), .A2(G390), .A3(new_n1030), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1319), .A2(new_n1328), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1321), .B1(new_n1323), .B2(new_n1329), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1083), .A2(new_n1084), .A3(new_n1322), .ZN(new_n1331));
  NAND4_X1  g1131(.A1(new_n1331), .A2(KEYINPUT126), .A3(new_n1319), .A4(new_n1328), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1320), .B1(new_n1330), .B2(new_n1332), .ZN(new_n1333));
  NOR3_X1   g1133(.A1(new_n1167), .A2(new_n1182), .A3(new_n1171), .ZN(new_n1334));
  OAI21_X1  g1134(.A(KEYINPUT57), .B1(new_n1334), .B2(new_n1230), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n718), .B1(new_n1335), .B2(new_n1241), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1336), .B1(new_n1238), .B2(new_n1237), .ZN(new_n1337));
  NOR3_X1   g1137(.A1(new_n1337), .A2(new_n1305), .A3(new_n1274), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1242), .A2(new_n769), .ZN(new_n1339));
  OAI211_X1 g1139(.A(new_n1273), .B(new_n1339), .C1(new_n1237), .C2(new_n1058), .ZN(new_n1340));
  AND2_X1   g1140(.A1(new_n1340), .A2(new_n1305), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1308), .B1(new_n1338), .B2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT60), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1300), .B1(new_n1183), .B2(new_n1343), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1230), .A2(KEYINPUT60), .A3(new_n1299), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1344), .A2(new_n718), .A3(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1297), .ZN(new_n1347));
  AND3_X1   g1147(.A1(new_n1346), .A2(G384), .A3(new_n1347), .ZN(new_n1348));
  AOI21_X1  g1148(.A(G384), .B1(new_n1346), .B2(new_n1347), .ZN(new_n1349));
  NOR2_X1   g1149(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1309), .A2(G2897), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1352));
  OAI211_X1 g1152(.A(G2897), .B(new_n1309), .C1(new_n1348), .C2(new_n1349), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1352), .A2(new_n1353), .ZN(new_n1354));
  INV_X1    g1154(.A(new_n1354), .ZN(new_n1355));
  AOI21_X1  g1155(.A(KEYINPUT61), .B1(new_n1342), .B2(new_n1355), .ZN(new_n1356));
  OAI211_X1 g1156(.A(new_n1308), .B(new_n1350), .C1(new_n1338), .C2(new_n1341), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1357), .A2(KEYINPUT62), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1356), .A2(new_n1358), .ZN(new_n1359));
  NOR2_X1   g1159(.A1(new_n1357), .A2(KEYINPUT62), .ZN(new_n1360));
  OAI21_X1  g1160(.A(new_n1333), .B1(new_n1359), .B2(new_n1360), .ZN(new_n1361));
  INV_X1    g1161(.A(KEYINPUT127), .ZN(new_n1362));
  INV_X1    g1162(.A(KEYINPUT63), .ZN(new_n1363));
  NOR3_X1   g1163(.A1(new_n1348), .A2(new_n1349), .A3(new_n1363), .ZN(new_n1364));
  OAI211_X1 g1164(.A(new_n1308), .B(new_n1364), .C1(new_n1338), .C2(new_n1341), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1330), .A2(new_n1332), .ZN(new_n1366));
  INV_X1    g1166(.A(new_n1320), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1366), .A2(new_n1367), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1365), .A2(new_n1368), .ZN(new_n1369));
  INV_X1    g1169(.A(KEYINPUT61), .ZN(new_n1370));
  NAND3_X1  g1170(.A1(new_n1244), .A2(G378), .A3(new_n1275), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1340), .A2(new_n1305), .ZN(new_n1372));
  AOI21_X1  g1172(.A(new_n1309), .B1(new_n1371), .B2(new_n1372), .ZN(new_n1373));
  OAI21_X1  g1173(.A(new_n1370), .B1(new_n1373), .B2(new_n1354), .ZN(new_n1374));
  NOR2_X1   g1174(.A1(new_n1369), .A2(new_n1374), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1357), .A2(new_n1363), .ZN(new_n1376));
  AOI21_X1  g1176(.A(new_n1362), .B1(new_n1375), .B2(new_n1376), .ZN(new_n1377));
  AOI21_X1  g1177(.A(new_n1333), .B1(new_n1373), .B2(new_n1364), .ZN(new_n1378));
  AND4_X1   g1178(.A1(new_n1362), .A2(new_n1356), .A3(new_n1378), .A4(new_n1376), .ZN(new_n1379));
  OAI21_X1  g1179(.A(new_n1361), .B1(new_n1377), .B2(new_n1379), .ZN(G405));
  AOI21_X1  g1180(.A(G378), .B1(new_n1244), .B2(new_n1275), .ZN(new_n1381));
  NOR2_X1   g1181(.A1(new_n1338), .A2(new_n1381), .ZN(new_n1382));
  XNOR2_X1  g1182(.A(new_n1382), .B(new_n1350), .ZN(new_n1383));
  XNOR2_X1  g1183(.A(new_n1383), .B(new_n1368), .ZN(G402));
endmodule


