//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n548, new_n549, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n563, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n594, new_n595,
    new_n598, new_n600, new_n601, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1184,
    new_n1185, new_n1186, new_n1187;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT65), .B(G2066), .ZN(G411));
  XNOR2_X1  g006(.A(KEYINPUT66), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  OAI21_X1  g035(.A(G125), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n458), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI211_X1 g038(.A(G137), .B(new_n458), .C1(new_n459), .C2(new_n460), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n463), .A2(new_n468), .ZN(G160));
  OR2_X1    g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(G2105), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G136), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n458), .B1(new_n470), .B2(new_n471), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  OR2_X1    g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n458), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n473), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G162));
  OAI211_X1 g054(.A(G126), .B(G2105), .C1(new_n459), .C2(new_n460), .ZN(new_n480));
  OR2_X1    g055(.A1(G102), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G114), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n481), .A2(new_n483), .A3(G2104), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n480), .A2(KEYINPUT67), .A3(new_n484), .ZN(new_n488));
  OAI211_X1 g063(.A(G138), .B(new_n458), .C1(new_n459), .C2(new_n460), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  XNOR2_X1  g065(.A(KEYINPUT3), .B(G2104), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n491), .A2(new_n492), .A3(G138), .A4(new_n458), .ZN(new_n493));
  AOI22_X1  g068(.A1(new_n487), .A2(new_n488), .B1(new_n490), .B2(new_n493), .ZN(G164));
  INV_X1    g069(.A(KEYINPUT6), .ZN(new_n495));
  OAI21_X1  g070(.A(KEYINPUT68), .B1(new_n495), .B2(G651), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n497));
  INV_X1    g072(.A(G651), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n497), .A2(new_n498), .A3(KEYINPUT6), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n495), .A2(G651), .ZN(new_n501));
  AND3_X1   g076(.A1(new_n500), .A2(G543), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G50), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n504));
  AND2_X1   g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  OAI21_X1  g081(.A(G62), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n504), .B1(new_n509), .B2(G651), .ZN(new_n510));
  AOI211_X1 g085(.A(KEYINPUT70), .B(new_n498), .C1(new_n507), .C2(new_n508), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n503), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT5), .B(G543), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n500), .A2(new_n501), .A3(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT69), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g091(.A1(new_n500), .A2(KEYINPUT69), .A3(new_n501), .A4(new_n513), .ZN(new_n517));
  AND3_X1   g092(.A1(new_n516), .A2(G88), .A3(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n512), .A2(new_n518), .ZN(G166));
  AND2_X1   g094(.A1(new_n516), .A2(new_n517), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G89), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n502), .A2(G51), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n525));
  AND2_X1   g100(.A1(G63), .A2(G651), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n524), .A2(new_n525), .B1(new_n513), .B2(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n521), .A2(new_n528), .ZN(G168));
  NAND2_X1  g104(.A1(new_n520), .A2(G90), .ZN(new_n530));
  NAND2_X1  g105(.A1(G77), .A2(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n505), .A2(new_n506), .ZN(new_n532));
  INV_X1    g107(.A(G64), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n502), .A2(G52), .B1(G651), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n530), .A2(new_n535), .ZN(G301));
  INV_X1    g111(.A(G301), .ZN(G171));
  NAND2_X1  g112(.A1(G68), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G56), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n532), .B2(new_n539), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n502), .A2(G43), .B1(G651), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n516), .A2(new_n517), .ZN(new_n542));
  INV_X1    g117(.A(G81), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(G188));
  NAND2_X1  g125(.A1(new_n502), .A2(G53), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT71), .ZN(new_n552));
  AOI21_X1  g127(.A(KEYINPUT72), .B1(new_n552), .B2(KEYINPUT9), .ZN(new_n553));
  NAND2_X1  g128(.A1(G78), .A2(G543), .ZN(new_n554));
  XOR2_X1   g129(.A(KEYINPUT73), .B(G65), .Z(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n555), .B2(new_n532), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n551), .A2(new_n553), .B1(G651), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n516), .A2(G91), .A3(new_n517), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n553), .B1(KEYINPUT72), .B2(KEYINPUT9), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n502), .A2(G53), .A3(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n557), .A2(new_n558), .A3(new_n560), .ZN(G299));
  INV_X1    g136(.A(G168), .ZN(G286));
  INV_X1    g137(.A(G88), .ZN(new_n563));
  OAI221_X1 g138(.A(new_n503), .B1(new_n510), .B2(new_n511), .C1(new_n542), .C2(new_n563), .ZN(G303));
  OR2_X1    g139(.A1(new_n513), .A2(G74), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n502), .A2(G49), .B1(new_n565), .B2(G651), .ZN(new_n566));
  INV_X1    g141(.A(G87), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n542), .B2(new_n567), .ZN(G288));
  NAND3_X1  g143(.A1(new_n516), .A2(G86), .A3(new_n517), .ZN(new_n569));
  NAND2_X1  g144(.A1(G73), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G61), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n532), .B2(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n502), .A2(G48), .B1(G651), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n569), .A2(new_n573), .ZN(G305));
  AOI22_X1  g149(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n575), .A2(new_n498), .ZN(new_n576));
  XOR2_X1   g151(.A(new_n576), .B(KEYINPUT74), .Z(new_n577));
  AOI21_X1  g152(.A(new_n577), .B1(G47), .B2(new_n502), .ZN(new_n578));
  INV_X1    g153(.A(G85), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n579), .B2(new_n542), .ZN(G290));
  NAND2_X1  g155(.A1(G301), .A2(G868), .ZN(new_n581));
  NAND2_X1  g156(.A1(G79), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G66), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n532), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n502), .A2(G54), .B1(G651), .B2(new_n584), .ZN(new_n585));
  XOR2_X1   g160(.A(new_n585), .B(KEYINPUT75), .Z(new_n586));
  INV_X1    g161(.A(G92), .ZN(new_n587));
  OAI21_X1  g162(.A(KEYINPUT10), .B1(new_n542), .B2(new_n587), .ZN(new_n588));
  OR3_X1    g163(.A1(new_n542), .A2(KEYINPUT10), .A3(new_n587), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n581), .B1(new_n591), .B2(G868), .ZN(G284));
  OAI21_X1  g167(.A(new_n581), .B1(new_n591), .B2(G868), .ZN(G321));
  INV_X1    g168(.A(G868), .ZN(new_n594));
  NAND2_X1  g169(.A1(G299), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(G168), .B2(new_n594), .ZN(G297));
  OAI21_X1  g171(.A(new_n595), .B1(G168), .B2(new_n594), .ZN(G280));
  XOR2_X1   g172(.A(KEYINPUT76), .B(G559), .Z(new_n598));
  OAI21_X1  g173(.A(new_n591), .B1(G860), .B2(new_n598), .ZN(G148));
  NAND2_X1  g174(.A1(new_n591), .A2(new_n598), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(G868), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(G868), .B2(new_n545), .ZN(G323));
  XNOR2_X1  g177(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g178(.A1(new_n491), .A2(new_n466), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT12), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT13), .ZN(new_n606));
  XNOR2_X1  g181(.A(KEYINPUT77), .B(G2100), .ZN(new_n607));
  OR2_X1    g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n606), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n472), .A2(G135), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n474), .A2(G123), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n458), .A2(G111), .ZN(new_n612));
  OAI21_X1  g187(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n610), .B(new_n611), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(G2096), .Z(new_n615));
  NAND3_X1  g190(.A1(new_n608), .A2(new_n609), .A3(new_n615), .ZN(G156));
  XNOR2_X1  g191(.A(G2427), .B(G2438), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(G2430), .ZN(new_n618));
  XNOR2_X1  g193(.A(KEYINPUT15), .B(G2435), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n619), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n620), .A2(KEYINPUT14), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(G1341), .B(G1348), .ZN(new_n623));
  XNOR2_X1  g198(.A(G2443), .B(G2446), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n622), .B(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n628));
  XNOR2_X1  g203(.A(G2451), .B(G2454), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(G14), .B1(new_n627), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n632), .B1(new_n631), .B2(new_n627), .ZN(G401));
  XOR2_X1   g208(.A(G2072), .B(G2078), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT79), .ZN(new_n635));
  XOR2_X1   g210(.A(KEYINPUT81), .B(KEYINPUT17), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2067), .B(G2678), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2084), .B(G2090), .ZN(new_n639));
  NOR3_X1   g214(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n639), .B1(new_n635), .B2(new_n638), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n641), .B1(new_n637), .B2(new_n638), .ZN(new_n642));
  INV_X1    g217(.A(new_n638), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n643), .A2(new_n639), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n635), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT80), .B(KEYINPUT18), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NOR3_X1   g222(.A1(new_n640), .A2(new_n642), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2096), .B(G2100), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(G227));
  XNOR2_X1  g225(.A(G1956), .B(G2474), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT82), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1961), .B(G1966), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1971), .B(G1976), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT19), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT20), .Z(new_n659));
  NOR2_X1   g234(.A1(new_n652), .A2(new_n654), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n661), .A2(new_n657), .A3(new_n655), .ZN(new_n662));
  OAI211_X1 g237(.A(new_n659), .B(new_n662), .C1(new_n657), .C2(new_n661), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1991), .B(G1996), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1981), .B(G1986), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G229));
  NAND2_X1  g244(.A1(new_n472), .A2(G140), .ZN(new_n670));
  INV_X1    g245(.A(G128), .ZN(new_n671));
  INV_X1    g246(.A(new_n474), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g248(.A(G2104), .B1(new_n458), .B2(G116), .ZN(new_n674));
  OR3_X1    g249(.A1(KEYINPUT85), .A2(G104), .A3(G2105), .ZN(new_n675));
  OAI21_X1  g250(.A(KEYINPUT85), .B1(G104), .B2(G2105), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n674), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(G29), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT86), .ZN(new_n680));
  INV_X1    g255(.A(G29), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(G26), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT28), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G2067), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT31), .B(G11), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT30), .B(G28), .Z(new_n687));
  OAI21_X1  g262(.A(new_n686), .B1(new_n687), .B2(G29), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n614), .A2(new_n681), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n688), .B1(new_n689), .B2(KEYINPUT92), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(KEYINPUT92), .B2(new_n689), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT93), .Z(new_n692));
  NOR2_X1   g267(.A1(new_n685), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(G1348), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n591), .A2(G16), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G4), .B2(G16), .ZN(new_n696));
  INV_X1    g271(.A(G1961), .ZN(new_n697));
  NAND2_X1  g272(.A1(G301), .A2(G16), .ZN(new_n698));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G5), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  OAI221_X1 g276(.A(new_n693), .B1(new_n694), .B2(new_n696), .C1(new_n697), .C2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n681), .A2(G35), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G162), .B2(new_n681), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT29), .Z(new_n705));
  INV_X1    g280(.A(G2090), .ZN(new_n706));
  NOR2_X1   g281(.A1(G164), .A2(new_n681), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G27), .B2(new_n681), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  AOI22_X1  g284(.A1(new_n705), .A2(new_n706), .B1(G2078), .B2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT27), .B(G1996), .ZN(new_n711));
  NAND3_X1  g286(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT26), .Z(new_n713));
  INV_X1    g288(.A(G129), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n672), .B2(new_n714), .ZN(new_n715));
  AOI22_X1  g290(.A1(new_n472), .A2(G141), .B1(G105), .B2(new_n466), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT89), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G29), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G29), .B2(G32), .ZN(new_n721));
  OAI221_X1 g296(.A(new_n710), .B1(new_n706), .B2(new_n705), .C1(new_n711), .C2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G2078), .ZN(new_n723));
  INV_X1    g298(.A(G2084), .ZN(new_n724));
  INV_X1    g299(.A(G34), .ZN(new_n725));
  AOI21_X1  g300(.A(G29), .B1(new_n725), .B2(KEYINPUT24), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(KEYINPUT24), .B2(new_n725), .ZN(new_n727));
  INV_X1    g302(.A(G160), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n727), .B1(new_n728), .B2(new_n681), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n708), .A2(new_n723), .B1(new_n724), .B2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n701), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(G1961), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n699), .A2(G19), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(new_n545), .B2(new_n699), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(G1341), .Z(new_n735));
  INV_X1    g310(.A(G1956), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n699), .A2(G20), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT23), .Z(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G299), .B2(G16), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n735), .B1(new_n736), .B2(new_n739), .ZN(new_n740));
  NOR4_X1   g315(.A1(new_n702), .A2(new_n722), .A3(new_n732), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n696), .A2(new_n694), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n729), .A2(new_n724), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT88), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n681), .A2(G33), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT25), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G139), .B2(new_n472), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n491), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n458), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT87), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n745), .B1(new_n751), .B2(G29), .ZN(new_n752));
  INV_X1    g327(.A(G2072), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n744), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n721), .A2(new_n711), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n754), .B(new_n755), .C1(new_n753), .C2(new_n752), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n742), .B1(new_n756), .B2(KEYINPUT90), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(KEYINPUT90), .B2(new_n756), .ZN(new_n758));
  NAND2_X1  g333(.A1(G168), .A2(G16), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT91), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n759), .B(new_n760), .C1(G16), .C2(G21), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n760), .B2(new_n759), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n762), .A2(G1966), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n762), .A2(G1966), .ZN(new_n764));
  AOI211_X1 g339(.A(new_n763), .B(new_n764), .C1(new_n736), .C2(new_n739), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n741), .A2(new_n758), .A3(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n699), .A2(G24), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G290), .B2(G16), .ZN(new_n769));
  INV_X1    g344(.A(G1986), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n472), .A2(G131), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n474), .A2(G119), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n458), .A2(G107), .ZN(new_n775));
  OAI21_X1  g350(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n773), .B(new_n774), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  MUX2_X1   g352(.A(G25), .B(new_n777), .S(G29), .Z(new_n778));
  XOR2_X1   g353(.A(KEYINPUT35), .B(G1991), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n771), .A2(new_n772), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n699), .A2(G22), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G166), .B2(new_n699), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(G1971), .Z(new_n784));
  NAND2_X1  g359(.A1(new_n784), .A2(KEYINPUT83), .ZN(new_n785));
  MUX2_X1   g360(.A(G6), .B(G305), .S(G16), .Z(new_n786));
  XOR2_X1   g361(.A(KEYINPUT32), .B(G1981), .Z(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  MUX2_X1   g363(.A(G23), .B(G288), .S(G16), .Z(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT33), .B(G1976), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n785), .A2(new_n788), .A3(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT84), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n784), .A2(KEYINPUT83), .ZN(new_n794));
  OR3_X1    g369(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n793), .B1(new_n792), .B2(new_n794), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT34), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n781), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT36), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n795), .A2(KEYINPUT34), .A3(new_n796), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n800), .B1(new_n799), .B2(new_n801), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n767), .B1(new_n803), .B2(new_n804), .ZN(G150));
  INV_X1    g380(.A(G150), .ZN(G311));
  XNOR2_X1  g381(.A(KEYINPUT97), .B(G860), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n544), .A2(KEYINPUT95), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT96), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n502), .A2(G55), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT94), .B(G93), .ZN(new_n814));
  OAI221_X1 g389(.A(new_n812), .B1(new_n498), .B2(new_n813), .C1(new_n542), .C2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT95), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n545), .B2(new_n816), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n811), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n811), .A2(new_n817), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT38), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n591), .A2(G559), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT39), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n808), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n824), .B2(new_n823), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n815), .A2(new_n808), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT37), .Z(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n828), .ZN(G145));
  XNOR2_X1  g404(.A(new_n728), .B(new_n614), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(new_n478), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n490), .A2(new_n493), .ZN(new_n832));
  INV_X1    g407(.A(new_n485), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n472), .A2(G142), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n474), .A2(G130), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n458), .A2(G118), .ZN(new_n837));
  OAI21_X1  g412(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n835), .B(new_n836), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT99), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n777), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n605), .B(KEYINPUT98), .Z(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n678), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n843), .A2(new_n844), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n834), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n847), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n485), .B1(new_n490), .B2(new_n493), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n849), .A2(new_n850), .A3(new_n845), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n751), .A2(new_n718), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n719), .B2(new_n751), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n848), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n853), .B1(new_n848), .B2(new_n851), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n831), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(G37), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n848), .A2(new_n851), .ZN(new_n859));
  INV_X1    g434(.A(new_n853), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n831), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n861), .A2(new_n862), .A3(new_n854), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n857), .A2(new_n858), .A3(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g440(.A(G290), .B(G166), .ZN(new_n866));
  XOR2_X1   g441(.A(G288), .B(G305), .Z(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(new_n868));
  XOR2_X1   g443(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n820), .B(new_n600), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n590), .A2(G299), .ZN(new_n872));
  INV_X1    g447(.A(G299), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n586), .A2(new_n873), .A3(new_n588), .A4(new_n589), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT100), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n871), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT41), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n872), .A2(new_n878), .A3(new_n874), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT101), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n879), .B(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n875), .ZN(new_n882));
  OAI21_X1  g457(.A(KEYINPUT102), .B1(new_n882), .B2(new_n878), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT102), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n875), .A2(new_n884), .A3(KEYINPUT41), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n881), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n877), .B1(new_n871), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT104), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT104), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n877), .B(new_n889), .C1(new_n871), .C2(new_n886), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n870), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n890), .A2(new_n870), .ZN(new_n892));
  OAI21_X1  g467(.A(G868), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n815), .A2(new_n594), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(G295));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n894), .ZN(G331));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n897));
  OAI21_X1  g472(.A(G168), .B1(new_n897), .B2(G301), .ZN(new_n898));
  NAND2_X1  g473(.A1(G301), .A2(new_n897), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n898), .B(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n819), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n811), .A2(new_n817), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n898), .B(new_n899), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n818), .A2(new_n905), .A3(new_n819), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n904), .A2(new_n906), .A3(new_n882), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n904), .A2(new_n906), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n907), .B1(new_n886), .B2(new_n908), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n909), .A2(new_n868), .ZN(new_n910));
  AOI21_X1  g485(.A(G37), .B1(new_n909), .B2(new_n868), .ZN(new_n911));
  AOI21_X1  g486(.A(KEYINPUT43), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n886), .A2(new_n908), .ZN(new_n913));
  INV_X1    g488(.A(new_n907), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n913), .A2(new_n868), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n868), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n876), .A2(new_n906), .A3(new_n904), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n875), .A2(KEYINPUT41), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n908), .A2(new_n879), .A3(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n916), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  AND4_X1   g495(.A1(KEYINPUT43), .A2(new_n915), .A3(new_n858), .A4(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(KEYINPUT44), .B1(new_n912), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n924), .B1(new_n910), .B2(new_n911), .ZN(new_n925));
  AND4_X1   g500(.A1(new_n924), .A2(new_n915), .A3(new_n858), .A4(new_n920), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n922), .A2(new_n927), .ZN(G397));
  INV_X1    g503(.A(G1384), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n834), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT106), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT45), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n932), .B1(new_n931), .B2(new_n930), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n464), .A2(new_n467), .ZN(new_n934));
  INV_X1    g509(.A(G125), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n935), .B1(new_n470), .B2(new_n471), .ZN(new_n936));
  INV_X1    g511(.A(new_n462), .ZN(new_n937));
  OAI21_X1  g512(.A(G2105), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n934), .A2(new_n938), .A3(G40), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(G160), .A2(KEYINPUT107), .A3(G40), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n933), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n945), .A2(G1996), .ZN(new_n946));
  XOR2_X1   g521(.A(new_n946), .B(KEYINPUT46), .Z(new_n947));
  INV_X1    g522(.A(new_n718), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n678), .B(G2067), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n944), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT47), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n951), .B(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT126), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n951), .B(KEYINPUT47), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT126), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n949), .B1(G1996), .B2(new_n948), .ZN(new_n958));
  INV_X1    g533(.A(new_n719), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n958), .B1(G1996), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n779), .ZN(new_n961));
  OR3_X1    g536(.A1(new_n960), .A2(new_n961), .A3(new_n777), .ZN(new_n962));
  OR2_X1    g537(.A1(new_n678), .A2(G2067), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n945), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n777), .B(new_n961), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n960), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT48), .ZN(new_n968));
  OR3_X1    g543(.A1(new_n945), .A2(G290), .A3(G1986), .ZN(new_n969));
  AOI22_X1  g544(.A1(new_n967), .A2(new_n944), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OR2_X1    g545(.A1(new_n969), .A2(new_n968), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n964), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n955), .A2(new_n957), .A3(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT51), .ZN(new_n974));
  INV_X1    g549(.A(G8), .ZN(new_n975));
  AOI21_X1  g550(.A(G1384), .B1(new_n832), .B2(new_n833), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT50), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n978), .A2(new_n941), .A3(new_n942), .ZN(new_n979));
  INV_X1    g554(.A(new_n488), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT67), .B1(new_n480), .B2(new_n484), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n832), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n977), .B1(new_n982), .B2(new_n929), .ZN(new_n983));
  XOR2_X1   g558(.A(KEYINPUT116), .B(G2084), .Z(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n979), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT115), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n976), .A2(KEYINPUT45), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n987), .B1(new_n943), .B2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n982), .A2(KEYINPUT45), .A3(new_n929), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT45), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n991), .B1(new_n850), .B2(G1384), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n992), .A2(KEYINPUT115), .A3(new_n941), .A4(new_n942), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n989), .A2(new_n990), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G1966), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n986), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n975), .B1(new_n996), .B2(G168), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n993), .A2(new_n990), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(G1966), .B1(new_n999), .B2(new_n989), .ZN(new_n1000));
  OAI21_X1  g575(.A(G286), .B1(new_n1000), .B2(new_n986), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n974), .B1(new_n997), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT107), .B1(G160), .B2(G40), .ZN(new_n1003));
  AND4_X1   g578(.A1(KEYINPUT107), .A2(new_n934), .A3(new_n938), .A4(G40), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT115), .B1(new_n1005), .B2(new_n992), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n995), .B1(new_n998), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n986), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1007), .A2(G168), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(G8), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1010), .A2(KEYINPUT51), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT62), .B1(new_n1002), .B2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n996), .A2(G168), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT51), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT62), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n997), .A2(new_n974), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT108), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1018), .B(new_n991), .C1(G164), .C2(G1384), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n834), .A2(KEYINPUT45), .A3(new_n929), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT108), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT45), .B1(new_n982), .B2(new_n929), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1019), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(G1971), .B1(new_n1023), .B2(new_n1005), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n976), .A2(new_n977), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(new_n1005), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n982), .A2(new_n929), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1028), .A2(KEYINPUT50), .ZN(new_n1029));
  NOR3_X1   g604(.A1(new_n1027), .A2(G2090), .A3(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(G8), .B1(new_n1024), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(G8), .B1(new_n512), .B2(new_n518), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT109), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT109), .ZN(new_n1036));
  NAND4_X1  g611(.A1(G303), .A2(new_n1036), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1034), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1031), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1023), .A2(new_n723), .A3(new_n1005), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n1042));
  INV_X1    g617(.A(new_n979), .ZN(new_n1043));
  INV_X1    g618(.A(new_n983), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n1041), .A2(new_n1042), .B1(new_n1045), .B2(new_n697), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1042), .A2(G2078), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n999), .A2(new_n1047), .A3(new_n989), .ZN(new_n1048));
  AOI21_X1  g623(.A(G301), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n979), .A2(G2090), .A3(new_n983), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1038), .B(G8), .C1(new_n1024), .C2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n941), .A2(new_n942), .A3(new_n976), .ZN(new_n1052));
  AND2_X1   g627(.A1(new_n1052), .A2(G8), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT113), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1054), .A2(KEYINPUT49), .ZN(new_n1055));
  INV_X1    g630(.A(G1981), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n569), .A2(new_n573), .A3(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g632(.A(KEYINPUT112), .B(G86), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n516), .A2(new_n517), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1056), .B1(new_n1059), .B2(new_n573), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1055), .B1(new_n1057), .B2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n569), .A2(new_n573), .A3(new_n1056), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1055), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n1059), .A2(new_n573), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1062), .B(new_n1063), .C1(new_n1064), .C2(new_n1056), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1053), .A2(new_n1061), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G1976), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1052), .B(G8), .C1(new_n1067), .C2(G288), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT52), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1070));
  OR2_X1    g645(.A1(G288), .A2(new_n1067), .ZN(new_n1071));
  XOR2_X1   g646(.A(KEYINPUT110), .B(G1976), .Z(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT52), .B1(G288), .B2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1053), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT111), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT111), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1053), .A2(new_n1076), .A3(new_n1071), .A4(new_n1073), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1070), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  AND4_X1   g653(.A1(new_n1040), .A2(new_n1049), .A3(new_n1051), .A4(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1012), .A2(new_n1017), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT125), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT125), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1012), .A2(new_n1017), .A3(new_n1079), .A4(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n1085));
  NOR2_X1   g660(.A1(G288), .A2(G1976), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1066), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(new_n1062), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT114), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT114), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1087), .A2(new_n1090), .A3(new_n1062), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1089), .A2(new_n1053), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1051), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1078), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(G286), .A2(new_n975), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n996), .A2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1078), .A2(new_n1040), .A3(new_n1051), .A4(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT63), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n991), .B1(G164), .B2(G1384), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1018), .B1(new_n976), .B2(KEYINPUT45), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n943), .B1(new_n1105), .B2(new_n1019), .ZN(new_n1106));
  OAI22_X1  g681(.A1(new_n1106), .A2(G1971), .B1(new_n1045), .B2(G2090), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1038), .B1(new_n1107), .B2(G8), .ZN(new_n1108));
  OAI211_X1 g683(.A(KEYINPUT63), .B(new_n1097), .C1(new_n1000), .C2(new_n986), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1070), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1051), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1085), .B(new_n1096), .C1(new_n1102), .C2(new_n1114), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1100), .A2(new_n1101), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1116));
  OAI21_X1  g691(.A(KEYINPUT117), .B1(new_n1116), .B2(new_n1095), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1084), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT118), .ZN(new_n1120));
  AND3_X1   g695(.A1(G299), .A2(new_n1120), .A3(KEYINPUT57), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT57), .B1(G299), .B2(new_n1120), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT119), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT56), .B(G2072), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1023), .A2(new_n1125), .A3(new_n1005), .A4(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n736), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1125), .B1(new_n1106), .B2(new_n1126), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1124), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1023), .A2(new_n1005), .A3(new_n1126), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(KEYINPUT119), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1133), .A2(new_n1123), .A3(new_n1128), .A4(new_n1127), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1131), .A2(KEYINPUT61), .A3(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n943), .A2(G1996), .ZN(new_n1136));
  XOR2_X1   g711(.A(KEYINPUT58), .B(G1341), .Z(new_n1137));
  AOI22_X1  g712(.A1(new_n1023), .A2(new_n1136), .B1(new_n1052), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n1139));
  OAI22_X1  g714(.A1(new_n1138), .A2(new_n544), .B1(new_n1139), .B2(KEYINPUT59), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(KEYINPUT59), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n1141), .B(KEYINPUT121), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1142), .ZN(new_n1144));
  OAI221_X1 g719(.A(new_n1144), .B1(new_n1139), .B2(KEYINPUT59), .C1(new_n1138), .C2(new_n544), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n1135), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT122), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT61), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1148), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  AOI211_X1 g726(.A(KEYINPUT122), .B(KEYINPUT61), .C1(new_n1131), .C2(new_n1134), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1147), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT123), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT123), .ZN(new_n1155));
  OAI211_X1 g730(.A(new_n1147), .B(new_n1155), .C1(new_n1151), .C2(new_n1152), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1045), .A2(new_n694), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(G2067), .B2(new_n1052), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(KEYINPUT60), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(new_n591), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1161), .B1(KEYINPUT60), .B2(new_n1159), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1154), .A2(new_n1156), .A3(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1131), .B1(new_n1159), .B2(new_n590), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n1134), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT54), .ZN(new_n1167));
  INV_X1    g742(.A(new_n939), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n933), .A2(new_n1168), .A3(new_n1020), .A4(new_n1047), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1046), .A2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1170), .A2(G171), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1167), .B1(new_n1171), .B2(new_n1049), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1172), .A2(new_n1173), .A3(new_n1040), .A4(new_n1113), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1046), .A2(G301), .A3(new_n1048), .ZN(new_n1175));
  XOR2_X1   g750(.A(new_n1175), .B(KEYINPUT124), .Z(new_n1176));
  AOI21_X1  g751(.A(new_n1167), .B1(new_n1170), .B2(G171), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1174), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1119), .B1(new_n1166), .B2(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g754(.A(G290), .B(new_n770), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n945), .B1(new_n966), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n973), .B1(new_n1179), .B2(new_n1181), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g757(.A(G319), .ZN(new_n1184));
  NOR3_X1   g758(.A1(G401), .A2(G227), .A3(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g759(.A(new_n1185), .B(KEYINPUT127), .ZN(new_n1186));
  NOR2_X1   g760(.A1(G229), .A2(new_n1186), .ZN(new_n1187));
  OAI211_X1 g761(.A(new_n864), .B(new_n1187), .C1(new_n925), .C2(new_n926), .ZN(G225));
  INV_X1    g762(.A(G225), .ZN(G308));
endmodule


