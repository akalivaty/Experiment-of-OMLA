//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n549, new_n551, new_n552,
    new_n553, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n614, new_n616, new_n617, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1206, new_n1207, new_n1208,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT66), .ZN(new_n452));
  XOR2_X1   g027(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n454), .ZN(new_n458));
  INV_X1    g033(.A(new_n455), .ZN(new_n459));
  AOI22_X1  g034(.A1(new_n458), .A2(G2106), .B1(G567), .B2(new_n459), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n468), .A2(new_n470), .A3(G137), .ZN(new_n471));
  NAND2_X1  g046(.A1(G101), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(G2105), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n466), .A2(new_n473), .ZN(G160));
  INV_X1    g049(.A(new_n463), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(new_n462), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n475), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  NOR2_X1   g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(new_n462), .B2(G112), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n477), .B(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  NAND4_X1  g058(.A1(new_n468), .A2(new_n470), .A3(G138), .A4(new_n462), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT4), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n463), .A2(new_n486), .A3(G138), .A4(new_n462), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n468), .A2(new_n470), .A3(G126), .A4(G2105), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n463), .A2(KEYINPUT68), .A3(G126), .A4(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(KEYINPUT69), .B1(new_n462), .B2(G114), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n497), .A2(new_n498), .A3(G2105), .ZN(new_n499));
  AND3_X1   g074(.A1(new_n495), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  AND3_X1   g076(.A1(new_n488), .A2(new_n493), .A3(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT70), .A3(KEYINPUT5), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n505), .A2(new_n507), .B1(new_n504), .B2(G543), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT6), .B(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  INV_X1    g089(.A(G50), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n512), .A2(G543), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n511), .A2(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  INV_X1    g094(.A(new_n516), .ZN(new_n520));
  AND2_X1   g095(.A1(G63), .A2(G651), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n520), .A2(G51), .B1(new_n508), .B2(new_n521), .ZN(new_n522));
  XOR2_X1   g097(.A(KEYINPUT71), .B(KEYINPUT7), .Z(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n523), .B(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n508), .A2(G89), .A3(new_n512), .ZN(new_n526));
  AND3_X1   g101(.A1(new_n522), .A2(new_n525), .A3(new_n526), .ZN(G168));
  AND2_X1   g102(.A1(new_n508), .A2(new_n512), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n528), .A2(G90), .B1(G52), .B2(new_n520), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  OAI21_X1  g105(.A(KEYINPUT72), .B1(new_n530), .B2(new_n510), .ZN(new_n531));
  NAND2_X1  g106(.A1(G77), .A2(G543), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n505), .A2(new_n507), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n504), .A2(G543), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(G64), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n532), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT72), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n537), .A2(new_n538), .A3(G651), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n529), .A2(new_n531), .A3(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  AOI22_X1  g116(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n510), .ZN(new_n543));
  INV_X1    g118(.A(G81), .ZN(new_n544));
  INV_X1    g119(.A(G43), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n513), .A2(new_n544), .B1(new_n545), .B2(new_n516), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  XOR2_X1   g128(.A(new_n553), .B(KEYINPUT73), .Z(G188));
  NAND3_X1  g129(.A1(new_n512), .A2(G53), .A3(G543), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(KEYINPUT9), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n512), .A2(new_n557), .A3(G53), .A4(G543), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n508), .A2(G91), .A3(new_n512), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n508), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n561));
  OAI211_X1 g136(.A(new_n559), .B(new_n560), .C1(new_n510), .C2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(KEYINPUT74), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n535), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G651), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n567), .A2(new_n568), .A3(new_n560), .A4(new_n559), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n563), .A2(new_n569), .ZN(G299));
  NAND3_X1  g145(.A1(new_n522), .A2(new_n525), .A3(new_n526), .ZN(G286));
  NAND2_X1  g146(.A1(new_n520), .A2(G49), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n508), .A2(G87), .A3(new_n512), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G288));
  AND3_X1   g150(.A1(new_n506), .A2(KEYINPUT70), .A3(KEYINPUT5), .ZN(new_n576));
  AOI21_X1  g151(.A(KEYINPUT70), .B1(new_n506), .B2(KEYINPUT5), .ZN(new_n577));
  OAI211_X1 g152(.A(G61), .B(new_n534), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n510), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n533), .A2(G86), .A3(new_n534), .A4(new_n512), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n512), .A2(G48), .A3(G543), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G305));
  AOI22_X1  g160(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(new_n510), .ZN(new_n587));
  INV_X1    g162(.A(G85), .ZN(new_n588));
  INV_X1    g163(.A(G47), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n513), .A2(new_n588), .B1(new_n589), .B2(new_n516), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n535), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(G651), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n520), .A2(G54), .ZN(new_n598));
  AND2_X1   g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n508), .A2(G92), .A3(new_n512), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(KEYINPUT75), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT75), .ZN(new_n602));
  NAND4_X1  g177(.A1(new_n508), .A2(new_n602), .A3(G92), .A4(new_n512), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n601), .A2(KEYINPUT10), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n601), .A2(new_n603), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AND3_X1   g182(.A1(new_n599), .A2(new_n604), .A3(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n593), .B1(new_n608), .B2(G868), .ZN(G284));
  OAI21_X1  g184(.A(new_n593), .B1(new_n608), .B2(G868), .ZN(G321));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  MUX2_X1   g186(.A(G286), .B(G299), .S(new_n611), .Z(G280));
  XOR2_X1   g187(.A(G280), .B(KEYINPUT76), .Z(G297));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n608), .B1(new_n614), .B2(G860), .ZN(G148));
  NAND2_X1  g190(.A1(new_n608), .A2(new_n614), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G868), .B2(new_n547), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT77), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g195(.A1(new_n478), .A2(KEYINPUT78), .A3(G135), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT78), .ZN(new_n622));
  INV_X1    g197(.A(new_n478), .ZN(new_n623));
  INV_X1    g198(.A(G135), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n476), .A2(G123), .ZN(new_n626));
  OR2_X1    g201(.A1(G99), .A2(G2105), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n627), .B(G2104), .C1(G111), .C2(new_n462), .ZN(new_n628));
  NAND4_X1  g203(.A1(new_n621), .A2(new_n625), .A3(new_n626), .A4(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(G2096), .Z(new_n630));
  NAND3_X1  g205(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2100), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n630), .A2(new_n634), .ZN(G156));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2435), .ZN(new_n637));
  XOR2_X1   g212(.A(G2427), .B(G2438), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(KEYINPUT14), .ZN(new_n640));
  XOR2_X1   g215(.A(G2451), .B(G2454), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n640), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G1341), .B(G1348), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n645), .B(new_n646), .Z(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(G14), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(G401));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2067), .B(G2678), .Z(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(KEYINPUT18), .ZN(new_n654));
  XOR2_X1   g229(.A(G2072), .B(G2078), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT79), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2096), .B(G2100), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT80), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n657), .B(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT17), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(new_n651), .B2(new_n652), .ZN(new_n662));
  AOI21_X1  g237(.A(KEYINPUT18), .B1(new_n653), .B2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n660), .B(new_n663), .Z(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(G227));
  XOR2_X1   g240(.A(G1956), .B(G2474), .Z(new_n666));
  XOR2_X1   g241(.A(G1961), .B(G1966), .Z(new_n667));
  NOR2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1971), .B(G1976), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n666), .A2(new_n667), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT20), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n672), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n669), .A2(new_n671), .A3(new_n673), .ZN(new_n677));
  OAI211_X1 g252(.A(new_n676), .B(new_n677), .C1(new_n675), .C2(new_n674), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT81), .B(G1986), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT82), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n678), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(G1996), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1981), .B(G1991), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n681), .B(new_n685), .ZN(G229));
  INV_X1    g261(.A(KEYINPUT34), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT85), .B(G1981), .Z(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(G305), .A2(G16), .ZN(new_n690));
  INV_X1    g265(.A(G16), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G6), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n690), .A2(KEYINPUT32), .A3(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(KEYINPUT32), .B1(new_n690), .B2(new_n692), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n689), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n690), .A2(new_n692), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT32), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n699), .A2(new_n688), .A3(new_n693), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(G303), .A2(G16), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n691), .A2(G22), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G1971), .ZN(new_n705));
  OR2_X1    g280(.A1(G16), .A2(G23), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G288), .B2(new_n691), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT33), .B(G1976), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G1971), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n702), .A2(new_n710), .A3(new_n703), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n705), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n687), .B1(new_n701), .B2(new_n712), .ZN(new_n713));
  AND3_X1   g288(.A1(new_n705), .A2(new_n711), .A3(new_n709), .ZN(new_n714));
  NAND4_X1  g289(.A1(new_n714), .A2(KEYINPUT34), .A3(new_n700), .A4(new_n696), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G25), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n476), .A2(G119), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n478), .A2(G131), .ZN(new_n720));
  OR2_X1    g295(.A1(G95), .A2(G2105), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n721), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n719), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n718), .B1(new_n724), .B2(new_n717), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT83), .Z(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT35), .B(G1991), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n591), .B(KEYINPUT84), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G16), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G16), .B2(G24), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G1986), .ZN(new_n732));
  INV_X1    g307(.A(G1986), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n730), .B(new_n733), .C1(G16), .C2(G24), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n732), .A2(new_n734), .B1(new_n727), .B2(new_n726), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n716), .A2(new_n728), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(KEYINPUT36), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT36), .ZN(new_n738));
  NAND4_X1  g313(.A1(new_n716), .A2(new_n738), .A3(new_n728), .A4(new_n735), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT27), .B(G1996), .Z(new_n741));
  OR2_X1    g316(.A1(G29), .A2(G32), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT92), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n463), .A2(G129), .A3(G2105), .ZN(new_n746));
  NAND3_X1  g321(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT26), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n463), .A2(G141), .A3(new_n462), .ZN(new_n750));
  NAND4_X1  g325(.A1(new_n745), .A2(new_n746), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT93), .ZN(new_n752));
  AND3_X1   g327(.A1(new_n752), .A2(KEYINPUT94), .A3(G29), .ZN(new_n753));
  AOI21_X1  g328(.A(KEYINPUT94), .B1(new_n752), .B2(G29), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n741), .B(new_n742), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(G164), .A2(G29), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G27), .B2(G29), .ZN(new_n757));
  INV_X1    g332(.A(G2078), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT30), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n760), .A2(G28), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(G28), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n761), .A2(new_n762), .A3(new_n717), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n755), .A2(new_n759), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(G299), .A2(G16), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n691), .A2(KEYINPUT23), .A3(G20), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT23), .ZN(new_n767));
  INV_X1    g342(.A(G20), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(new_n768), .B2(G16), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n765), .A2(new_n766), .A3(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(G1956), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n764), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OR3_X1    g349(.A1(G286), .A2(KEYINPUT95), .A3(new_n691), .ZN(new_n775));
  NOR2_X1   g350(.A1(G286), .A2(new_n691), .ZN(new_n776));
  OAI21_X1  g351(.A(KEYINPUT95), .B1(G16), .B2(G21), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(G1966), .ZN(new_n779));
  INV_X1    g354(.A(G1966), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n775), .B(new_n780), .C1(new_n776), .C2(new_n777), .ZN(new_n781));
  INV_X1    g356(.A(G1341), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n547), .A2(G16), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G16), .B2(G19), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n779), .B(new_n781), .C1(new_n782), .C2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT28), .ZN(new_n786));
  INV_X1    g361(.A(G26), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(new_n787), .B2(G29), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n787), .A2(G29), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n463), .A2(G128), .A3(G2105), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n463), .A2(G140), .A3(new_n462), .ZN(new_n791));
  OR2_X1    g366(.A1(G104), .A2(G2105), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n792), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n790), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n789), .B1(new_n794), .B2(G29), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n788), .B1(new_n795), .B2(new_n786), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT87), .ZN(new_n797));
  INV_X1    g372(.A(G2067), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n785), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n608), .A2(G16), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G4), .B2(G16), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT86), .B(G1348), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n691), .A2(G5), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G171), .B2(new_n691), .ZN(new_n806));
  INV_X1    g381(.A(G1961), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n774), .A2(new_n800), .A3(new_n804), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n717), .A2(G35), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G162), .B2(new_n717), .ZN(new_n811));
  MUX2_X1   g386(.A(new_n810), .B(new_n811), .S(KEYINPUT97), .Z(new_n812));
  XOR2_X1   g387(.A(KEYINPUT29), .B(G2090), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT24), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n717), .B1(new_n815), .B2(G34), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n816), .A2(KEYINPUT91), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n816), .A2(KEYINPUT91), .ZN(new_n818));
  AOI211_X1 g393(.A(new_n817), .B(new_n818), .C1(new_n815), .C2(G34), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(G160), .B2(G29), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n820), .A2(G2084), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT96), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT31), .B(G11), .Z(new_n823));
  INV_X1    g398(.A(new_n757), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n823), .B1(new_n824), .B2(G2078), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n814), .A2(new_n822), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n742), .B1(new_n753), .B2(new_n754), .ZN(new_n827));
  INV_X1    g402(.A(new_n741), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n827), .A2(new_n828), .B1(G2084), .B2(new_n820), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n802), .A2(new_n803), .ZN(new_n831));
  NOR4_X1   g406(.A1(new_n809), .A2(new_n826), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n717), .A2(G33), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n478), .A2(G139), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n835), .A2(new_n462), .ZN(new_n836));
  XNOR2_X1  g411(.A(KEYINPUT88), .B(KEYINPUT25), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n834), .A2(new_n836), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n833), .B1(new_n840), .B2(new_n717), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT89), .ZN(new_n842));
  INV_X1    g417(.A(G2072), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT90), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n784), .A2(new_n782), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n740), .A2(new_n832), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n842), .A2(new_n843), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n629), .A2(new_n717), .ZN(new_n849));
  NOR3_X1   g424(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(G311));
  OR3_X1    g425(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(G150));
  AOI22_X1  g426(.A1(new_n528), .A2(G93), .B1(G55), .B2(new_n520), .ZN(new_n852));
  AOI22_X1  g427(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n852), .B1(new_n510), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(G860), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(KEYINPUT37), .Z(new_n856));
  NAND2_X1  g431(.A1(new_n608), .A2(G559), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT38), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT39), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n852), .B(KEYINPUT98), .C1(new_n510), .C2(new_n853), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT98), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n853), .A2(new_n510), .ZN(new_n862));
  INV_X1    g437(.A(G93), .ZN(new_n863));
  INV_X1    g438(.A(G55), .ZN(new_n864));
  OAI22_X1  g439(.A1(new_n513), .A2(new_n863), .B1(new_n864), .B2(new_n516), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n861), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n860), .A2(new_n547), .A3(new_n866), .ZN(new_n867));
  OAI221_X1 g442(.A(new_n861), .B1(new_n543), .B2(new_n546), .C1(new_n862), .C2(new_n865), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n859), .B(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n856), .B1(new_n871), .B2(G860), .ZN(G145));
  XNOR2_X1  g447(.A(new_n629), .B(G160), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(G162), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n794), .A2(KEYINPUT99), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT99), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n790), .A2(new_n791), .A3(new_n876), .A4(new_n793), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(G164), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n488), .A2(new_n493), .A3(new_n501), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n880), .A2(new_n875), .A3(new_n877), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n751), .B(KEYINPUT93), .Z(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n752), .A2(new_n879), .A3(new_n881), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(new_n840), .A3(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT100), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n751), .B1(new_n879), .B2(new_n881), .ZN(new_n888));
  INV_X1    g463(.A(new_n840), .ZN(new_n889));
  INV_X1    g464(.A(new_n751), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n889), .B1(new_n882), .B2(new_n890), .ZN(new_n891));
  OAI211_X1 g466(.A(new_n886), .B(new_n887), .C1(new_n888), .C2(new_n891), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n884), .A2(KEYINPUT100), .A3(new_n840), .A4(new_n885), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n476), .A2(G130), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n478), .A2(G142), .ZN(new_n896));
  NOR2_X1   g471(.A1(G106), .A2(G2105), .ZN(new_n897));
  OAI21_X1  g472(.A(G2104), .B1(new_n462), .B2(G118), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n895), .B(new_n896), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  XOR2_X1   g474(.A(new_n899), .B(new_n632), .Z(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(new_n724), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n874), .B1(new_n894), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n892), .A2(new_n901), .A3(new_n893), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT102), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT102), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n892), .A2(new_n901), .A3(new_n906), .A4(new_n893), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n903), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT103), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT103), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n903), .A2(new_n905), .A3(new_n910), .A4(new_n907), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(G37), .ZN(new_n913));
  AOI211_X1 g488(.A(KEYINPUT101), .B(new_n901), .C1(new_n892), .C2(new_n893), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT101), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n915), .B1(new_n894), .B2(new_n902), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n904), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n874), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n912), .A2(new_n913), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT40), .ZN(new_n920));
  AOI21_X1  g495(.A(G37), .B1(new_n909), .B2(new_n911), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT40), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(new_n922), .A3(new_n918), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n920), .A2(new_n923), .ZN(G395));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n563), .A2(new_n925), .A3(new_n569), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n608), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n925), .B1(new_n563), .B2(new_n569), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n599), .A2(new_n607), .A3(new_n604), .ZN(new_n930));
  NAND3_X1  g505(.A1(G299), .A2(new_n930), .A3(KEYINPUT104), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT41), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(G299), .A2(KEYINPUT104), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n934), .A2(new_n608), .A3(new_n926), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT41), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n935), .A2(new_n936), .A3(new_n931), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n933), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n929), .A2(new_n932), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n616), .B(new_n869), .ZN(new_n940));
  MUX2_X1   g515(.A(new_n938), .B(new_n939), .S(new_n940), .Z(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(KEYINPUT105), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT105), .B1(new_n940), .B2(new_n939), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(G303), .B(G288), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n945), .A2(G305), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n945), .A2(G305), .ZN(new_n947));
  OAI21_X1  g522(.A(G290), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  OR2_X1    g523(.A1(new_n945), .A2(G305), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n945), .A2(G305), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(new_n591), .A3(new_n950), .ZN(new_n951));
  AND2_X1   g526(.A1(KEYINPUT106), .A2(KEYINPUT42), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n948), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(KEYINPUT106), .A2(KEYINPUT42), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n955), .B(KEYINPUT107), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n954), .B(new_n957), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n942), .A2(new_n944), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n958), .B1(new_n942), .B2(new_n944), .ZN(new_n960));
  OAI21_X1  g535(.A(G868), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n854), .A2(new_n611), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(G295));
  NAND2_X1  g538(.A1(new_n961), .A2(new_n962), .ZN(G331));
  NAND2_X1  g539(.A1(new_n948), .A2(new_n951), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT109), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n933), .A2(new_n966), .A3(new_n937), .ZN(new_n967));
  NAND3_X1  g542(.A1(G171), .A2(KEYINPUT108), .A3(G168), .ZN(new_n968));
  NAND2_X1  g543(.A1(G168), .A2(KEYINPUT108), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT108), .ZN(new_n970));
  NAND2_X1  g545(.A1(G286), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n969), .A2(new_n971), .A3(G301), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n968), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n869), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n968), .A2(new_n972), .A3(new_n868), .A4(new_n867), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n935), .A2(new_n936), .A3(new_n931), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT109), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n967), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n939), .A2(new_n975), .A3(new_n974), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n965), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n936), .B1(new_n935), .B2(new_n931), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n976), .B1(new_n977), .B2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n983), .A2(new_n965), .A3(new_n980), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n913), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT43), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n981), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  AND4_X1   g562(.A1(new_n931), .A2(new_n974), .A3(new_n935), .A4(new_n975), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(new_n938), .B2(new_n976), .ZN(new_n989));
  AOI21_X1  g564(.A(G37), .B1(new_n989), .B2(new_n965), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n983), .A2(new_n980), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n991), .A2(new_n951), .A3(new_n948), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT43), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(KEYINPUT44), .B1(new_n987), .B2(new_n993), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n981), .A2(new_n985), .A3(KEYINPUT43), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n986), .B1(new_n990), .B2(new_n992), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n994), .B1(new_n997), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g573(.A(G1384), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n880), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G40), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n466), .A2(new_n1001), .A3(new_n473), .ZN(new_n1002));
  XOR2_X1   g577(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1000), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n794), .B(new_n798), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G1996), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1007), .B1(new_n752), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(new_n1008), .B2(new_n890), .ZN(new_n1010));
  OR3_X1    g585(.A1(new_n1010), .A2(new_n727), .A3(new_n723), .ZN(new_n1011));
  OR2_X1    g586(.A1(new_n794), .A2(G2067), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1005), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1005), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1014), .B1(new_n751), .B2(new_n1007), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1014), .A2(KEYINPUT46), .A3(new_n1008), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT46), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1017), .B1(new_n1005), .B2(G1996), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1015), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  XOR2_X1   g594(.A(new_n1019), .B(KEYINPUT47), .Z(new_n1020));
  XOR2_X1   g595(.A(new_n723), .B(new_n727), .Z(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1014), .B1(new_n1010), .B2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1014), .A2(new_n733), .A3(new_n591), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n1024), .B(KEYINPUT48), .ZN(new_n1025));
  AOI211_X1 g600(.A(new_n1013), .B(new_n1020), .C1(new_n1023), .C2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(KEYINPUT113), .A2(KEYINPUT49), .ZN(new_n1027));
  OAI21_X1  g602(.A(G1981), .B1(new_n580), .B2(new_n583), .ZN(new_n1028));
  OR2_X1    g603(.A1(KEYINPUT113), .A2(KEYINPUT49), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NOR3_X1   g605(.A1(new_n580), .A2(new_n583), .A3(G1981), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1027), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G1981), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n584), .A2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1034), .A2(KEYINPUT113), .A3(KEYINPUT49), .A4(new_n1028), .ZN(new_n1035));
  INV_X1    g610(.A(G8), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n500), .B1(new_n491), .B2(new_n492), .ZN(new_n1037));
  AOI21_X1  g612(.A(G1384), .B1(new_n1037), .B2(new_n488), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1036), .B1(new_n1038), .B2(new_n1002), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1032), .A2(new_n1035), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G288), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(G1976), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1039), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT52), .ZN(new_n1044));
  XNOR2_X1  g619(.A(KEYINPUT112), .B(G1976), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT52), .B1(G288), .B2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1039), .A2(new_n1042), .A3(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1040), .A2(new_n1044), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT116), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1040), .A2(new_n1044), .A3(new_n1050), .A4(new_n1047), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT115), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT50), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1054), .B1(new_n880), .B2(new_n999), .ZN(new_n1055));
  INV_X1    g630(.A(new_n473), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n464), .A2(new_n465), .ZN(new_n1057));
  OAI211_X1 g632(.A(G40), .B(new_n1056), .C1(new_n1057), .C2(new_n462), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1053), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G2090), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1038), .A2(new_n1054), .ZN(new_n1061));
  OAI211_X1 g636(.A(KEYINPUT115), .B(new_n1002), .C1(new_n1038), .C2(new_n1054), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1058), .B1(new_n1038), .B2(KEYINPUT45), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1000), .A2(new_n1004), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n710), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1063), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(G8), .ZN(new_n1069));
  NAND2_X1  g644(.A1(G303), .A2(G8), .ZN(new_n1070));
  XNOR2_X1  g645(.A(new_n1070), .B(KEYINPUT55), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1071), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1058), .B1(new_n1055), .B2(KEYINPUT111), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT111), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1075), .B1(new_n1038), .B2(new_n1054), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1074), .A2(new_n1061), .A3(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1067), .B1(new_n1077), .B2(G2090), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1073), .A2(G8), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G2084), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1074), .A2(new_n1080), .A3(new_n1061), .A4(new_n1076), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1002), .B1(new_n1000), .B2(new_n1004), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1038), .A2(KEYINPUT45), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n780), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AOI211_X1 g659(.A(new_n1036), .B(G286), .C1(new_n1081), .C2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1052), .A2(new_n1072), .A3(new_n1079), .A4(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT63), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1078), .A2(G8), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1087), .B1(new_n1089), .B2(new_n1071), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1048), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1090), .A2(new_n1079), .A3(new_n1091), .A4(new_n1085), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1088), .A2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1079), .A2(new_n1048), .ZN(new_n1094));
  INV_X1    g669(.A(G1976), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1040), .A2(new_n1095), .A3(new_n1041), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n1031), .B(KEYINPUT114), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1094), .B1(new_n1039), .B2(new_n1098), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1052), .A2(new_n1079), .A3(new_n1072), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1064), .A2(new_n1065), .A3(new_n758), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1000), .A2(KEYINPUT111), .A3(KEYINPUT50), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(new_n1002), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1061), .B1(new_n1055), .B2(KEYINPUT111), .ZN(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT120), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT120), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1074), .A2(new_n1108), .A3(new_n1061), .A4(new_n1076), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1107), .A2(new_n807), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT125), .ZN(new_n1111));
  OR4_X1    g686(.A1(new_n1102), .A2(new_n1082), .A3(G2078), .A4(new_n1083), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1111), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1103), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1081), .A2(G168), .A3(new_n1084), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(G8), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT51), .ZN(new_n1118));
  AOI21_X1  g693(.A(G168), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT51), .ZN(new_n1120));
  OAI211_X1 g695(.A(G8), .B(new_n1116), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT62), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1118), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1100), .A2(new_n1115), .A3(G171), .A4(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1122), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1093), .B(new_n1099), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT125), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n1129), .A2(new_n1130), .B1(new_n1102), .B2(new_n1101), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1127), .B1(new_n1131), .B2(G301), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1110), .A2(KEYINPUT126), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1101), .B(KEYINPUT53), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT126), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1107), .A2(new_n1135), .A3(new_n1109), .A4(new_n807), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1133), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT127), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT127), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1133), .A2(new_n1139), .A3(new_n1134), .A4(new_n1136), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1138), .A2(G171), .A3(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1107), .A2(new_n803), .A3(new_n1109), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1038), .A2(new_n1002), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT118), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1038), .A2(KEYINPUT118), .A3(new_n1002), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1145), .A2(new_n798), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(KEYINPUT119), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT119), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1145), .A2(new_n1149), .A3(new_n798), .A4(new_n1146), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1142), .A2(new_n1151), .A3(new_n930), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n930), .B1(new_n1142), .B2(new_n1151), .ZN(new_n1153));
  OAI21_X1  g728(.A(KEYINPUT60), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n1142), .A2(new_n1151), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n930), .A2(KEYINPUT60), .ZN(new_n1156));
  XOR2_X1   g731(.A(KEYINPUT122), .B(G1996), .Z(new_n1157));
  INV_X1    g732(.A(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1064), .A2(new_n1065), .A3(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  XOR2_X1   g735(.A(KEYINPUT58), .B(G1341), .Z(new_n1161));
  INV_X1    g736(.A(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1162), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1163));
  OAI211_X1 g738(.A(KEYINPUT123), .B(new_n547), .C1(new_n1160), .C2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(KEYINPUT59), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1146), .ZN(new_n1166));
  AOI21_X1  g741(.A(KEYINPUT118), .B1(new_n1038), .B2(new_n1002), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1161), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(new_n1159), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT59), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1169), .A2(KEYINPUT123), .A3(new_n1170), .A4(new_n547), .ZN(new_n1171));
  AOI22_X1  g746(.A1(new_n1155), .A2(new_n1156), .B1(new_n1165), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT61), .ZN(new_n1173));
  XOR2_X1   g748(.A(KEYINPUT56), .B(G2072), .Z(new_n1174));
  OAI21_X1  g749(.A(KEYINPUT117), .B1(new_n1066), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT117), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1174), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1064), .A2(new_n1065), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1175), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1059), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(new_n771), .ZN(new_n1181));
  XOR2_X1   g756(.A(new_n562), .B(KEYINPUT57), .Z(new_n1182));
  NAND3_X1  g757(.A1(new_n1179), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1182), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1173), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  AND2_X1   g761(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n1182), .B(KEYINPUT121), .ZN(new_n1188));
  OAI211_X1 g763(.A(KEYINPUT61), .B(new_n1183), .C1(new_n1187), .C2(new_n1188), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1154), .A2(new_n1172), .A3(new_n1186), .A4(new_n1189), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1191), .B1(new_n1153), .B2(new_n1183), .ZN(new_n1192));
  AOI22_X1  g767(.A1(new_n1132), .A2(new_n1141), .B1(new_n1190), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1100), .A2(new_n1194), .ZN(new_n1195));
  OR2_X1    g770(.A1(new_n1137), .A2(G171), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1196), .B1(new_n1131), .B2(G301), .ZN(new_n1197));
  XOR2_X1   g772(.A(KEYINPUT124), .B(KEYINPUT54), .Z(new_n1198));
  AOI21_X1  g773(.A(new_n1195), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1126), .B1(new_n1193), .B2(new_n1199), .ZN(new_n1200));
  NOR2_X1   g775(.A1(new_n1010), .A2(new_n1022), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n591), .B(G1986), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1005), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1026), .B1(new_n1200), .B2(new_n1203), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g779(.A(G229), .ZN(new_n1206));
  NAND3_X1  g780(.A1(new_n919), .A2(new_n664), .A3(new_n1206), .ZN(new_n1207));
  OAI211_X1 g781(.A(G319), .B(new_n648), .C1(new_n995), .C2(new_n996), .ZN(new_n1208));
  NOR2_X1   g782(.A1(new_n1207), .A2(new_n1208), .ZN(G308));
  INV_X1    g783(.A(G319), .ZN(new_n1210));
  AND2_X1   g784(.A1(new_n979), .A2(new_n980), .ZN(new_n1211));
  OAI211_X1 g785(.A(new_n986), .B(new_n990), .C1(new_n1211), .C2(new_n965), .ZN(new_n1212));
  NOR2_X1   g786(.A1(new_n989), .A2(new_n965), .ZN(new_n1213));
  OAI21_X1  g787(.A(KEYINPUT43), .B1(new_n1213), .B2(new_n985), .ZN(new_n1214));
  AOI21_X1  g788(.A(new_n1210), .B1(new_n1212), .B2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g789(.A(G227), .B1(new_n921), .B2(new_n918), .ZN(new_n1216));
  NAND4_X1  g790(.A1(new_n1215), .A2(new_n1216), .A3(new_n648), .A4(new_n1206), .ZN(G225));
endmodule


