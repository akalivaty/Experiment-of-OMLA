//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 1 1 0 0 1 1 0 1 1 0 0 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 1 0 0 1 1 0 0 1 0 0 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014;
  XNOR2_X1  g000(.A(G125), .B(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT16), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  OR3_X1    g003(.A1(new_n189), .A2(KEYINPUT16), .A3(G140), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n188), .A2(G146), .A3(new_n190), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G119), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT72), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G119), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G128), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT72), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n199), .B1(new_n197), .B2(new_n202), .ZN(new_n203));
  XOR2_X1   g017(.A(KEYINPUT24), .B(G110), .Z(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n197), .A2(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n196), .A2(KEYINPUT23), .A3(G119), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n201), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G110), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n195), .A2(new_n205), .A3(new_n210), .ZN(new_n211));
  OAI22_X1  g025(.A1(new_n203), .A2(new_n204), .B1(new_n209), .B2(G110), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT73), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n194), .A2(new_n213), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n188), .A2(KEYINPUT73), .A3(G146), .A4(new_n190), .ZN(new_n215));
  OR2_X1    g029(.A1(KEYINPUT64), .A2(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(KEYINPUT64), .A2(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(new_n187), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n212), .A2(new_n214), .A3(new_n215), .A4(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n211), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT22), .B(G137), .ZN(new_n222));
  INV_X1    g036(.A(G953), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n223), .A2(G221), .A3(G234), .ZN(new_n224));
  XOR2_X1   g038(.A(new_n222), .B(new_n224), .Z(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n221), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n211), .A2(new_n220), .A3(new_n225), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  OR3_X1    g044(.A1(new_n230), .A2(KEYINPUT25), .A3(G902), .ZN(new_n231));
  INV_X1    g045(.A(G217), .ZN(new_n232));
  INV_X1    g046(.A(G902), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n232), .B1(G234), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(KEYINPUT25), .B1(new_n230), .B2(G902), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n231), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n234), .A2(G902), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n229), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT74), .ZN(new_n239));
  OR2_X1    g053(.A1(new_n238), .A2(KEYINPUT74), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n236), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(G472), .A2(G902), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n242), .B(KEYINPUT70), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G134), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G137), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT66), .ZN(new_n247));
  INV_X1    g061(.A(G137), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G134), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n246), .A2(KEYINPUT66), .ZN(new_n251));
  OAI21_X1  g065(.A(G131), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT11), .B1(new_n245), .B2(G137), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT11), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(new_n248), .A3(G134), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G131), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n256), .A2(new_n257), .A3(new_n246), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n252), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G143), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n261), .B1(new_n216), .B2(new_n217), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT1), .ZN(new_n263));
  OAI21_X1  g077(.A(G128), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n261), .A2(G146), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n266), .B1(new_n218), .B2(G143), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  AND2_X1   g082(.A1(KEYINPUT64), .A2(G146), .ZN(new_n269));
  NOR2_X1   g083(.A1(KEYINPUT64), .A2(G146), .ZN(new_n270));
  OAI21_X1  g084(.A(G143), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n192), .A2(G143), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n271), .A2(new_n263), .A3(G128), .A4(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(KEYINPUT67), .B1(new_n268), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n196), .B1(new_n271), .B2(KEYINPUT1), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n269), .A2(new_n270), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n265), .B1(new_n277), .B2(new_n261), .ZN(new_n278));
  OAI211_X1 g092(.A(KEYINPUT67), .B(new_n274), .C1(new_n276), .C2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n260), .B1(new_n275), .B2(new_n280), .ZN(new_n281));
  AND3_X1   g095(.A1(new_n256), .A2(new_n257), .A3(new_n246), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n257), .B1(new_n256), .B2(new_n246), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  XOR2_X1   g098(.A(KEYINPUT0), .B(G128), .Z(new_n285));
  NOR3_X1   g099(.A1(new_n269), .A2(new_n270), .A3(G143), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n285), .B1(new_n286), .B2(new_n265), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n271), .A2(KEYINPUT0), .A3(G128), .A4(new_n273), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n284), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n281), .A2(KEYINPUT30), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT30), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n287), .A2(KEYINPUT65), .A3(new_n288), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT65), .B1(new_n287), .B2(new_n288), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n294), .A2(new_n295), .A3(new_n284), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n259), .B1(new_n268), .B2(new_n274), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n293), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  XOR2_X1   g112(.A(G116), .B(G119), .Z(new_n299));
  XNOR2_X1  g113(.A(KEYINPUT2), .B(G113), .ZN(new_n300));
  OR2_X1    g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n300), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n292), .A2(new_n298), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n303), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n281), .A2(new_n305), .A3(new_n291), .ZN(new_n306));
  NOR2_X1   g120(.A1(G237), .A2(G953), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G210), .ZN(new_n308));
  INV_X1    g122(.A(G101), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n308), .B(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n311));
  XOR2_X1   g125(.A(new_n310), .B(new_n311), .Z(new_n312));
  NAND3_X1  g126(.A1(new_n304), .A2(new_n306), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT31), .ZN(new_n314));
  XOR2_X1   g128(.A(KEYINPUT68), .B(KEYINPUT31), .Z(new_n315));
  NAND4_X1  g129(.A1(new_n304), .A2(new_n306), .A3(new_n312), .A4(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT69), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT65), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n289), .A2(new_n319), .ZN(new_n320));
  OR2_X1    g134(.A1(new_n282), .A2(new_n283), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n287), .A2(KEYINPUT65), .A3(new_n288), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n274), .B1(new_n276), .B2(new_n278), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n260), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n305), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n306), .B1(new_n318), .B2(new_n326), .ZN(new_n327));
  AOI211_X1 g141(.A(KEYINPUT69), .B(new_n305), .C1(new_n323), .C2(new_n325), .ZN(new_n328));
  OAI21_X1  g142(.A(KEYINPUT28), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT67), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n324), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n259), .B1(new_n331), .B2(new_n279), .ZN(new_n332));
  NOR3_X1   g146(.A1(new_n332), .A2(new_n290), .A3(new_n303), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n333), .A2(KEYINPUT28), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n312), .B1(new_n329), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n244), .B1(new_n317), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT32), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n296), .A2(new_n297), .ZN(new_n340));
  OAI21_X1  g154(.A(KEYINPUT69), .B1(new_n340), .B2(new_n305), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n326), .A2(new_n318), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n341), .A2(new_n306), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n334), .B1(new_n343), .B2(KEYINPUT28), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n314), .B(new_n316), .C1(new_n344), .C2(new_n312), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(KEYINPUT32), .A3(new_n244), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n339), .A2(KEYINPUT71), .A3(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT71), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n337), .A2(new_n348), .A3(new_n338), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n344), .A2(new_n312), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT29), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n304), .A2(new_n306), .ZN(new_n353));
  INV_X1    g167(.A(new_n312), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n351), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT28), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n303), .B1(new_n332), .B2(new_n290), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n357), .B1(new_n306), .B2(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n359), .A2(new_n334), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n354), .A2(new_n352), .ZN(new_n361));
  AOI21_X1  g175(.A(G902), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n356), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G472), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n241), .B1(new_n350), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G952), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n366), .A2(G953), .ZN(new_n367));
  NAND2_X1  g181(.A1(G234), .A2(G237), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  XOR2_X1   g184(.A(KEYINPUT21), .B(G898), .Z(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n368), .A2(G902), .A3(G953), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n370), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(G214), .B1(G237), .B2(G902), .ZN(new_n377));
  OAI21_X1  g191(.A(G210), .B1(G237), .B2(G902), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n289), .A2(G125), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n379), .B1(G125), .B2(new_n324), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n223), .A2(G224), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(KEYINPUT79), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n380), .B(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT6), .ZN(new_n385));
  INV_X1    g199(.A(G104), .ZN(new_n386));
  OAI21_X1  g200(.A(KEYINPUT3), .B1(new_n386), .B2(G107), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT3), .ZN(new_n388));
  INV_X1    g202(.A(G107), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n389), .A3(G104), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n386), .A2(G107), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n387), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G101), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n387), .A2(new_n390), .A3(new_n309), .A4(new_n391), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(KEYINPUT4), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT75), .ZN(new_n396));
  OR2_X1    g210(.A1(new_n393), .A2(KEYINPUT4), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT75), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n393), .A2(new_n398), .A3(KEYINPUT4), .A4(new_n394), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n396), .A2(new_n303), .A3(new_n397), .A4(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT76), .ZN(new_n401));
  XNOR2_X1  g215(.A(G104), .B(G107), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n401), .B1(new_n402), .B2(new_n309), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n389), .A2(G104), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n391), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(KEYINPUT76), .A3(G101), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n403), .A2(new_n406), .A3(new_n394), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT5), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(new_n200), .A3(G116), .ZN(new_n409));
  OAI211_X1 g223(.A(G113), .B(new_n409), .C1(new_n299), .C2(new_n408), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n407), .A2(new_n301), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n400), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT78), .ZN(new_n413));
  XOR2_X1   g227(.A(G110), .B(G122), .Z(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n414), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n400), .A2(new_n416), .A3(new_n411), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n385), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  AOI211_X1 g232(.A(KEYINPUT78), .B(new_n416), .C1(new_n400), .C2(new_n411), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n419), .A2(KEYINPUT6), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n384), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT80), .ZN(new_n422));
  INV_X1    g236(.A(new_n417), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT6), .B1(new_n419), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n415), .A2(new_n385), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT80), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n427), .A3(new_n384), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n422), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT8), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n410), .A2(new_n301), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n407), .B(new_n431), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n412), .B(new_n416), .C1(new_n430), .C2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n414), .B1(new_n432), .B2(KEYINPUT8), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n382), .A2(KEYINPUT7), .ZN(new_n436));
  XOR2_X1   g250(.A(new_n380), .B(new_n436), .Z(new_n437));
  NAND2_X1  g251(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n233), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n378), .B1(new_n429), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n378), .ZN(new_n442));
  AOI211_X1 g256(.A(new_n442), .B(new_n439), .C1(new_n422), .C2(new_n428), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n376), .B(new_n377), .C1(new_n441), .C2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G469), .ZN(new_n445));
  XNOR2_X1  g259(.A(G110), .B(G140), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n223), .A2(G227), .ZN(new_n447));
  XOR2_X1   g261(.A(new_n446), .B(new_n447), .Z(new_n448));
  OAI211_X1 g262(.A(KEYINPUT10), .B(new_n407), .C1(new_n275), .C2(new_n280), .ZN(new_n449));
  OAI21_X1  g263(.A(G128), .B1(new_n265), .B2(new_n263), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n450), .B(KEYINPUT77), .C1(new_n262), .C2(new_n272), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n274), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n271), .A2(new_n273), .ZN(new_n453));
  AOI21_X1  g267(.A(KEYINPUT77), .B1(new_n453), .B2(new_n450), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n407), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT10), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n289), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n396), .A2(new_n458), .A3(new_n397), .A4(new_n399), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n449), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n321), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n449), .A2(new_n284), .A3(new_n457), .A4(new_n459), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n448), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n448), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n403), .A2(new_n406), .A3(new_n394), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n268), .A2(new_n274), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n455), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(KEYINPUT12), .B1(new_n467), .B2(new_n321), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT12), .ZN(new_n469));
  AOI211_X1 g283(.A(new_n469), .B(new_n284), .C1(new_n455), .C2(new_n466), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n464), .A2(new_n471), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n445), .B(new_n233), .C1(new_n463), .C2(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n445), .A2(new_n233), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n462), .B1(new_n470), .B2(new_n468), .ZN(new_n476));
  INV_X1    g290(.A(new_n448), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n461), .A2(new_n462), .A3(new_n448), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n478), .A2(G469), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n473), .A2(new_n475), .A3(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(G221), .ZN(new_n482));
  XOR2_X1   g296(.A(KEYINPUT9), .B(G234), .Z(new_n483));
  AOI21_X1  g297(.A(new_n482), .B1(new_n483), .B2(new_n233), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n481), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT20), .ZN(new_n487));
  NOR2_X1   g301(.A1(G475), .A2(G902), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(KEYINPUT84), .ZN(new_n489));
  INV_X1    g303(.A(G237), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n490), .A2(new_n223), .A3(G214), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n261), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n307), .A2(G143), .A3(G214), .ZN(new_n493));
  NAND2_X1  g307(.A1(KEYINPUT18), .A2(G131), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n492), .A2(new_n493), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(KEYINPUT18), .A3(G131), .ZN(new_n497));
  XOR2_X1   g311(.A(G125), .B(G140), .Z(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G146), .ZN(new_n499));
  AND3_X1   g313(.A1(new_n499), .A2(KEYINPUT81), .A3(new_n219), .ZN(new_n500));
  AOI21_X1  g314(.A(KEYINPUT81), .B1(new_n499), .B2(new_n219), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n495), .B(new_n497), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n496), .A2(G131), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n492), .A2(new_n257), .A3(new_n493), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n498), .A2(KEYINPUT19), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT19), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n187), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n506), .A2(new_n218), .A3(new_n508), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n505), .A2(new_n214), .A3(new_n215), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n502), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT82), .ZN(new_n512));
  XNOR2_X1  g326(.A(G113), .B(G122), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(new_n386), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT82), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n502), .A2(new_n510), .A3(new_n516), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n512), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n195), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n496), .A2(KEYINPUT17), .A3(G131), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n519), .B(new_n520), .C1(KEYINPUT17), .C2(new_n505), .ZN(new_n521));
  XOR2_X1   g335(.A(new_n514), .B(KEYINPUT83), .Z(new_n522));
  AND3_X1   g336(.A1(new_n521), .A2(new_n502), .A3(new_n522), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n487), .B(new_n489), .C1(new_n518), .C2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT85), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n514), .B1(new_n511), .B2(KEYINPUT82), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n523), .B1(new_n517), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n488), .ZN(new_n529));
  OAI21_X1  g343(.A(KEYINPUT20), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n523), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n527), .A2(new_n517), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n533), .A2(KEYINPUT85), .A3(new_n487), .A4(new_n489), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n526), .A2(new_n530), .A3(new_n534), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n521), .A2(new_n502), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n536), .A2(new_n514), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n233), .B1(new_n537), .B2(new_n523), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(G475), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT13), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n542), .B1(new_n196), .B2(G143), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT86), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n196), .A2(G143), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n261), .A2(G128), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT86), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n547), .A3(new_n542), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n544), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT87), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n196), .A2(G143), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT13), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n544), .A2(new_n548), .A3(KEYINPUT87), .A4(new_n545), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n551), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(G134), .ZN(new_n556));
  XNOR2_X1  g370(.A(G116), .B(G122), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(new_n389), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT89), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT88), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n261), .A2(G128), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n560), .B1(new_n552), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n546), .A2(new_n545), .A3(KEYINPUT88), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n559), .B1(new_n564), .B2(new_n245), .ZN(new_n565));
  AOI211_X1 g379(.A(KEYINPUT89), .B(G134), .C1(new_n562), .C2(new_n563), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n556), .A2(new_n558), .A3(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n564), .B(new_n245), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT14), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n557), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(G116), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n572), .A2(KEYINPUT14), .A3(G122), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n571), .A2(G107), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT90), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n571), .A2(KEYINPUT90), .A3(G107), .A4(new_n573), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n557), .A2(new_n389), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n569), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n568), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n483), .A2(G217), .A3(new_n223), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n582), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n568), .A2(new_n584), .A3(new_n580), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n233), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT15), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n587), .A2(new_n588), .A3(G478), .ZN(new_n589));
  INV_X1    g403(.A(G478), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n586), .B(new_n233), .C1(KEYINPUT15), .C2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n541), .A2(new_n593), .ZN(new_n594));
  NOR3_X1   g408(.A1(new_n444), .A2(new_n486), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n365), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(G101), .ZN(G3));
  INV_X1    g411(.A(new_n337), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT91), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n599), .B(new_n233), .C1(new_n317), .C2(new_n336), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n600), .A2(G472), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n599), .B1(new_n345), .B2(new_n233), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n598), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n241), .ZN(new_n605));
  AND2_X1   g419(.A1(new_n481), .A2(new_n485), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n604), .A2(KEYINPUT92), .A3(new_n605), .A4(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT92), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n600), .A2(G472), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n606), .B(new_n337), .C1(new_n609), .C2(new_n602), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n608), .B1(new_n610), .B2(new_n241), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n585), .A2(KEYINPUT93), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT93), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n568), .A2(new_n614), .A3(new_n580), .A4(new_n584), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n613), .A2(new_n583), .A3(KEYINPUT33), .A4(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT94), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n615), .A2(KEYINPUT33), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n619), .A2(KEYINPUT94), .A3(new_n583), .A4(new_n613), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT33), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n586), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n621), .A2(G478), .A3(new_n233), .A4(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT95), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n587), .A2(new_n590), .ZN(new_n627));
  AOI22_X1  g441(.A1(new_n618), .A2(new_n620), .B1(new_n622), .B2(new_n586), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n628), .A2(KEYINPUT95), .A3(G478), .A4(new_n233), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n626), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n540), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n631), .A2(new_n444), .A3(KEYINPUT96), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT96), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n630), .A2(new_n540), .ZN(new_n634));
  INV_X1    g448(.A(new_n444), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n612), .B1(new_n632), .B2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT34), .B(G104), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G6));
  INV_X1    g453(.A(KEYINPUT97), .ZN(new_n640));
  OAI221_X1 g454(.A(new_n377), .B1(new_n640), .B2(new_n375), .C1(new_n441), .C2(new_n443), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n533), .A2(new_n487), .A3(new_n488), .ZN(new_n642));
  AOI22_X1  g456(.A1(new_n530), .A2(new_n642), .B1(G475), .B2(new_n538), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n592), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n375), .A2(new_n640), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n641), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n612), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G107), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT98), .B(KEYINPUT35), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G9));
  NOR2_X1   g465(.A1(new_n226), .A2(KEYINPUT36), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n221), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n237), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n236), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n444), .A2(new_n594), .A3(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n610), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(new_n659), .B(G110), .Z(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT99), .B(KEYINPUT37), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G12));
  NAND2_X1  g476(.A1(new_n350), .A2(new_n364), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n441), .A2(new_n443), .ZN(new_n664));
  INV_X1    g478(.A(new_n377), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n664), .A2(new_n665), .A3(new_n656), .ZN(new_n666));
  INV_X1    g480(.A(G900), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n370), .B1(new_n374), .B2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n644), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n663), .A2(new_n606), .A3(new_n666), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G128), .ZN(G30));
  AOI22_X1  g485(.A1(new_n535), .A2(new_n539), .B1(new_n589), .B2(new_n591), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n668), .B(KEYINPUT39), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n486), .A2(new_n674), .ZN(new_n675));
  OR2_X1    g489(.A1(new_n675), .A2(KEYINPUT40), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(KEYINPUT40), .ZN(new_n677));
  AOI211_X1 g491(.A(new_n665), .B(new_n673), .C1(new_n676), .C2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n353), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n679), .A2(new_n354), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n306), .A2(new_n358), .A3(new_n354), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n233), .ZN(new_n682));
  OAI21_X1  g496(.A(G472), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n350), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n427), .B1(new_n426), .B2(new_n384), .ZN(new_n685));
  AOI211_X1 g499(.A(KEYINPUT80), .B(new_n383), .C1(new_n424), .C2(new_n425), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n440), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n442), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n429), .A2(new_n378), .A3(new_n440), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT38), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n678), .A2(new_n656), .A3(new_n684), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G143), .ZN(G45));
  INV_X1    g507(.A(new_n668), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n630), .A2(new_n540), .A3(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n663), .A2(new_n695), .A3(new_n666), .A4(new_n606), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G146), .ZN(G48));
  INV_X1    g511(.A(G472), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n698), .B1(new_n356), .B2(new_n362), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n699), .B1(new_n347), .B2(new_n349), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n233), .B1(new_n463), .B2(new_n472), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(G469), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n702), .A2(new_n485), .A3(new_n473), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n700), .A2(new_n241), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n705), .B1(new_n636), .B2(new_n632), .ZN(new_n706));
  XNOR2_X1  g520(.A(KEYINPUT41), .B(G113), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G15));
  NAND2_X1  g522(.A1(new_n705), .A2(new_n647), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT100), .B(G116), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G18));
  OAI211_X1 g525(.A(new_n703), .B(new_n377), .C1(new_n441), .C2(new_n443), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT101), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n690), .A2(KEYINPUT101), .A3(new_n377), .A4(new_n703), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n594), .A2(new_n656), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n716), .A2(new_n663), .A3(new_n376), .A4(new_n717), .ZN(new_n718));
  XOR2_X1   g532(.A(KEYINPUT102), .B(G119), .Z(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G21));
  NOR2_X1   g534(.A1(new_n641), .A2(new_n646), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT103), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n722), .B1(new_n359), .B2(new_n334), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n354), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n359), .A2(new_n334), .A3(new_n722), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n244), .B1(new_n726), .B2(new_n317), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT104), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n345), .A2(new_n233), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(G472), .ZN(new_n731));
  OAI211_X1 g545(.A(KEYINPUT104), .B(new_n244), .C1(new_n726), .C2(new_n317), .ZN(new_n732));
  AND4_X1   g546(.A1(new_n605), .A2(new_n729), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n721), .A2(new_n672), .A3(new_n703), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G122), .ZN(G24));
  NAND3_X1  g549(.A1(new_n630), .A2(new_n540), .A3(new_n694), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n729), .A2(new_n731), .A3(new_n655), .A4(new_n732), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n716), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G125), .ZN(G27));
  INV_X1    g554(.A(KEYINPUT105), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n688), .A2(new_n377), .A3(new_n689), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n741), .B1(new_n742), .B2(new_n486), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n664), .A2(KEYINPUT105), .A3(new_n606), .A4(new_n377), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(new_n365), .A3(new_n695), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT42), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n736), .B1(new_n743), .B2(new_n744), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n364), .A2(new_n339), .A3(new_n346), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n605), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n750), .A2(new_n747), .ZN(new_n751));
  AOI22_X1  g565(.A1(new_n746), .A2(new_n747), .B1(new_n748), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(new_n257), .ZN(G33));
  NAND3_X1  g567(.A1(new_n745), .A2(new_n365), .A3(new_n669), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G134), .ZN(G36));
  NAND2_X1  g569(.A1(new_n630), .A2(new_n541), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT43), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n756), .B(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n604), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(new_n759), .A3(new_n655), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT107), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(new_n762), .A3(KEYINPUT44), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT44), .ZN(new_n764));
  OAI21_X1  g578(.A(KEYINPUT107), .B1(new_n760), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n742), .B1(new_n760), .B2(new_n764), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n478), .A2(new_n479), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(KEYINPUT45), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(G469), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT106), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n769), .A2(KEYINPUT106), .A3(G469), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n474), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n774), .A2(KEYINPUT46), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n473), .B1(new_n774), .B2(KEYINPUT46), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n485), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n777), .A2(new_n674), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n766), .A2(new_n767), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G137), .ZN(G39));
  INV_X1    g595(.A(KEYINPUT47), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n777), .A2(new_n782), .ZN(new_n783));
  OAI211_X1 g597(.A(KEYINPUT47), .B(new_n485), .C1(new_n775), .C2(new_n776), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n441), .A2(new_n443), .A3(new_n665), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n663), .A2(new_n605), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n785), .A2(new_n695), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G140), .ZN(G42));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n672), .B(new_n377), .C1(new_n441), .C2(new_n443), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n486), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n684), .A2(new_n792), .A3(new_n656), .A4(new_n694), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n670), .A2(new_n739), .A3(new_n696), .A4(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n700), .A2(new_n486), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n797), .B(new_n666), .C1(new_n669), .C2(new_n695), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n798), .A2(KEYINPUT52), .A3(new_n739), .A4(new_n793), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT53), .B1(new_n800), .B2(KEYINPUT109), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n706), .A2(new_n709), .A3(new_n718), .A4(new_n734), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n365), .A2(new_n595), .B1(new_n657), .B2(new_n658), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n541), .A2(new_n592), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n631), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n607), .A2(new_n611), .A3(new_n721), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n802), .A2(new_n807), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n700), .A2(new_n486), .A3(new_n656), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n592), .A2(new_n668), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n786), .A2(KEYINPUT108), .A3(new_n643), .A4(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT108), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n688), .A2(new_n377), .A3(new_n689), .A4(new_n643), .ZN(new_n813));
  INV_X1    g627(.A(new_n810), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n809), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n737), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n745), .A2(new_n695), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n817), .A2(new_n754), .A3(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n752), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n800), .A2(new_n808), .A3(new_n821), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n801), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n801), .A2(new_n822), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n790), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n826));
  INV_X1    g640(.A(new_n807), .ZN(new_n827));
  AND4_X1   g641(.A1(new_n706), .A2(new_n709), .A3(new_n718), .A4(new_n734), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n821), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n796), .A2(new_n799), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n826), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n800), .A2(new_n808), .A3(KEYINPUT53), .A4(new_n821), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n831), .A2(new_n790), .A3(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(KEYINPUT110), .B1(new_n825), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n758), .A2(new_n370), .A3(new_n733), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(new_n716), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n758), .A2(new_n370), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n691), .A2(new_n377), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n839), .A2(new_n703), .A3(new_n733), .A4(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT50), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n837), .A2(KEYINPUT50), .A3(new_n703), .A4(new_n840), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n702), .A2(new_n473), .ZN(new_n846));
  XOR2_X1   g660(.A(new_n846), .B(KEYINPUT111), .Z(new_n847));
  AND2_X1   g661(.A1(new_n847), .A2(new_n484), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n786), .B(new_n837), .C1(new_n785), .C2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n742), .A2(new_n704), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n241), .A2(new_n369), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n850), .A2(new_n350), .A3(new_n683), .A4(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT112), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n852), .A2(new_n853), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n854), .A2(new_n855), .A3(new_n630), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n541), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n839), .A2(new_n818), .A3(new_n850), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n845), .A2(new_n849), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT51), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI22_X1  g675(.A1(new_n843), .A2(new_n844), .B1(new_n856), .B2(new_n541), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n862), .A2(KEYINPUT51), .A3(new_n858), .A4(new_n849), .ZN(new_n863));
  INV_X1    g677(.A(new_n750), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n839), .A2(new_n864), .A3(new_n850), .ZN(new_n865));
  XNOR2_X1  g679(.A(KEYINPUT113), .B(KEYINPUT48), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  OR2_X1    g681(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n865), .A2(new_n867), .ZN(new_n869));
  OR3_X1    g683(.A1(new_n854), .A2(new_n855), .A3(new_n631), .ZN(new_n870));
  AND4_X1   g684(.A1(new_n367), .A2(new_n868), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  AND4_X1   g685(.A1(new_n838), .A2(new_n861), .A3(new_n863), .A4(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT110), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n801), .A2(new_n822), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n801), .A2(new_n822), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n873), .B(new_n833), .C1(new_n876), .C2(new_n790), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n835), .A2(new_n872), .A3(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT114), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n366), .A2(new_n223), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n835), .A2(new_n872), .A3(new_n877), .A4(KEYINPUT114), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n846), .B(KEYINPUT49), .Z(new_n884));
  NOR3_X1   g698(.A1(new_n691), .A2(new_n884), .A3(new_n241), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n684), .A2(new_n484), .A3(new_n756), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n885), .A2(new_n377), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n883), .A2(new_n887), .ZN(G75));
  XNOR2_X1  g702(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  NOR4_X1   g704(.A1(new_n802), .A2(new_n752), .A3(new_n820), .A4(new_n807), .ZN(new_n891));
  AOI21_X1  g705(.A(KEYINPUT53), .B1(new_n891), .B2(new_n800), .ZN(new_n892));
  AND4_X1   g706(.A1(KEYINPUT53), .A2(new_n800), .A3(new_n808), .A4(new_n821), .ZN(new_n893));
  OAI211_X1 g707(.A(G210), .B(G902), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT56), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n426), .B(new_n383), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n896), .B1(new_n894), .B2(new_n895), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n890), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n896), .ZN(new_n900));
  INV_X1    g714(.A(G210), .ZN(new_n901));
  AOI211_X1 g715(.A(new_n901), .B(new_n233), .C1(new_n831), .C2(new_n832), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n900), .B1(new_n902), .B2(KEYINPUT56), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n903), .A2(new_n889), .A3(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n223), .A2(G952), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n899), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(KEYINPUT116), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT116), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n899), .A2(new_n905), .A3(new_n910), .A4(new_n907), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n909), .A2(new_n911), .ZN(G51));
  NAND2_X1  g726(.A1(new_n831), .A2(new_n832), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(KEYINPUT54), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n833), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n474), .B(KEYINPUT57), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n917), .B1(new_n463), .B2(new_n472), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n233), .B1(new_n831), .B2(new_n832), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n919), .A2(new_n772), .A3(new_n773), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n906), .B1(new_n918), .B2(new_n920), .ZN(G54));
  NAND2_X1  g735(.A1(KEYINPUT58), .A2(G475), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT117), .ZN(new_n923));
  OR2_X1    g737(.A1(new_n922), .A2(KEYINPUT117), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n919), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n925), .A2(new_n528), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n925), .A2(new_n528), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n926), .A2(new_n927), .A3(new_n906), .ZN(G60));
  XNOR2_X1  g742(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n590), .A2(new_n233), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n929), .B(new_n930), .Z(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n915), .A2(new_n628), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n931), .B1(new_n835), .B2(new_n877), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n907), .B(new_n933), .C1(new_n934), .C2(new_n628), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(G63));
  NAND2_X1  g750(.A1(G217), .A2(G902), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT60), .Z(new_n938));
  NAND2_X1  g752(.A1(new_n913), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(KEYINPUT119), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT119), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n913), .A2(new_n941), .A3(new_n938), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n653), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n940), .A2(new_n230), .A3(new_n942), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n944), .A2(new_n945), .A3(new_n907), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT61), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n944), .A2(new_n945), .A3(KEYINPUT61), .A4(new_n907), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(G66));
  INV_X1    g764(.A(new_n808), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT120), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n223), .B1(new_n371), .B2(G224), .ZN(new_n953));
  AOI22_X1  g767(.A1(new_n951), .A2(new_n223), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n954), .B1(new_n952), .B2(new_n953), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n424), .B(new_n425), .C1(G898), .C2(new_n223), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(G69));
  INV_X1    g771(.A(KEYINPUT124), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n292), .A2(new_n298), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n506), .A2(new_n508), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n959), .B(new_n960), .Z(new_n961));
  INV_X1    g775(.A(KEYINPUT123), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n739), .A2(new_n696), .A3(new_n670), .ZN(new_n963));
  NAND2_X1  g777(.A1(KEYINPUT121), .A2(KEYINPUT62), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n692), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(KEYINPUT121), .A2(KEYINPUT62), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n780), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n965), .B1(KEYINPUT121), .B2(KEYINPUT62), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n365), .A2(new_n675), .A3(new_n786), .A4(new_n805), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT122), .Z(new_n972));
  NAND3_X1  g786(.A1(new_n788), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n962), .B1(new_n969), .B2(new_n973), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n788), .A2(new_n970), .A3(new_n972), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n778), .B1(new_n763), .B2(new_n765), .ZN(new_n976));
  AOI22_X1  g790(.A1(new_n976), .A2(new_n767), .B1(new_n967), .B2(new_n966), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n975), .A2(new_n977), .A3(KEYINPUT123), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n974), .A2(new_n978), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n958), .B(new_n961), .C1(new_n979), .C2(G953), .ZN(new_n980));
  AOI21_X1  g794(.A(G953), .B1(new_n974), .B2(new_n978), .ZN(new_n981));
  INV_X1    g795(.A(new_n961), .ZN(new_n982));
  OAI21_X1  g796(.A(KEYINPUT124), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(G900), .A2(G953), .ZN(new_n984));
  INV_X1    g798(.A(new_n752), .ZN(new_n985));
  OR3_X1    g799(.A1(new_n778), .A2(new_n750), .A3(new_n791), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n986), .A2(new_n754), .A3(new_n788), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n780), .A2(KEYINPUT125), .A3(new_n963), .ZN(new_n988));
  AOI21_X1  g802(.A(KEYINPUT125), .B1(new_n780), .B2(new_n963), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n985), .B(new_n987), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n984), .B(new_n982), .C1(new_n990), .C2(G953), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n980), .A2(new_n983), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n223), .B1(G227), .B2(G900), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n993), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n980), .A2(new_n983), .A3(new_n995), .A4(new_n991), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n994), .A2(new_n996), .ZN(G72));
  NAND2_X1  g811(.A1(G472), .A2(G902), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT63), .Z(new_n999));
  OAI21_X1  g813(.A(new_n999), .B1(new_n990), .B2(new_n951), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n1000), .A2(new_n354), .A3(new_n679), .ZN(new_n1001));
  INV_X1    g815(.A(new_n999), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n876), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT127), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n313), .A2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(new_n355), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n906), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1001), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n974), .A2(new_n978), .A3(new_n808), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT126), .ZN(new_n1010));
  AND3_X1   g824(.A1(new_n1009), .A2(new_n1010), .A3(new_n999), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1010), .B1(new_n1009), .B2(new_n999), .ZN(new_n1012));
  INV_X1    g826(.A(new_n680), .ZN(new_n1013));
  NOR3_X1   g827(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n1008), .A2(new_n1014), .ZN(G57));
endmodule


