//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 1 0 1 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 1 1 1 1 1 0 0 1 1 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  XOR2_X1   g002(.A(G110), .B(G140), .Z(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT73), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(KEYINPUT74), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  AND2_X1   g006(.A1(new_n192), .A2(G227), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n191), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G137), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G134), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(G134), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n199));
  AND2_X1   g013(.A1(new_n199), .A2(KEYINPUT11), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n196), .B1(new_n198), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G131), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(KEYINPUT11), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n199), .A2(KEYINPUT11), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(new_n197), .ZN(new_n205));
  AND3_X1   g019(.A1(new_n201), .A2(new_n202), .A3(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n202), .B1(new_n201), .B2(new_n205), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT76), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G143), .ZN(new_n212));
  INV_X1    g026(.A(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G146), .ZN(new_n214));
  AOI21_X1  g028(.A(G128), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n213), .A2(KEYINPUT1), .A3(G146), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT66), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n219));
  XNOR2_X1  g033(.A(G143), .B(G146), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n219), .B(new_n216), .C1(new_n220), .C2(G128), .ZN(new_n221));
  INV_X1    g035(.A(G128), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n223), .A2(new_n212), .A3(new_n214), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n218), .A2(new_n221), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT10), .ZN(new_n227));
  INV_X1    g041(.A(G104), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT3), .B1(new_n228), .B2(G107), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n230));
  INV_X1    g044(.A(G107), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n230), .A2(new_n231), .A3(G104), .ZN(new_n232));
  INV_X1    g046(.A(G101), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n228), .A2(G107), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n229), .A2(new_n232), .A3(new_n233), .A4(new_n234), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n231), .A2(G104), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n228), .A2(G107), .ZN(new_n237));
  OAI21_X1  g051(.A(G101), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n235), .A2(new_n238), .A3(KEYINPUT75), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT75), .B1(new_n235), .B2(new_n238), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n210), .B1(new_n227), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n235), .A2(new_n238), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT75), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n235), .A2(new_n238), .A3(KEYINPUT75), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n247), .A2(KEYINPUT76), .A3(KEYINPUT10), .A4(new_n226), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n242), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT10), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n216), .B1(new_n220), .B2(G128), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n251), .A2(new_n224), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n250), .B1(new_n252), .B2(new_n243), .ZN(new_n253));
  AND2_X1   g067(.A1(KEYINPUT0), .A2(G128), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n220), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(KEYINPUT0), .A2(G128), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n256), .B1(new_n220), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n229), .A2(new_n232), .A3(new_n234), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n261), .A3(G101), .ZN(new_n262));
  AND2_X1   g076(.A1(new_n260), .A2(G101), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n235), .A2(KEYINPUT4), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n259), .B(new_n262), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n253), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(KEYINPUT78), .B1(new_n249), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT78), .ZN(new_n269));
  AOI211_X1 g083(.A(new_n269), .B(new_n266), .C1(new_n242), .C2(new_n248), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n209), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n249), .A2(new_n208), .A3(new_n267), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n194), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT77), .ZN(new_n274));
  INV_X1    g088(.A(new_n243), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n274), .B1(new_n226), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n275), .B1(new_n251), .B2(new_n224), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n224), .B1(new_n251), .B2(KEYINPUT66), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n278), .A2(KEYINPUT77), .A3(new_n221), .A4(new_n243), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n276), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n280), .A2(KEYINPUT12), .A3(new_n209), .ZN(new_n281));
  AOI21_X1  g095(.A(KEYINPUT12), .B1(new_n280), .B2(new_n209), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n194), .B(new_n272), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n187), .B(new_n188), .C1(new_n273), .C2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n272), .B1(new_n281), .B2(new_n282), .ZN(new_n286));
  INV_X1    g100(.A(new_n194), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NOR3_X1   g102(.A1(new_n227), .A2(new_n241), .A3(new_n210), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n250), .B1(new_n278), .B2(new_n221), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT76), .B1(new_n290), .B2(new_n247), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n267), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n269), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n249), .A2(KEYINPUT78), .A3(new_n267), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n208), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n194), .A2(new_n272), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n288), .B(G469), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n187), .A2(new_n188), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n285), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT9), .B(G234), .ZN(new_n301));
  OAI21_X1  g115(.A(G221), .B1(new_n301), .B2(G902), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(G214), .B1(G237), .B2(G902), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT20), .ZN(new_n306));
  NOR2_X1   g120(.A1(G475), .A2(G902), .ZN(new_n307));
  NOR2_X1   g121(.A1(G237), .A2(G953), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(G143), .A3(G214), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(G143), .B1(new_n308), .B2(G214), .ZN(new_n311));
  OAI21_X1  g125(.A(G131), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT17), .ZN(new_n313));
  INV_X1    g127(.A(G237), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n314), .A2(new_n192), .A3(G214), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n213), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(new_n202), .A3(new_n309), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n312), .A2(new_n313), .A3(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT16), .ZN(new_n319));
  INV_X1    g133(.A(G125), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G140), .ZN(new_n321));
  INV_X1    g135(.A(G140), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G125), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT71), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n321), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n320), .A2(KEYINPUT71), .A3(G140), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n319), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n323), .A2(KEYINPUT16), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n211), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n328), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n320), .A2(KEYINPUT71), .A3(G140), .ZN(new_n331));
  XNOR2_X1  g145(.A(G125), .B(G140), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n331), .B1(new_n332), .B2(new_n324), .ZN(new_n333));
  OAI211_X1 g147(.A(G146), .B(new_n330), .C1(new_n333), .C2(new_n319), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n316), .A2(new_n309), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(KEYINPUT17), .A3(G131), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n318), .A2(new_n329), .A3(new_n334), .A4(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT83), .ZN(new_n338));
  OAI211_X1 g152(.A(KEYINPUT18), .B(G131), .C1(new_n335), .C2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n332), .A2(new_n211), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n325), .A2(new_n326), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n340), .B1(new_n341), .B2(new_n211), .ZN(new_n342));
  NAND2_X1  g156(.A1(KEYINPUT18), .A2(G131), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n316), .A2(KEYINPUT83), .A3(new_n343), .A4(new_n309), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n339), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(G113), .B(G122), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(new_n228), .ZN(new_n347));
  AND3_X1   g161(.A1(new_n337), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n312), .A2(new_n317), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT19), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n332), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n351), .B1(new_n341), .B2(new_n350), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n334), .B(new_n349), .C1(new_n352), .C2(G146), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n347), .B1(new_n353), .B2(new_n345), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n306), .B(new_n307), .C1(new_n348), .C2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT84), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n337), .A2(new_n345), .A3(new_n347), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n353), .A2(new_n345), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n357), .B1(new_n358), .B2(new_n347), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT84), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n359), .A2(new_n360), .A3(new_n306), .A4(new_n307), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n307), .B1(new_n348), .B2(new_n354), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(KEYINPUT20), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n356), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n337), .A2(new_n345), .ZN(new_n365));
  INV_X1    g179(.A(new_n347), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT85), .ZN(new_n367));
  OR2_X1    g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n365), .A2(new_n367), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n188), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G475), .ZN(new_n371));
  AND3_X1   g185(.A1(new_n364), .A2(KEYINPUT86), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(KEYINPUT86), .B1(new_n364), .B2(new_n371), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(G210), .B1(G237), .B2(G902), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n375), .B(KEYINPUT82), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT81), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  XOR2_X1   g192(.A(KEYINPUT2), .B(G113), .Z(new_n379));
  OR2_X1    g193(.A1(KEYINPUT67), .A2(G116), .ZN(new_n380));
  NAND2_X1  g194(.A1(KEYINPUT67), .A2(G116), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(G119), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G116), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n379), .B(new_n382), .C1(new_n383), .C2(G119), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT2), .B(G113), .ZN(new_n385));
  AND2_X1   g199(.A1(KEYINPUT67), .A2(G116), .ZN(new_n386));
  NOR2_X1   g200(.A1(KEYINPUT67), .A2(G116), .ZN(new_n387));
  INV_X1    g201(.A(G119), .ZN(new_n388));
  NOR3_X1   g202(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n383), .A2(G119), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n385), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n384), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n260), .A2(G101), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(KEYINPUT4), .A3(new_n235), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n392), .A2(new_n394), .A3(new_n262), .ZN(new_n395));
  XNOR2_X1  g209(.A(G110), .B(G122), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n382), .B(KEYINPUT5), .C1(new_n383), .C2(G119), .ZN(new_n397));
  INV_X1    g211(.A(G113), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT5), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n398), .B1(new_n390), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n384), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n395), .B(new_n396), .C1(new_n241), .C2(new_n402), .ZN(new_n403));
  AOI22_X1  g217(.A1(new_n261), .A2(new_n263), .B1(new_n384), .B2(new_n391), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n389), .A2(new_n390), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n397), .A2(new_n400), .B1(new_n405), .B2(new_n379), .ZN(new_n406));
  AOI22_X1  g220(.A1(new_n404), .A2(new_n394), .B1(new_n247), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n396), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT79), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n403), .B(KEYINPUT6), .C1(new_n407), .C2(new_n409), .ZN(new_n410));
  OR2_X1    g224(.A1(new_n258), .A2(new_n220), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n320), .B1(new_n411), .B2(new_n256), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n412), .B1(new_n226), .B2(new_n320), .ZN(new_n413));
  INV_X1    g227(.A(G224), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(G953), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n413), .B(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n395), .B1(new_n241), .B2(new_n402), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT6), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n417), .A2(KEYINPUT79), .A3(new_n418), .A4(new_n408), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n410), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT7), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n421), .A2(KEYINPUT80), .ZN(new_n422));
  AOI21_X1  g236(.A(G125), .B1(new_n278), .B2(new_n221), .ZN(new_n423));
  OAI221_X1 g237(.A(new_n422), .B1(new_n414), .B2(G953), .C1(new_n423), .C2(new_n412), .ZN(new_n424));
  AND2_X1   g238(.A1(KEYINPUT80), .A2(KEYINPUT7), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n415), .B1(new_n413), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n396), .B(KEYINPUT8), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n401), .A2(new_n384), .A3(new_n275), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n275), .B1(new_n401), .B2(new_n384), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n413), .A2(new_n421), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(new_n403), .A3(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n188), .B1(new_n427), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n378), .B1(new_n420), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n402), .A2(new_n243), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n406), .A2(new_n275), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n438), .A2(new_n428), .B1(new_n421), .B2(new_n413), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n439), .A2(new_n403), .A3(new_n426), .A4(new_n424), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n410), .A2(new_n416), .A3(new_n419), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n440), .A2(new_n441), .A3(new_n188), .A4(new_n377), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n435), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G478), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n444), .A2(KEYINPUT15), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(G128), .B(G143), .ZN(new_n447));
  INV_X1    g261(.A(G134), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n447), .B(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(KEYINPUT87), .B1(new_n383), .B2(G122), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT87), .ZN(new_n451));
  INV_X1    g265(.A(G122), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n452), .A3(G116), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n380), .A2(G122), .A3(new_n381), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(new_n455), .A3(new_n231), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n449), .A2(new_n456), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n455), .A2(KEYINPUT14), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n454), .B1(new_n455), .B2(KEYINPUT14), .ZN(new_n459));
  OAI21_X1  g273(.A(G107), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n454), .A2(new_n455), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G107), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n456), .ZN(new_n463));
  AOI21_X1  g277(.A(KEYINPUT13), .B1(new_n222), .B2(G143), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(new_n448), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n465), .B(new_n447), .ZN(new_n466));
  AOI22_X1  g280(.A1(new_n457), .A2(new_n460), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(G217), .ZN(new_n469));
  NOR3_X1   g283(.A1(new_n301), .A2(new_n469), .A3(G953), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n468), .A2(KEYINPUT88), .A3(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT88), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n473), .B1(new_n467), .B2(new_n470), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n467), .A2(new_n470), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n472), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n446), .B1(new_n476), .B2(new_n188), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n476), .A2(new_n188), .A3(new_n446), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(G234), .A2(G237), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n481), .A2(G952), .A3(new_n192), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n481), .A2(G902), .A3(G953), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT21), .B(G898), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n480), .A2(new_n485), .ZN(new_n486));
  AND4_X1   g300(.A1(new_n305), .A2(new_n374), .A3(new_n443), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n304), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(KEYINPUT23), .B1(new_n222), .B2(G119), .ZN(new_n489));
  AOI21_X1  g303(.A(KEYINPUT70), .B1(new_n222), .B2(G119), .ZN(new_n490));
  XOR2_X1   g304(.A(new_n489), .B(new_n490), .Z(new_n491));
  INV_X1    g305(.A(G110), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OR3_X1    g307(.A1(new_n222), .A2(KEYINPUT69), .A3(G119), .ZN(new_n494));
  OAI21_X1  g308(.A(KEYINPUT69), .B1(new_n222), .B2(G119), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n494), .B(new_n495), .C1(new_n388), .C2(G128), .ZN(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT24), .B(G110), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n334), .B(new_n340), .C1(new_n493), .C2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n329), .A2(new_n334), .ZN(new_n500));
  OR2_X1    g314(.A1(new_n496), .A2(new_n497), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n500), .B(new_n501), .C1(new_n492), .C2(new_n491), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n192), .A2(G221), .A3(G234), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(KEYINPUT72), .ZN(new_n505));
  XOR2_X1   g319(.A(KEYINPUT22), .B(G137), .Z(new_n506));
  XNOR2_X1  g320(.A(new_n505), .B(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n505), .ZN(new_n509));
  AND2_X1   g323(.A1(new_n509), .A2(new_n506), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n509), .A2(new_n506), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n502), .B(new_n499), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n508), .A2(new_n188), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT25), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT25), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n508), .A2(new_n515), .A3(new_n188), .A4(new_n512), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n469), .B1(G234), .B2(new_n188), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AND2_X1   g332(.A1(new_n508), .A2(new_n512), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n517), .A2(G902), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n201), .A2(new_n202), .A3(new_n205), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n196), .A2(KEYINPUT65), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n448), .A2(KEYINPUT65), .A3(G137), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n197), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G131), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n226), .A2(new_n523), .A3(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n259), .B1(new_n206), .B2(new_n207), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT30), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n530), .B1(new_n528), .B2(new_n529), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n392), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n528), .A2(new_n529), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n534), .A2(new_n392), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n308), .A2(G210), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(KEYINPUT27), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT26), .B(G101), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n538), .B(new_n539), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n533), .A2(KEYINPUT31), .A3(new_n536), .A4(new_n540), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n541), .A2(new_n188), .ZN(new_n542));
  INV_X1    g356(.A(G472), .ZN(new_n543));
  INV_X1    g357(.A(new_n392), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT68), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n528), .A2(new_n529), .A3(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n545), .B1(new_n528), .B2(new_n529), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n544), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT28), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n544), .B1(new_n528), .B2(new_n529), .ZN(new_n552));
  OAI21_X1  g366(.A(KEYINPUT28), .B1(new_n535), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n540), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n533), .A2(new_n540), .A3(new_n536), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT31), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n542), .B(new_n543), .C1(new_n554), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT32), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n541), .A2(new_n188), .ZN(new_n560));
  INV_X1    g374(.A(new_n548), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n392), .B1(new_n561), .B2(new_n546), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n553), .B1(new_n562), .B2(KEYINPUT28), .ZN(new_n563));
  INV_X1    g377(.A(new_n540), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n534), .A2(KEYINPUT30), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n535), .B1(new_n568), .B2(new_n392), .ZN(new_n569));
  AOI21_X1  g383(.A(KEYINPUT31), .B1(new_n569), .B2(new_n540), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n560), .B1(new_n565), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT32), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n571), .A2(new_n572), .A3(new_n543), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n559), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n533), .A2(new_n536), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n564), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT29), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n576), .B(new_n577), .C1(new_n563), .C2(new_n564), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n551), .A2(KEYINPUT29), .A3(new_n540), .A4(new_n553), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n578), .A2(new_n188), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(G472), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n522), .B1(new_n574), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n488), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(new_n233), .ZN(G3));
  OAI21_X1  g399(.A(new_n542), .B1(new_n554), .B2(new_n557), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n586), .A2(KEYINPUT89), .A3(G472), .ZN(new_n587));
  NAND2_X1  g401(.A1(KEYINPUT89), .A2(G472), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n571), .A2(new_n588), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NOR3_X1   g405(.A1(new_n591), .A2(new_n303), .A3(new_n522), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n470), .A2(KEYINPUT90), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n468), .A2(new_n593), .ZN(new_n594));
  NOR3_X1   g408(.A1(new_n467), .A2(KEYINPUT90), .A3(new_n470), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT33), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n596), .B1(new_n476), .B2(KEYINPUT33), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n597), .A2(G478), .A3(new_n188), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n476), .A2(new_n188), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n444), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n601), .B1(new_n372), .B2(new_n373), .ZN(new_n602));
  INV_X1    g416(.A(new_n305), .ZN(new_n603));
  INV_X1    g417(.A(new_n434), .ZN(new_n604));
  INV_X1    g418(.A(new_n376), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n604), .A2(new_n441), .A3(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n376), .B1(new_n420), .B2(new_n434), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n603), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n485), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n602), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n592), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT34), .B(G104), .Z(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G6));
  INV_X1    g428(.A(new_n479), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n615), .A2(new_n477), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n363), .A2(new_n355), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n371), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n610), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n592), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT35), .B(G107), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G9));
  INV_X1    g436(.A(KEYINPUT92), .ZN(new_n623));
  OAI21_X1  g437(.A(KEYINPUT91), .B1(new_n507), .B2(KEYINPUT36), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT91), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT36), .ZN(new_n626));
  OAI211_X1 g440(.A(new_n625), .B(new_n626), .C1(new_n510), .C2(new_n511), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n503), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n499), .A2(new_n502), .A3(new_n624), .A4(new_n627), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n623), .B1(new_n631), .B2(new_n520), .ZN(new_n632));
  INV_X1    g446(.A(new_n520), .ZN(new_n633));
  AOI211_X1 g447(.A(KEYINPUT92), .B(new_n633), .C1(new_n629), .C2(new_n630), .ZN(new_n634));
  OR2_X1    g448(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT93), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n635), .A2(new_n636), .A3(new_n518), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n513), .A2(KEYINPUT25), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n516), .A2(new_n517), .ZN(new_n639));
  OAI22_X1  g453(.A1(new_n638), .A2(new_n639), .B1(new_n632), .B2(new_n634), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(KEYINPUT93), .ZN(new_n641));
  AND4_X1   g455(.A1(new_n587), .A2(new_n637), .A3(new_n641), .A4(new_n589), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n304), .A2(new_n487), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT37), .B(G110), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G12));
  AOI22_X1  g459(.A1(new_n559), .A2(new_n573), .B1(new_n580), .B2(G472), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n637), .A2(new_n641), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n608), .ZN(new_n649));
  INV_X1    g463(.A(new_n618), .ZN(new_n650));
  XNOR2_X1  g464(.A(KEYINPUT94), .B(G900), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n482), .B1(new_n652), .B2(new_n483), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n480), .A2(new_n650), .A3(new_n654), .ZN(new_n655));
  OAI21_X1  g469(.A(KEYINPUT95), .B1(new_n649), .B2(new_n655), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n616), .A2(new_n618), .A3(new_n653), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT95), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n657), .A2(new_n658), .A3(new_n608), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n648), .A2(new_n304), .A3(new_n656), .A4(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G128), .ZN(G30));
  XNOR2_X1  g475(.A(new_n443), .B(KEYINPUT38), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n364), .A2(new_n371), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT86), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n364), .A2(KEYINPUT86), .A3(new_n371), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n640), .A2(new_n603), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n667), .A2(new_n668), .A3(new_n480), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT98), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n662), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n564), .B1(new_n535), .B2(new_n552), .ZN(new_n672));
  XOR2_X1   g486(.A(new_n672), .B(KEYINPUT96), .Z(new_n673));
  INV_X1    g487(.A(new_n555), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n188), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(G472), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n574), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT97), .ZN(new_n678));
  AOI211_X1 g492(.A(new_n671), .B(new_n678), .C1(new_n670), .C2(new_n669), .ZN(new_n679));
  XOR2_X1   g493(.A(new_n653), .B(KEYINPUT39), .Z(new_n680));
  NAND2_X1  g494(.A1(new_n304), .A2(new_n680), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n681), .A2(KEYINPUT40), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(KEYINPUT40), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n679), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(new_n213), .ZN(G45));
  OAI211_X1 g499(.A(new_n601), .B(new_n654), .C1(new_n372), .C2(new_n373), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n648), .A2(new_n304), .A3(new_n608), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G146), .ZN(G48));
  OAI21_X1  g503(.A(new_n188), .B1(new_n273), .B2(new_n284), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(G469), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n285), .ZN(new_n692));
  INV_X1    g506(.A(new_n302), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n583), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n611), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT41), .B(G113), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G15));
  NAND2_X1  g513(.A1(new_n696), .A2(new_n619), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G116), .ZN(G18));
  NAND2_X1  g515(.A1(new_n374), .A2(new_n486), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n646), .A2(new_n702), .A3(new_n647), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n691), .A2(new_n302), .A3(new_n285), .A4(new_n608), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT99), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n704), .A2(new_n705), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n703), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(KEYINPUT100), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT100), .ZN(new_n710));
  OAI211_X1 g524(.A(new_n703), .B(new_n710), .C1(new_n706), .C2(new_n707), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G119), .ZN(G21));
  INV_X1    g527(.A(new_n522), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n586), .A2(G472), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n714), .A2(new_n715), .A3(new_n558), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n610), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT101), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n718), .B1(new_n374), .B2(new_n616), .ZN(new_n719));
  OAI211_X1 g533(.A(KEYINPUT101), .B(new_n480), .C1(new_n372), .C2(new_n373), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n694), .A2(new_n717), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G122), .ZN(G24));
  AND2_X1   g536(.A1(new_n715), .A2(new_n558), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n640), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n724), .A2(new_n686), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n725), .B1(new_n706), .B2(new_n707), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G125), .ZN(G27));
  INV_X1    g541(.A(KEYINPUT104), .ZN(new_n728));
  INV_X1    g542(.A(new_n272), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n287), .B1(new_n295), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(G902), .B1(new_n730), .B2(new_n283), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n298), .B1(new_n731), .B2(new_n187), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT102), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n297), .A2(new_n733), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n194), .A2(new_n272), .ZN(new_n735));
  AOI22_X1  g549(.A1(new_n271), .A2(new_n735), .B1(new_n286), .B2(new_n287), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(KEYINPUT102), .A3(G469), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n693), .B1(new_n732), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n435), .A2(new_n305), .A3(new_n442), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT103), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n728), .B1(new_n739), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n297), .A2(new_n733), .ZN(new_n744));
  AOI21_X1  g558(.A(KEYINPUT102), .B1(new_n736), .B2(G469), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n285), .B(new_n299), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  AND4_X1   g560(.A1(new_n728), .A2(new_n746), .A3(new_n742), .A4(new_n302), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n582), .B(new_n687), .C1(new_n743), .C2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(KEYINPUT105), .A2(KEYINPUT42), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT105), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT42), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n748), .A2(new_n749), .A3(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n746), .A2(new_n742), .A3(new_n302), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT104), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n739), .A2(new_n728), .A3(new_n742), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n583), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n757), .A2(new_n750), .A3(new_n751), .A4(new_n687), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n753), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(new_n202), .ZN(G33));
  XNOR2_X1  g574(.A(new_n657), .B(KEYINPUT106), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n582), .B(new_n761), .C1(new_n743), .C2(new_n747), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G134), .ZN(G36));
  XOR2_X1   g577(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n764));
  INV_X1    g578(.A(KEYINPUT43), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT107), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n374), .A2(new_n601), .ZN(new_n767));
  MUX2_X1   g581(.A(new_n764), .B(new_n766), .S(new_n767), .Z(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(new_n591), .A3(new_n640), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(KEYINPUT44), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n736), .B(KEYINPUT45), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n771), .A2(new_n187), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n298), .ZN(new_n773));
  AOI22_X1  g587(.A1(new_n773), .A2(KEYINPUT46), .B1(new_n187), .B2(new_n731), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n774), .B1(KEYINPUT46), .B2(new_n773), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n775), .A2(new_n302), .A3(new_n680), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n770), .A2(new_n742), .A3(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G137), .ZN(G39));
  NAND2_X1  g592(.A1(new_n775), .A2(new_n302), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(KEYINPUT47), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n646), .A2(new_n687), .A3(new_n522), .A4(new_n742), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G140), .ZN(G42));
  XOR2_X1   g597(.A(new_n692), .B(KEYINPUT109), .Z(new_n784));
  XOR2_X1   g598(.A(new_n784), .B(KEYINPUT49), .Z(new_n785));
  INV_X1    g599(.A(new_n662), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n767), .A2(new_n714), .A3(new_n302), .A4(new_n305), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT108), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n785), .A2(new_n786), .A3(new_n678), .A4(new_n788), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n487), .B(new_n304), .C1(new_n582), .C2(new_n642), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n582), .B(new_n694), .C1(new_n619), .C2(new_n611), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n443), .A2(new_n305), .A3(new_n609), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n665), .A2(new_n666), .A3(new_n480), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n792), .B1(new_n602), .B2(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n304), .A2(new_n794), .A3(new_n714), .A4(new_n590), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n790), .A2(new_n791), .A3(new_n721), .A4(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n796), .B1(new_n711), .B2(new_n709), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n725), .B1(new_n743), .B2(new_n747), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT110), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n478), .A2(new_n479), .A3(new_n654), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n799), .B1(new_n800), .B2(new_n618), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n616), .A2(new_n650), .A3(KEYINPUT110), .A4(new_n654), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n803), .A2(new_n742), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n648), .A2(new_n804), .A3(new_n304), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n762), .A2(new_n798), .A3(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n797), .A2(new_n806), .A3(new_n758), .A4(new_n753), .ZN(new_n807));
  OR2_X1    g621(.A1(new_n807), .A2(KEYINPUT111), .ZN(new_n808));
  AOI21_X1  g622(.A(KEYINPUT101), .B1(new_n667), .B2(new_n480), .ZN(new_n809));
  INV_X1    g623(.A(new_n720), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n635), .A2(new_n518), .A3(new_n654), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n812), .B1(new_n574), .B2(new_n676), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n811), .A2(new_n608), .A3(new_n739), .A4(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n726), .A2(new_n660), .A3(new_n688), .A4(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT52), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT112), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n574), .A2(new_n581), .ZN(new_n820));
  INV_X1    g634(.A(new_n647), .ZN(new_n821));
  AND4_X1   g635(.A1(new_n820), .A2(new_n821), .A3(new_n656), .A4(new_n659), .ZN(new_n822));
  NOR4_X1   g636(.A1(new_n646), .A2(new_n647), .A3(new_n686), .A4(new_n649), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n304), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n824), .A2(KEYINPUT52), .A3(new_n726), .A4(new_n814), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n817), .A2(new_n819), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n815), .A2(new_n818), .A3(new_n816), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(KEYINPUT53), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n808), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n807), .A2(KEYINPUT111), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n755), .A2(new_n756), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n648), .A2(new_n804), .ZN(new_n833));
  AOI22_X1  g647(.A1(new_n832), .A2(new_n725), .B1(new_n833), .B2(new_n304), .ZN(new_n834));
  AND4_X1   g648(.A1(new_n721), .A2(new_n790), .A3(new_n791), .A4(new_n795), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n712), .A2(new_n834), .A3(new_n835), .A4(new_n762), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n836), .A2(new_n759), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT113), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n838), .B1(new_n817), .B2(new_n825), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n817), .A2(new_n825), .A3(new_n838), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n837), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI22_X1  g655(.A1(new_n830), .A2(new_n831), .B1(KEYINPUT53), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT54), .ZN(new_n843));
  INV_X1    g657(.A(new_n759), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n844), .A2(KEYINPUT53), .A3(new_n797), .A4(new_n806), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT115), .B1(new_n845), .B2(new_n828), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n836), .A2(new_n759), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT115), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n848), .A2(new_n849), .A3(new_n827), .A4(new_n826), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n817), .A2(new_n825), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT113), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n817), .A2(new_n825), .A3(new_n838), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n807), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n856), .A2(KEYINPUT114), .A3(KEYINPUT53), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT114), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n858), .B1(new_n841), .B2(new_n847), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n851), .B(new_n852), .C1(new_n857), .C2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n843), .A2(new_n860), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n694), .A2(new_n742), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n768), .A2(new_n482), .A3(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n863), .A2(new_n724), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n768), .A2(new_n482), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n865), .A2(new_n716), .ZN(new_n866));
  AND4_X1   g680(.A1(new_n603), .A2(new_n866), .A3(new_n786), .A4(new_n694), .ZN(new_n867));
  OR2_X1    g681(.A1(new_n867), .A2(KEYINPUT50), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(KEYINPUT50), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n864), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n780), .B1(new_n302), .B2(new_n784), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n871), .A2(new_n742), .A3(new_n866), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n678), .A2(new_n862), .A3(new_n714), .A4(new_n482), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(KEYINPUT116), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(new_n374), .A3(new_n600), .A4(new_n598), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n870), .A2(new_n872), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT51), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n876), .A2(new_n877), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n863), .A2(new_n583), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(KEYINPUT48), .Z(new_n881));
  NAND3_X1  g695(.A1(new_n874), .A2(new_n667), .A3(new_n601), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n192), .A2(G952), .ZN(new_n883));
  INV_X1    g697(.A(new_n706), .ZN(new_n884));
  INV_X1    g698(.A(new_n707), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n883), .B1(new_n866), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n881), .A2(new_n882), .A3(new_n887), .ZN(new_n888));
  NOR4_X1   g702(.A1(new_n861), .A2(new_n878), .A3(new_n879), .A4(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(G952), .A2(G953), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n789), .B1(new_n889), .B2(new_n890), .ZN(G75));
  NAND2_X1  g705(.A1(new_n410), .A2(new_n419), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(new_n416), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT55), .Z(new_n894));
  INV_X1    g708(.A(KEYINPUT117), .ZN(new_n895));
  OAI21_X1  g709(.A(KEYINPUT114), .B1(new_n856), .B2(KEYINPUT53), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n841), .A2(new_n858), .A3(new_n847), .ZN(new_n897));
  AOI22_X1  g711(.A1(new_n896), .A2(new_n897), .B1(new_n850), .B2(new_n846), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n895), .B1(new_n898), .B2(new_n188), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n851), .B1(new_n857), .B2(new_n859), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n900), .A2(KEYINPUT117), .A3(G902), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  AOI211_X1 g717(.A(KEYINPUT56), .B(new_n894), .C1(new_n903), .C2(new_n376), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n898), .A2(new_n188), .A3(new_n605), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n894), .B1(new_n905), .B2(KEYINPUT56), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n192), .A2(G952), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n904), .A2(new_n909), .ZN(G51));
  NOR2_X1   g724(.A1(new_n273), .A2(new_n284), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n900), .A2(KEYINPUT54), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n860), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n298), .B(KEYINPUT57), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n911), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n899), .A2(new_n772), .A3(new_n901), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n908), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT118), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI211_X1 g733(.A(KEYINPUT118), .B(new_n908), .C1(new_n915), .C2(new_n916), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(G54));
  NAND2_X1  g735(.A1(KEYINPUT58), .A2(G475), .ZN(new_n922));
  OAI221_X1 g736(.A(new_n357), .B1(new_n347), .B2(new_n358), .C1(new_n902), .C2(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n903), .A2(KEYINPUT58), .A3(G475), .A4(new_n359), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n923), .A2(new_n924), .A3(new_n908), .ZN(G60));
  XNOR2_X1  g739(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n926));
  NAND2_X1  g740(.A1(G478), .A2(G902), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n926), .B(new_n927), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n913), .A2(new_n597), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n597), .B1(new_n861), .B2(new_n928), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n929), .A2(new_n930), .A3(new_n907), .ZN(G63));
  OAI21_X1  g745(.A(KEYINPUT60), .B1(new_n469), .B2(new_n188), .ZN(new_n932));
  OR3_X1    g746(.A1(new_n469), .A2(new_n188), .A3(KEYINPUT60), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n900), .A2(new_n631), .A3(new_n932), .A4(new_n933), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n900), .A2(new_n932), .A3(new_n933), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n908), .B(new_n934), .C1(new_n935), .C2(new_n519), .ZN(new_n936));
  XOR2_X1   g750(.A(KEYINPUT120), .B(KEYINPUT61), .Z(new_n937));
  XNOR2_X1  g751(.A(new_n936), .B(new_n937), .ZN(G66));
  OAI21_X1  g752(.A(G953), .B1(new_n484), .B2(new_n414), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT121), .ZN(new_n940));
  INV_X1    g754(.A(new_n797), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n940), .B1(new_n941), .B2(new_n192), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n892), .B1(G898), .B2(new_n192), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n942), .B(new_n943), .Z(G69));
  XNOR2_X1  g758(.A(new_n568), .B(new_n352), .ZN(new_n945));
  INV_X1    g759(.A(new_n824), .ZN(new_n946));
  INV_X1    g760(.A(new_n726), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n684), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT62), .ZN(new_n951));
  INV_X1    g765(.A(new_n681), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n602), .A2(new_n793), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n952), .A2(new_n582), .A3(new_n742), .A4(new_n953), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT123), .Z(new_n955));
  AND2_X1   g769(.A1(new_n782), .A2(new_n777), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n951), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n957), .A2(new_n192), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT122), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n945), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n958), .A2(KEYINPUT122), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n776), .A2(new_n582), .A3(new_n608), .A4(new_n811), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT125), .Z(new_n963));
  NAND4_X1  g777(.A1(new_n956), .A2(new_n762), .A3(new_n948), .A4(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n192), .B1(new_n964), .B2(new_n759), .ZN(new_n965));
  INV_X1    g779(.A(G900), .ZN(new_n966));
  AOI21_X1  g780(.A(KEYINPUT124), .B1(new_n966), .B2(G953), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n966), .A2(KEYINPUT124), .A3(G953), .ZN(new_n968));
  NOR3_X1   g782(.A1(new_n945), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n965), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n960), .B1(new_n961), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n192), .B1(G227), .B2(G900), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n960), .B(new_n972), .C1(new_n961), .C2(new_n970), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(G72));
  NAND2_X1  g790(.A1(G472), .A2(G902), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT63), .Z(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n979), .B1(new_n576), .B2(new_n555), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT126), .Z(new_n981));
  NAND2_X1  g795(.A1(new_n842), .A2(new_n981), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT127), .Z(new_n983));
  NOR3_X1   g797(.A1(new_n964), .A2(new_n759), .A3(new_n941), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n564), .B(new_n569), .C1(new_n984), .C2(new_n979), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n978), .B1(new_n957), .B2(new_n941), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n986), .A2(new_n540), .A3(new_n575), .ZN(new_n987));
  AND4_X1   g801(.A1(new_n908), .A2(new_n983), .A3(new_n985), .A4(new_n987), .ZN(G57));
endmodule


