//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 1 1 0 1 1 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 1 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 0 1 0 1 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954;
  XNOR2_X1  g000(.A(KEYINPUT66), .B(G131), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  NOR2_X1   g002(.A1(G237), .A2(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n189), .A2(G143), .A3(G214), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  AOI21_X1  g005(.A(G143), .B1(new_n189), .B2(G214), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n188), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n192), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(new_n187), .A3(new_n190), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n193), .A2(new_n195), .A3(KEYINPUT91), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n191), .A2(new_n192), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT91), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(new_n187), .ZN(new_n199));
  AOI21_X1  g013(.A(KEYINPUT17), .B1(new_n196), .B2(new_n199), .ZN(new_n200));
  OR2_X1    g014(.A1(new_n200), .A2(KEYINPUT94), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT16), .ZN(new_n202));
  OR2_X1    g016(.A1(G125), .A2(G140), .ZN(new_n203));
  NAND2_X1  g017(.A1(G125), .A2(G140), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G125), .ZN(new_n206));
  NOR3_X1   g020(.A1(new_n206), .A2(KEYINPUT16), .A3(G140), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G146), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n210), .B1(new_n205), .B2(new_n207), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n209), .A2(KEYINPUT79), .A3(new_n211), .ZN(new_n212));
  OR3_X1    g026(.A1(new_n208), .A2(KEYINPUT79), .A3(G146), .ZN(new_n213));
  INV_X1    g027(.A(new_n193), .ZN(new_n214));
  AOI22_X1  g028(.A1(new_n212), .A2(new_n213), .B1(KEYINPUT17), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n200), .A2(KEYINPUT94), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n201), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(G113), .B(G122), .ZN(new_n218));
  INV_X1    g032(.A(G104), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n218), .B(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT18), .A2(G131), .ZN(new_n221));
  OR2_X1    g035(.A1(new_n197), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n203), .A2(new_n204), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n223), .B(new_n210), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n197), .A2(new_n221), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n222), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n217), .A2(new_n220), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n196), .A2(new_n199), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT92), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT19), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n223), .B1(KEYINPUT93), .B2(new_n230), .ZN(new_n231));
  OR2_X1    g045(.A1(new_n230), .A2(KEYINPUT93), .ZN(new_n232));
  XNOR2_X1  g046(.A(new_n231), .B(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(new_n210), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT92), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n196), .A2(new_n199), .A3(new_n235), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n229), .A2(new_n234), .A3(new_n209), .A4(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(new_n226), .ZN(new_n238));
  INV_X1    g052(.A(new_n220), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n227), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G475), .ZN(new_n242));
  INV_X1    g056(.A(G902), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT20), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AND3_X1   g060(.A1(new_n217), .A2(new_n220), .A3(new_n226), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n220), .B1(new_n217), .B2(new_n226), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n243), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G475), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n241), .A2(KEYINPUT20), .A3(new_n242), .A4(new_n243), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n246), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G953), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n253), .A2(G952), .ZN(new_n254));
  INV_X1    g068(.A(G234), .ZN(new_n255));
  INV_X1    g069(.A(G237), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT21), .B(G898), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n259), .B(KEYINPUT99), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  AOI211_X1 g075(.A(new_n243), .B(new_n253), .C1(G234), .C2(G237), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n258), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  XOR2_X1   g077(.A(KEYINPUT9), .B(G234), .Z(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G217), .ZN(new_n266));
  NOR3_X1   g080(.A1(new_n265), .A2(new_n266), .A3(G953), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G107), .ZN(new_n269));
  INV_X1    g083(.A(G116), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G122), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT95), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n271), .B(new_n272), .ZN(new_n273));
  OR2_X1    g087(.A1(new_n270), .A2(G122), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n273), .A2(KEYINPUT96), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT96), .B1(new_n273), .B2(new_n274), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n269), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n273), .A2(KEYINPUT14), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n274), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n273), .A2(KEYINPUT14), .ZN(new_n281));
  OAI21_X1  g095(.A(G107), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G128), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G143), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT97), .ZN(new_n285));
  INV_X1    g099(.A(G143), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n285), .B1(G128), .B2(new_n286), .ZN(new_n287));
  NOR3_X1   g101(.A1(new_n283), .A2(KEYINPUT97), .A3(G143), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n284), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n289), .B(G134), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n278), .A2(new_n282), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G134), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT13), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n293), .B1(new_n284), .B2(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n289), .B(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n277), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n297), .A2(G107), .A3(new_n275), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n296), .B1(new_n278), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n268), .B1(new_n292), .B2(new_n299), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n278), .A2(new_n298), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n291), .B(new_n267), .C1(new_n301), .C2(new_n296), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT98), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n300), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  OAI211_X1 g118(.A(KEYINPUT98), .B(new_n268), .C1(new_n292), .C2(new_n299), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n243), .A3(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G478), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n307), .A2(KEYINPUT15), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n308), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n304), .A2(new_n243), .A3(new_n305), .A4(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n252), .A2(new_n263), .A3(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(G214), .B1(G237), .B2(G902), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  XOR2_X1   g129(.A(G110), .B(G122), .Z(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT3), .B1(new_n219), .B2(G107), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT82), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n219), .A2(G107), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT3), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n269), .A2(G104), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  OAI211_X1 g139(.A(KEYINPUT82), .B(KEYINPUT3), .C1(new_n219), .C2(G107), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n320), .A2(new_n323), .A3(new_n325), .A4(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G101), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n324), .B1(new_n322), .B2(new_n321), .ZN(new_n329));
  INV_X1    g143(.A(G101), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n329), .A2(new_n330), .A3(new_n320), .A4(new_n326), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n328), .A2(KEYINPUT4), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT71), .ZN(new_n333));
  NAND2_X1  g147(.A1(KEYINPUT2), .A2(G113), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT70), .B1(KEYINPUT2), .B2(G113), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NOR3_X1   g150(.A1(KEYINPUT70), .A2(KEYINPUT2), .A3(G113), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n334), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(G116), .B(G119), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  OR3_X1    g155(.A1(KEYINPUT70), .A2(KEYINPUT2), .A3(G113), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n335), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n339), .B1(new_n343), .B2(new_n334), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n333), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n338), .A2(new_n340), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n343), .A2(new_n334), .A3(new_n339), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n347), .A3(KEYINPUT71), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT4), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n327), .A2(new_n349), .A3(G101), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n332), .A2(new_n345), .A3(new_n348), .A4(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(G101), .B1(new_n324), .B2(new_n321), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n331), .A2(new_n352), .ZN(new_n353));
  NOR3_X1   g167(.A1(new_n270), .A2(KEYINPUT5), .A3(G119), .ZN(new_n354));
  OR2_X1    g168(.A1(new_n354), .A2(KEYINPUT86), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n339), .A2(KEYINPUT5), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(KEYINPUT86), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n355), .A2(G113), .A3(new_n356), .A4(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n353), .A2(new_n347), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n317), .B1(new_n351), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n351), .A2(new_n359), .A3(new_n317), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n361), .A2(KEYINPUT87), .A3(KEYINPUT6), .A4(new_n362), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n351), .A2(new_n359), .A3(new_n317), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT6), .ZN(new_n365));
  NOR3_X1   g179(.A1(new_n364), .A2(new_n360), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n351), .A2(new_n359), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(new_n365), .A3(new_n316), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT87), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n363), .B1(new_n366), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n210), .A2(G143), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n286), .A2(KEYINPUT64), .A3(G146), .ZN(new_n373));
  AOI21_X1  g187(.A(KEYINPUT64), .B1(new_n286), .B2(G146), .ZN(new_n374));
  OAI211_X1 g188(.A(G128), .B(new_n372), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n286), .A2(G146), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n210), .A2(G143), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n375), .B(KEYINPUT0), .C1(G128), .C2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT0), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n380), .B1(new_n378), .B2(new_n283), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n206), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT1), .B1(new_n286), .B2(G146), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT68), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n372), .A2(KEYINPUT68), .A3(KEYINPUT1), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(G128), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n378), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT64), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n390), .B1(new_n210), .B2(G143), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n286), .A2(KEYINPUT64), .A3(G146), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n376), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT1), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(new_n394), .A3(G128), .ZN(new_n395));
  AOI21_X1  g209(.A(G125), .B1(new_n389), .B2(new_n395), .ZN(new_n396));
  OR3_X1    g210(.A1(new_n382), .A2(KEYINPUT89), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n253), .A2(G224), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n398), .B(KEYINPUT88), .ZN(new_n399));
  OAI21_X1  g213(.A(KEYINPUT89), .B1(new_n382), .B2(new_n396), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n397), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n399), .B1(new_n397), .B2(new_n400), .ZN(new_n402));
  OR2_X1    g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n371), .A2(new_n403), .ZN(new_n404));
  XOR2_X1   g218(.A(new_n316), .B(KEYINPUT8), .Z(new_n405));
  INV_X1    g219(.A(new_n359), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n353), .B1(new_n347), .B2(new_n358), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n382), .ZN(new_n409));
  INV_X1    g223(.A(new_n396), .ZN(new_n410));
  AND4_X1   g224(.A1(KEYINPUT7), .A2(new_n409), .A3(new_n410), .A4(new_n399), .ZN(new_n411));
  AOI22_X1  g225(.A1(new_n409), .A2(new_n410), .B1(KEYINPUT7), .B2(new_n399), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n408), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(KEYINPUT90), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT90), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n415), .B(new_n408), .C1(new_n411), .C2(new_n412), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n414), .A2(new_n416), .A3(new_n362), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n404), .A2(new_n417), .A3(new_n243), .ZN(new_n418));
  OAI21_X1  g232(.A(G210), .B1(G237), .B2(G902), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(G902), .B1(new_n371), .B2(new_n403), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n422), .A2(new_n419), .A3(new_n417), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n315), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(G221), .B1(new_n265), .B2(G902), .ZN(new_n425));
  INV_X1    g239(.A(G469), .ZN(new_n426));
  XNOR2_X1  g240(.A(G110), .B(G140), .ZN(new_n427));
  INV_X1    g241(.A(G227), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n428), .A2(G953), .ZN(new_n429));
  XOR2_X1   g243(.A(new_n427), .B(new_n429), .Z(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT10), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n383), .A2(G128), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(KEYINPUT83), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT83), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n283), .B1(new_n372), .B2(KEYINPUT1), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n436), .B1(new_n393), .B2(new_n437), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n435), .A2(new_n438), .A3(new_n395), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n331), .A2(new_n352), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n432), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n379), .A2(new_n381), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n332), .A2(new_n442), .A3(new_n350), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT65), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n444), .B1(new_n293), .B2(G137), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(KEYINPUT11), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n293), .A2(G137), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT11), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n444), .B(new_n448), .C1(new_n293), .C2(G137), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n446), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n450), .A2(KEYINPUT67), .A3(G131), .ZN(new_n451));
  AOI21_X1  g265(.A(KEYINPUT67), .B1(new_n450), .B2(G131), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n446), .A2(new_n187), .A3(new_n447), .A4(new_n449), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NOR3_X1   g268(.A1(new_n451), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n432), .B1(new_n389), .B2(new_n395), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n353), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n441), .A2(new_n443), .A3(new_n455), .A4(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(KEYINPUT84), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n435), .A2(new_n438), .A3(new_n395), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n353), .A2(new_n460), .ZN(new_n461));
  AOI22_X1  g275(.A1(new_n461), .A2(new_n432), .B1(new_n353), .B2(new_n456), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT84), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n462), .A2(new_n463), .A3(new_n455), .A4(new_n443), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n431), .B1(new_n459), .B2(new_n464), .ZN(new_n465));
  AOI211_X1 g279(.A(new_n283), .B(new_n376), .C1(new_n391), .C2(new_n392), .ZN(new_n466));
  AOI22_X1  g280(.A1(new_n466), .A2(new_n394), .B1(new_n387), .B2(new_n388), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n440), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n461), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n450), .A2(G131), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT67), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n450), .A2(KEYINPUT67), .A3(G131), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n453), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n469), .A2(KEYINPUT12), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(KEYINPUT85), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n469), .A2(new_n474), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT12), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT85), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n469), .A2(new_n480), .A3(KEYINPUT12), .A4(new_n474), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n476), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n465), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n459), .A2(new_n464), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n462), .A2(new_n443), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n474), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n430), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n426), .B(new_n243), .C1(new_n483), .C2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(G469), .A2(G902), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n465), .A2(new_n486), .ZN(new_n490));
  AND2_X1   g304(.A1(new_n482), .A2(new_n484), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n490), .B1(new_n491), .B2(new_n430), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n488), .B(new_n489), .C1(new_n426), .C2(new_n492), .ZN(new_n493));
  AND4_X1   g307(.A1(new_n313), .A2(new_n424), .A3(new_n425), .A4(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT32), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT31), .ZN(new_n496));
  INV_X1    g310(.A(new_n447), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n293), .A2(G137), .ZN(new_n498));
  OAI21_X1  g312(.A(G131), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n453), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(KEYINPUT69), .B1(new_n467), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n389), .A2(new_n395), .ZN(new_n502));
  INV_X1    g316(.A(new_n500), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT69), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n442), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n501), .B(new_n505), .C1(new_n455), .C2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT30), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n345), .A2(new_n348), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  AOI22_X1  g325(.A1(new_n474), .A2(new_n442), .B1(new_n502), .B2(new_n503), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT30), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n509), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT72), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n509), .A2(KEYINPUT72), .A3(new_n511), .A4(new_n513), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n510), .A2(KEYINPUT73), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT73), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n345), .A2(new_n520), .A3(new_n348), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n512), .ZN(new_n523));
  XOR2_X1   g337(.A(KEYINPUT74), .B(KEYINPUT27), .Z(new_n524));
  NAND2_X1  g338(.A1(new_n189), .A2(G210), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n524), .B(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT26), .B(G101), .ZN(new_n527));
  XOR2_X1   g341(.A(new_n526), .B(new_n527), .Z(new_n528));
  NAND2_X1  g342(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n496), .B1(new_n518), .B2(new_n530), .ZN(new_n531));
  AOI211_X1 g345(.A(KEYINPUT31), .B(new_n529), .C1(new_n516), .C2(new_n517), .ZN(new_n532));
  INV_X1    g346(.A(new_n523), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n533), .A2(KEYINPUT28), .ZN(new_n534));
  INV_X1    g348(.A(new_n507), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n523), .B1(new_n535), .B2(new_n510), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT28), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n528), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n531), .A2(new_n532), .A3(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(G472), .A2(G902), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n495), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n518), .A2(new_n530), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT31), .ZN(new_n544));
  INV_X1    g358(.A(new_n538), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n518), .A2(new_n496), .A3(new_n530), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n547), .A2(KEYINPUT32), .A3(new_n540), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n534), .A2(new_n537), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n528), .ZN(new_n550));
  INV_X1    g364(.A(new_n528), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n518), .A2(new_n523), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT29), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n522), .ZN(new_n554));
  INV_X1    g368(.A(new_n512), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n556), .A2(KEYINPUT75), .A3(new_n523), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT75), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n554), .A2(new_n555), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n557), .A2(KEYINPUT28), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n534), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n528), .A2(KEYINPUT29), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n243), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(G472), .B1(new_n553), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n542), .A2(new_n548), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(G119), .ZN(new_n566));
  OAI21_X1  g380(.A(KEYINPUT77), .B1(new_n566), .B2(G128), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT23), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(G128), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT23), .ZN(new_n570));
  OAI211_X1 g384(.A(KEYINPUT77), .B(new_n570), .C1(new_n566), .C2(G128), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n568), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G110), .ZN(new_n573));
  XOR2_X1   g387(.A(new_n573), .B(KEYINPUT78), .Z(new_n574));
  INV_X1    g388(.A(KEYINPUT76), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n569), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n566), .A2(KEYINPUT76), .A3(G128), .ZN(new_n577));
  AOI22_X1  g391(.A1(new_n576), .A2(new_n577), .B1(G119), .B2(new_n283), .ZN(new_n578));
  XOR2_X1   g392(.A(KEYINPUT24), .B(G110), .Z(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n574), .A2(new_n580), .A3(new_n213), .A4(new_n212), .ZN(new_n581));
  OR3_X1    g395(.A1(new_n578), .A2(KEYINPUT80), .A3(new_n579), .ZN(new_n582));
  OAI21_X1  g396(.A(KEYINPUT80), .B1(new_n578), .B2(new_n579), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n582), .B(new_n583), .C1(G110), .C2(new_n572), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n223), .A2(new_n210), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n584), .A2(new_n209), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n253), .A2(G221), .A3(G234), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(KEYINPUT22), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(G137), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n581), .A2(new_n586), .A3(new_n590), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n243), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n266), .B1(G234), .B2(new_n243), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n599));
  INV_X1    g413(.A(new_n597), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n592), .A2(new_n243), .A3(new_n600), .A4(new_n593), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n598), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n596), .B1(new_n602), .B2(new_n595), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n494), .A2(new_n565), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G101), .ZN(G3));
  NAND2_X1  g419(.A1(new_n547), .A2(new_n243), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n606), .A2(KEYINPUT100), .A3(G472), .ZN(new_n607));
  NAND2_X1  g421(.A1(KEYINPUT100), .A2(G472), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n547), .A2(new_n243), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n425), .ZN(new_n611));
  AOI211_X1 g425(.A(new_n596), .B(new_n611), .C1(new_n602), .C2(new_n595), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n493), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT33), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n304), .A2(new_n615), .A3(new_n305), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n300), .A2(new_n302), .A3(KEYINPUT33), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n616), .A2(G478), .A3(new_n243), .A4(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n306), .A2(new_n307), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n252), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n621), .A2(new_n263), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n614), .A2(new_n424), .A3(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT34), .B(G104), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G6));
  XNOR2_X1  g439(.A(new_n263), .B(KEYINPUT101), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n422), .A2(new_n419), .A3(new_n417), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n419), .B1(new_n422), .B2(new_n417), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n314), .B(new_n626), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n312), .A2(new_n250), .A3(new_n246), .A4(new_n251), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n614), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT35), .B(G107), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  NAND2_X1  g448(.A1(new_n602), .A2(new_n595), .ZN(new_n635));
  XOR2_X1   g449(.A(new_n587), .B(KEYINPUT102), .Z(new_n636));
  OR2_X1    g450(.A1(new_n591), .A2(KEYINPUT36), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n595), .A2(G902), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n635), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n494), .A2(new_n609), .A3(new_n607), .A4(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(new_n642), .B(KEYINPUT37), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G110), .ZN(G12));
  NAND2_X1  g458(.A1(new_n493), .A2(new_n425), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n314), .B1(new_n627), .B2(new_n628), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(G900), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n262), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n257), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n630), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n565), .A2(new_n647), .A3(new_n641), .A4(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G128), .ZN(G30));
  NAND2_X1  g468(.A1(new_n421), .A2(new_n423), .ZN(new_n655));
  XOR2_X1   g469(.A(new_n655), .B(KEYINPUT38), .Z(new_n656));
  INV_X1    g470(.A(new_n312), .ZN(new_n657));
  INV_X1    g471(.A(new_n252), .ZN(new_n658));
  OR3_X1    g472(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(new_n650), .B(KEYINPUT39), .Z(new_n660));
  OR2_X1    g474(.A1(new_n645), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT40), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n542), .A2(new_n548), .ZN(new_n663));
  AND2_X1   g477(.A1(new_n557), .A2(new_n559), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n243), .B1(new_n664), .B2(new_n528), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n551), .B1(new_n518), .B2(new_n523), .ZN(new_n666));
  OAI21_X1  g480(.A(G472), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n641), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR4_X1   g484(.A1(new_n659), .A2(new_n662), .A3(new_n315), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT103), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G143), .ZN(G45));
  NAND3_X1  g487(.A1(new_n252), .A2(new_n620), .A3(new_n650), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n565), .A2(new_n647), .A3(new_n641), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G146), .ZN(G48));
  NAND2_X1  g491(.A1(new_n484), .A2(new_n486), .ZN(new_n678));
  AOI22_X1  g492(.A1(new_n678), .A2(new_n431), .B1(new_n465), .B2(new_n482), .ZN(new_n679));
  OAI21_X1  g493(.A(G469), .B1(new_n679), .B2(G902), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n680), .A2(new_n425), .A3(new_n488), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT104), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n680), .A2(KEYINPUT104), .A3(new_n488), .A4(new_n425), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n683), .A2(new_n424), .A3(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n686), .A2(new_n565), .A3(new_n603), .A4(new_n622), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT41), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G113), .ZN(G15));
  AND2_X1   g503(.A1(new_n565), .A2(new_n603), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT105), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n683), .A2(new_n684), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n690), .A2(new_n691), .A3(new_n631), .A4(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n565), .A2(new_n692), .A3(new_n631), .A4(new_n603), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(KEYINPUT105), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G116), .ZN(G18));
  NAND2_X1  g511(.A1(new_n685), .A2(KEYINPUT106), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n683), .A2(new_n424), .A3(new_n699), .A4(new_n684), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n701), .A2(new_n565), .A3(new_n313), .A4(new_n641), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G119), .ZN(G21));
  NOR2_X1   g517(.A1(new_n658), .A2(new_n657), .ZN(new_n704));
  AND4_X1   g518(.A1(new_n424), .A2(new_n704), .A3(new_n683), .A4(new_n684), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n561), .A2(new_n551), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT107), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n706), .A2(new_n544), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n528), .B1(new_n560), .B2(new_n534), .ZN(new_n709));
  OAI21_X1  g523(.A(KEYINPUT107), .B1(new_n709), .B2(new_n531), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n708), .A2(new_n710), .A3(new_n546), .ZN(new_n711));
  AOI22_X1  g525(.A1(new_n711), .A2(new_n540), .B1(new_n606), .B2(G472), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n705), .A2(new_n603), .A3(new_n626), .A4(new_n712), .ZN(new_n713));
  XOR2_X1   g527(.A(new_n713), .B(KEYINPUT108), .Z(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G122), .ZN(G24));
  AOI21_X1  g529(.A(new_n674), .B1(new_n698), .B2(new_n700), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n712), .A2(new_n641), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(KEYINPUT109), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G125), .ZN(G27));
  NAND3_X1  g534(.A1(new_n421), .A2(new_n314), .A3(new_n423), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n645), .A2(new_n721), .A3(new_n674), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n722), .A2(new_n565), .A3(new_n603), .ZN(new_n723));
  NOR2_X1   g537(.A1(KEYINPUT110), .A2(KEYINPUT42), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n724), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n722), .A2(new_n565), .A3(new_n603), .A4(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(KEYINPUT111), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n725), .A2(KEYINPUT111), .A3(new_n727), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(KEYINPUT112), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G131), .ZN(G33));
  INV_X1    g547(.A(new_n613), .ZN(new_n734));
  INV_X1    g548(.A(new_n721), .ZN(new_n735));
  AND4_X1   g549(.A1(new_n565), .A2(new_n734), .A3(new_n652), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(new_n293), .ZN(G36));
  NAND2_X1  g551(.A1(new_n658), .A2(new_n620), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT43), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n738), .B1(KEYINPUT113), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(KEYINPUT113), .B(KEYINPUT43), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n740), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n610), .A3(new_n641), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT44), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n744), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(new_n735), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT114), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n492), .B(KEYINPUT45), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(G469), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n489), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT46), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n488), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n751), .A2(new_n752), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n425), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(new_n660), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT114), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n745), .A2(new_n758), .A3(new_n735), .A4(new_n746), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n748), .A2(new_n757), .A3(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G137), .ZN(G39));
  XNOR2_X1  g575(.A(new_n756), .B(KEYINPUT47), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n735), .A2(new_n675), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n565), .A2(new_n603), .ZN(new_n764));
  OR3_X1    g578(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G140), .ZN(G42));
  INV_X1    g580(.A(new_n668), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n680), .A2(new_n488), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n658), .B(new_n620), .C1(new_n768), .C2(KEYINPUT49), .ZN(new_n769));
  AOI211_X1 g583(.A(new_n315), .B(new_n769), .C1(KEYINPUT49), .C2(new_n768), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n767), .A2(new_n770), .A3(new_n612), .A4(new_n656), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n653), .A2(new_n676), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n772), .B1(new_n717), .B2(new_n716), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n646), .A2(new_n657), .A3(new_n658), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n650), .A2(KEYINPUT116), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n650), .A2(KEYINPUT116), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n645), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n668), .A2(new_n669), .A3(new_n774), .A4(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT52), .B1(new_n773), .B2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n772), .ZN(new_n780));
  AND4_X1   g594(.A1(KEYINPUT52), .A2(new_n780), .A3(new_n718), .A4(new_n778), .ZN(new_n781));
  OAI21_X1  g595(.A(KEYINPUT53), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n694), .B(new_n691), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n698), .A2(new_n700), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n565), .A2(new_n313), .A3(new_n641), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n687), .B(new_n713), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n725), .A2(new_n727), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n712), .A2(new_n722), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n252), .A2(new_n312), .A3(new_n651), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n565), .A2(new_n735), .A3(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n789), .B1(new_n791), .B2(new_n645), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n736), .B1(new_n792), .B2(new_n641), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n621), .A2(new_n630), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(new_n629), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n795), .A2(new_n609), .A3(new_n607), .A4(new_n734), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n642), .A2(new_n604), .A3(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n787), .A2(new_n788), .A3(new_n793), .A4(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n782), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n642), .A2(new_n796), .A3(new_n604), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n783), .A2(new_n786), .A3(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n801), .A2(KEYINPUT115), .A3(new_n731), .A4(new_n793), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n725), .A2(KEYINPUT111), .A3(new_n727), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n793), .B1(new_n804), .B2(new_n728), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n713), .A2(new_n687), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n696), .A2(new_n806), .A3(new_n797), .A4(new_n702), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n803), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n773), .A2(KEYINPUT52), .A3(new_n778), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n780), .A2(new_n718), .A3(new_n778), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n802), .A2(new_n808), .A3(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n799), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n815), .B1(new_n809), .B2(new_n812), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n802), .A2(new_n819), .A3(new_n808), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n802), .A2(new_n819), .A3(new_n808), .A4(KEYINPUT117), .ZN(new_n823));
  AOI22_X1  g637(.A1(new_n822), .A2(new_n823), .B1(new_n815), .B2(new_n814), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n818), .B1(new_n824), .B2(new_n817), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT51), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n768), .B(KEYINPUT119), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n762), .B1(new_n425), .B2(new_n827), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n742), .A2(new_n258), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n712), .A2(new_n603), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(KEYINPUT118), .B1(new_n831), .B2(new_n721), .ZN(new_n832));
  OR3_X1    g646(.A1(new_n831), .A2(KEYINPUT118), .A3(new_n721), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n828), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n829), .A2(new_n692), .A3(new_n830), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n656), .A2(new_n315), .ZN(new_n836));
  OR4_X1    g650(.A1(KEYINPUT120), .A2(new_n835), .A3(KEYINPUT50), .A4(new_n836), .ZN(new_n837));
  OAI22_X1  g651(.A1(new_n835), .A2(new_n836), .B1(KEYINPUT120), .B2(KEYINPUT50), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n692), .A2(new_n735), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n829), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(new_n717), .ZN(new_n841));
  AND4_X1   g655(.A1(new_n603), .A2(new_n767), .A3(new_n258), .A4(new_n839), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n842), .A2(new_n658), .A3(new_n619), .A4(new_n618), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n837), .A2(new_n838), .A3(new_n841), .A4(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n826), .B1(new_n834), .B2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT121), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT48), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n840), .A2(new_n690), .A3(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n846), .A2(KEYINPUT48), .ZN(new_n849));
  XOR2_X1   g663(.A(new_n848), .B(new_n849), .Z(new_n850));
  AND3_X1   g664(.A1(new_n837), .A2(new_n841), .A3(new_n843), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n828), .A2(new_n832), .A3(new_n833), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n851), .A2(new_n852), .A3(KEYINPUT51), .A4(new_n838), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n845), .A2(new_n254), .A3(new_n850), .A4(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n831), .A2(new_n784), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n842), .A2(new_n252), .A3(new_n620), .ZN(new_n856));
  NOR4_X1   g670(.A1(new_n825), .A2(new_n854), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(G952), .A2(G953), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n771), .B1(new_n857), .B2(new_n858), .ZN(G75));
  NAND2_X1  g673(.A1(new_n814), .A2(new_n815), .ZN(new_n860));
  INV_X1    g674(.A(new_n799), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n862), .A2(new_n863), .A3(G902), .ZN(new_n864));
  OAI21_X1  g678(.A(KEYINPUT122), .B1(new_n816), .B2(new_n243), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n864), .A2(new_n865), .A3(new_n420), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT56), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n371), .B(new_n403), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(KEYINPUT55), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n866), .A2(new_n867), .A3(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n253), .A2(G952), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n872), .B(KEYINPUT123), .Z(new_n873));
  NAND3_X1  g687(.A1(new_n862), .A2(G210), .A3(G902), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n867), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n873), .B1(new_n875), .B2(new_n869), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n871), .A2(new_n876), .ZN(G51));
  NAND2_X1  g691(.A1(new_n489), .A2(KEYINPUT57), .ZN(new_n878));
  INV_X1    g692(.A(new_n818), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n816), .A2(new_n817), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n489), .A2(KEYINPUT57), .ZN(new_n882));
  OAI22_X1  g696(.A1(new_n881), .A2(new_n882), .B1(new_n487), .B2(new_n483), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n864), .A2(new_n865), .A3(G469), .A4(new_n749), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n872), .B1(new_n883), .B2(new_n884), .ZN(G54));
  INV_X1    g699(.A(new_n872), .ZN(new_n886));
  AND2_X1   g700(.A1(KEYINPUT58), .A2(G475), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n864), .A2(new_n865), .A3(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n241), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n886), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n888), .A2(new_n889), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n888), .A2(KEYINPUT124), .A3(new_n889), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n890), .B1(new_n893), .B2(new_n894), .ZN(G60));
  AND2_X1   g709(.A1(new_n616), .A2(new_n617), .ZN(new_n896));
  NAND2_X1  g710(.A1(G478), .A2(G902), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT59), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n896), .B(new_n898), .C1(new_n879), .C2(new_n880), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n896), .B1(new_n825), .B2(new_n898), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n900), .A2(new_n901), .A3(new_n873), .ZN(G63));
  NAND2_X1  g716(.A1(G217), .A2(G902), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT60), .Z(new_n904));
  NAND2_X1  g718(.A1(new_n862), .A2(new_n904), .ZN(new_n905));
  OR2_X1    g719(.A1(new_n905), .A2(new_n638), .ZN(new_n906));
  INV_X1    g720(.A(new_n873), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n592), .A2(new_n593), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n906), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT61), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n906), .A2(KEYINPUT61), .A3(new_n907), .A4(new_n909), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(G66));
  AOI21_X1  g728(.A(new_n253), .B1(new_n260), .B2(G224), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n915), .B1(new_n807), .B2(new_n253), .ZN(new_n916));
  INV_X1    g730(.A(new_n371), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n917), .B1(G898), .B2(new_n253), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n916), .B(new_n918), .Z(G69));
  NAND3_X1  g733(.A1(new_n757), .A2(new_n690), .A3(new_n774), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n765), .A2(new_n760), .A3(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n736), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n731), .A2(new_n922), .A3(new_n773), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n253), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n509), .A2(new_n513), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT125), .Z(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(new_n233), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n648), .A2(G953), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n924), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n773), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT62), .ZN(new_n931));
  OR3_X1    g745(.A1(new_n671), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n931), .B1(new_n671), .B2(new_n930), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n661), .A2(new_n794), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n690), .A2(new_n935), .A3(new_n735), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n934), .A2(new_n760), .A3(new_n765), .A4(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(new_n927), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n937), .A2(new_n253), .A3(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n929), .A2(new_n939), .A3(KEYINPUT126), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n428), .B1(new_n938), .B2(KEYINPUT126), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n253), .B1(new_n941), .B2(G900), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n940), .B(new_n942), .Z(G72));
  NOR2_X1   g757(.A1(new_n937), .A2(new_n807), .ZN(new_n944));
  XNOR2_X1  g758(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n945));
  NAND2_X1  g759(.A1(G472), .A2(G902), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n666), .B1(new_n944), .B2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n552), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n921), .A2(new_n807), .A3(new_n923), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n949), .B1(new_n950), .B2(new_n947), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n948), .A2(new_n886), .A3(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n824), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n949), .A2(new_n666), .A3(new_n947), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(G57));
endmodule


