//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 1 1 0 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 0 0 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985;
  XOR2_X1   g000(.A(G15gat), .B(G43gat), .Z(new_n202));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT25), .ZN(new_n205));
  INV_X1    g004(.A(G169gat), .ZN(new_n206));
  INV_X1    g005(.A(G176gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n206), .A2(new_n207), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT23), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(G176gat), .ZN(new_n212));
  OR2_X1    g011(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NOR2_X1   g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216));
  INV_X1    g015(.A(G183gat), .ZN(new_n217));
  INV_X1    g016(.A(G190gat), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT24), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT24), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n220), .A2(G183gat), .A3(G190gat), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n216), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n223));
  OAI211_X1 g022(.A(new_n211), .B(new_n215), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n222), .A2(new_n223), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n205), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI211_X1 g027(.A(KEYINPUT66), .B(new_n205), .C1(new_n224), .C2(new_n225), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n205), .B1(new_n212), .B2(new_n206), .ZN(new_n230));
  OR2_X1    g029(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(G190gat), .ZN(new_n234));
  AND2_X1   g033(.A1(new_n219), .A2(new_n221), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n211), .B(new_n230), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n228), .A2(new_n229), .A3(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G127gat), .B(G134gat), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT72), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n238), .B(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT1), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(G113gat), .B2(G120gat), .ZN(new_n242));
  XOR2_X1   g041(.A(KEYINPUT71), .B(G113gat), .Z(new_n243));
  AOI21_X1  g042(.A(new_n242), .B1(new_n243), .B2(G120gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n240), .A2(new_n244), .ZN(new_n245));
  AND2_X1   g044(.A1(G113gat), .A2(G120gat), .ZN(new_n246));
  OR2_X1    g045(.A1(new_n242), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n238), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n245), .A2(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n208), .B1(new_n209), .B2(KEYINPUT26), .ZN(new_n251));
  OR2_X1    g050(.A1(new_n251), .A2(KEYINPUT70), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n208), .A2(KEYINPUT26), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n253), .B1(new_n251), .B2(KEYINPUT70), .ZN(new_n254));
  AOI22_X1  g053(.A1(new_n252), .A2(new_n254), .B1(G183gat), .B2(G190gat), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT27), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n256), .B1(new_n231), .B2(new_n232), .ZN(new_n257));
  NOR2_X1   g056(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n218), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  AND2_X1   g058(.A1(new_n259), .A2(KEYINPUT68), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT28), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n261), .B1(new_n259), .B2(KEYINPUT68), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT27), .B(G183gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n264), .A2(KEYINPUT28), .A3(new_n218), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(KEYINPUT69), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n255), .B1(new_n263), .B2(new_n266), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n237), .A2(new_n250), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n250), .B1(new_n237), .B2(new_n267), .ZN(new_n269));
  INV_X1    g068(.A(G227gat), .ZN(new_n270));
  INV_X1    g069(.A(G233gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NOR3_X1   g072(.A1(new_n268), .A2(new_n269), .A3(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n204), .B1(new_n274), .B2(KEYINPUT33), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n273), .B1(new_n268), .B2(new_n269), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT34), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT34), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n278), .B(new_n273), .C1(new_n268), .C2(new_n269), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n275), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n237), .A2(new_n267), .ZN(new_n281));
  AOI22_X1  g080(.A1(new_n240), .A2(new_n244), .B1(new_n247), .B2(new_n248), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n237), .A2(new_n267), .A3(new_n250), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(new_n272), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT32), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n204), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT33), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n288), .B1(new_n285), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n283), .A2(new_n284), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n278), .B1(new_n291), .B2(new_n273), .ZN(new_n292));
  INV_X1    g091(.A(new_n279), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n290), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AND3_X1   g093(.A1(new_n280), .A2(new_n287), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n287), .B1(new_n280), .B2(new_n294), .ZN(new_n296));
  XNOR2_X1  g095(.A(G78gat), .B(G106gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n297), .B(G22gat), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT31), .B(G50gat), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(G155gat), .A2(G162gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT2), .ZN(new_n303));
  INV_X1    g102(.A(G141gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G148gat), .ZN(new_n305));
  INV_X1    g104(.A(G148gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G141gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G155gat), .ZN(new_n309));
  INV_X1    g108(.A(G162gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AND3_X1   g110(.A1(new_n311), .A2(KEYINPUT78), .A3(new_n302), .ZN(new_n312));
  AOI21_X1  g111(.A(KEYINPUT78), .B1(new_n311), .B2(new_n302), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n303), .B(new_n308), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n308), .A2(new_n303), .ZN(new_n315));
  OR2_X1    g114(.A1(new_n302), .A2(KEYINPUT77), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n302), .A2(KEYINPUT77), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n315), .A2(new_n311), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT3), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n314), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT29), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT74), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT22), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n323), .A2(new_n324), .B1(G211gat), .B2(G218gat), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n325), .B1(new_n323), .B2(new_n324), .ZN(new_n326));
  XNOR2_X1  g125(.A(G197gat), .B(G204gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  XOR2_X1   g127(.A(G211gat), .B(G218gat), .Z(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n329), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n331), .A2(new_n326), .A3(new_n327), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n322), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT83), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n335), .B(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(G228gat), .A2(G233gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT80), .ZN(new_n339));
  AND3_X1   g138(.A1(new_n314), .A2(new_n318), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n339), .B1(new_n314), .B2(new_n318), .ZN(new_n341));
  OR2_X1    g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n332), .A2(KEYINPUT82), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n343), .A2(KEYINPUT29), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n330), .A2(KEYINPUT82), .A3(new_n332), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT3), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n337), .B(new_n338), .C1(new_n342), .C2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n314), .A2(new_n318), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT29), .B1(new_n330), .B2(new_n332), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n348), .B1(new_n349), .B2(KEYINPUT3), .ZN(new_n350));
  AOI22_X1  g149(.A1(new_n350), .A2(KEYINPUT84), .B1(new_n334), .B2(new_n322), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT84), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n352), .B(new_n348), .C1(new_n349), .C2(KEYINPUT3), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n338), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n301), .B1(new_n347), .B2(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n335), .B(KEYINPUT83), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n338), .B1(new_n346), .B2(new_n342), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NOR3_X1   g158(.A1(new_n359), .A2(new_n354), .A3(new_n300), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n299), .B1(new_n356), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n347), .A2(new_n355), .A3(new_n301), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n300), .B1(new_n359), .B2(new_n354), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n362), .A2(new_n363), .A3(new_n298), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  NOR3_X1   g164(.A1(new_n295), .A2(new_n296), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(G226gat), .A2(G233gat), .ZN(new_n367));
  XOR2_X1   g166(.A(new_n367), .B(KEYINPUT75), .Z(new_n368));
  NOR2_X1   g167(.A1(new_n368), .A2(KEYINPUT29), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n369), .B1(new_n237), .B2(new_n267), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n368), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n237), .A2(new_n267), .A3(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n371), .A2(new_n333), .A3(new_n373), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n237), .A2(new_n267), .A3(new_n372), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n334), .B1(new_n375), .B2(new_n370), .ZN(new_n376));
  XNOR2_X1  g175(.A(G8gat), .B(G36gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(G64gat), .B(G92gat), .ZN(new_n378));
  XOR2_X1   g177(.A(new_n377), .B(new_n378), .Z(new_n379));
  NAND3_X1  g178(.A1(new_n374), .A2(new_n376), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT76), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT30), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT30), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n380), .A2(KEYINPUT76), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n374), .A2(new_n376), .ZN(new_n385));
  INV_X1    g184(.A(new_n379), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n382), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  XOR2_X1   g187(.A(G1gat), .B(G29gat), .Z(new_n389));
  XNOR2_X1  g188(.A(new_n389), .B(KEYINPUT0), .ZN(new_n390));
  XNOR2_X1  g189(.A(G57gat), .B(G85gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n390), .B(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT5), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n250), .A2(new_n348), .ZN(new_n394));
  INV_X1    g193(.A(new_n348), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n282), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(G225gat), .A2(G233gat), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n393), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT79), .ZN(new_n401));
  AOI22_X1  g200(.A1(KEYINPUT3), .A2(new_n348), .B1(new_n245), .B2(new_n249), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n401), .B1(new_n402), .B2(new_n320), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n348), .A2(KEYINPUT3), .ZN(new_n404));
  AND4_X1   g203(.A1(new_n401), .A2(new_n404), .A3(new_n250), .A4(new_n320), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n398), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n342), .A2(KEYINPUT4), .A3(new_n282), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT4), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n396), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n400), .B1(new_n406), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n404), .A2(new_n250), .A3(new_n320), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT79), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n402), .A2(new_n401), .A3(new_n320), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n399), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT81), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n396), .A2(KEYINPUT4), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n408), .B(new_n282), .C1(new_n340), .C2(new_n341), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT5), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AND3_X1   g218(.A1(new_n415), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n416), .B1(new_n415), .B2(new_n419), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n392), .B(new_n411), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT6), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n417), .A2(new_n418), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n393), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT81), .B1(new_n406), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n415), .A2(new_n416), .A3(new_n419), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n392), .B1(new_n429), .B2(new_n411), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n424), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n411), .B1(new_n420), .B2(new_n421), .ZN(new_n432));
  INV_X1    g231(.A(new_n392), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n434), .A2(new_n423), .A3(new_n422), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n388), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n366), .A2(new_n436), .A3(KEYINPUT88), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT88), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n280), .A2(new_n294), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n286), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n280), .A2(new_n294), .A3(new_n287), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n361), .A2(new_n364), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  AOI22_X1  g242(.A1(new_n381), .A2(KEYINPUT30), .B1(new_n385), .B2(new_n386), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n424), .A2(new_n430), .ZN(new_n445));
  AOI211_X1 g244(.A(new_n423), .B(new_n392), .C1(new_n429), .C2(new_n411), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n384), .B(new_n444), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n438), .B1(new_n443), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n437), .A2(new_n448), .A3(KEYINPUT35), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT86), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n392), .B1(new_n450), .B2(KEYINPUT40), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n413), .A2(new_n414), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n398), .B1(new_n452), .B2(new_n425), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT39), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n451), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n394), .A2(new_n398), .A3(new_n396), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n413), .A2(new_n414), .B1(new_n417), .B2(new_n418), .ZN(new_n457));
  OAI211_X1 g256(.A(KEYINPUT39), .B(new_n456), .C1(new_n457), .C2(new_n398), .ZN(new_n458));
  NOR2_X1   g257(.A1(KEYINPUT85), .A2(KEYINPUT40), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n459), .A2(KEYINPUT86), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n455), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n460), .B1(new_n455), .B2(new_n458), .ZN(new_n462));
  NOR3_X1   g261(.A1(new_n461), .A2(new_n430), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n388), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT37), .ZN(new_n465));
  INV_X1    g264(.A(new_n376), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT87), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n333), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n465), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n374), .A2(new_n376), .A3(new_n467), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT38), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n386), .B1(new_n385), .B2(KEYINPUT37), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n465), .B1(new_n374), .B2(new_n376), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT38), .B1(new_n472), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n435), .A2(new_n431), .A3(new_n380), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n464), .B(new_n442), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n295), .A2(new_n296), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT36), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(KEYINPUT73), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(KEYINPUT73), .ZN(new_n483));
  OR2_X1    g282(.A1(new_n481), .A2(KEYINPUT73), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n483), .B(new_n484), .C1(new_n295), .C2(new_n296), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n447), .A2(new_n365), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n479), .A2(new_n482), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT35), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n438), .B(new_n488), .C1(new_n443), .C2(new_n447), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n449), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G15gat), .B(G22gat), .ZN(new_n491));
  INV_X1    g290(.A(G1gat), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(KEYINPUT16), .A3(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT91), .ZN(new_n494));
  INV_X1    g293(.A(G8gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n493), .B(new_n496), .C1(new_n492), .C2(new_n491), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n494), .A2(new_n495), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n497), .B(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(G29gat), .A2(G36gat), .ZN(new_n500));
  OR2_X1    g299(.A1(new_n500), .A2(KEYINPUT89), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(KEYINPUT89), .ZN(new_n502));
  NOR2_X1   g301(.A1(G29gat), .A2(G36gat), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT14), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n501), .A2(new_n502), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G43gat), .B(G50gat), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n507), .A2(KEYINPUT15), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n507), .A2(KEYINPUT15), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(new_n508), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n507), .A2(KEYINPUT15), .ZN(new_n513));
  OAI211_X1 g312(.A(KEYINPUT17), .B(new_n510), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n499), .A2(new_n514), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n507), .A2(KEYINPUT15), .A3(new_n509), .ZN(new_n516));
  INV_X1    g315(.A(new_n513), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n509), .B1(new_n507), .B2(KEYINPUT15), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR3_X1   g318(.A1(new_n519), .A2(KEYINPUT90), .A3(KEYINPUT17), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT90), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT17), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n515), .B1(new_n520), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(G229gat), .A2(G233gat), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n499), .A2(new_n519), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT18), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n525), .A2(KEYINPUT18), .A3(new_n526), .A4(new_n527), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n499), .A2(new_n519), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n526), .B(KEYINPUT13), .Z(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n530), .A2(new_n531), .A3(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G113gat), .B(G141gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(G197gat), .ZN(new_n538));
  XOR2_X1   g337(.A(KEYINPUT11), .B(G169gat), .Z(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(KEYINPUT12), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n536), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n530), .A2(new_n541), .A3(new_n531), .A4(new_n535), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AND2_X1   g344(.A1(new_n490), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(G85gat), .A2(G92gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(KEYINPUT7), .ZN(new_n548));
  NAND2_X1  g347(.A1(G99gat), .A2(G106gat), .ZN(new_n549));
  INV_X1    g348(.A(G85gat), .ZN(new_n550));
  INV_X1    g349(.A(G92gat), .ZN(new_n551));
  AOI22_X1  g350(.A1(KEYINPUT8), .A2(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G99gat), .B(G106gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n514), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(KEYINPUT90), .B1(new_n519), .B2(KEYINPUT17), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n522), .A2(new_n521), .A3(new_n523), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G190gat), .B(G218gat), .ZN(new_n561));
  AND2_X1   g360(.A1(G232gat), .A2(G233gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT41), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n563), .B1(new_n519), .B2(new_n556), .ZN(new_n564));
  OR3_X1    g363(.A1(new_n560), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n561), .B1(new_n560), .B2(new_n564), .ZN(new_n566));
  XNOR2_X1  g365(.A(G134gat), .B(G162gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(KEYINPUT96), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n562), .A2(KEYINPUT41), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n568), .B(new_n569), .Z(new_n570));
  AND4_X1   g369(.A1(KEYINPUT97), .A2(new_n565), .A3(new_n566), .A4(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT97), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n566), .A2(new_n572), .ZN(new_n573));
  AOI22_X1  g372(.A1(new_n573), .A2(new_n570), .B1(new_n565), .B2(new_n566), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(G71gat), .A2(G78gat), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT92), .ZN(new_n577));
  NAND2_X1  g376(.A1(G71gat), .A2(G78gat), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G57gat), .B(G64gat), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n577), .A2(KEYINPUT9), .ZN(new_n581));
  OAI221_X1 g380(.A(new_n579), .B1(new_n577), .B2(new_n578), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT95), .ZN(new_n583));
  INV_X1    g382(.A(G57gat), .ZN(new_n584));
  OAI21_X1  g383(.A(KEYINPUT93), .B1(new_n584), .B2(G64gat), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT93), .ZN(new_n586));
  INV_X1    g385(.A(G64gat), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(new_n587), .A3(G57gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n584), .A2(G64gat), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n585), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT94), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n585), .A2(new_n588), .A3(KEYINPUT94), .A4(new_n589), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n578), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n595), .B1(KEYINPUT9), .B2(new_n576), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n583), .B1(new_n594), .B2(new_n597), .ZN(new_n598));
  AOI211_X1 g397(.A(KEYINPUT95), .B(new_n596), .C1(new_n592), .C2(new_n593), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n582), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n601), .A2(KEYINPUT21), .ZN(new_n602));
  NAND2_X1  g401(.A1(G231gat), .A2(G233gat), .ZN(new_n603));
  OR2_X1    g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n603), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(G127gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n601), .A2(KEYINPUT21), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(new_n499), .ZN(new_n609));
  INV_X1    g408(.A(G127gat), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n604), .A2(new_n610), .A3(new_n605), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n607), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n609), .B1(new_n607), .B2(new_n611), .ZN(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(new_n309), .ZN(new_n616));
  XNOR2_X1  g415(.A(G183gat), .B(G211gat), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n616), .B(new_n617), .Z(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  OR3_X1    g418(.A1(new_n613), .A2(new_n614), .A3(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n619), .B1(new_n613), .B2(new_n614), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n575), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n600), .A2(new_n556), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT10), .ZN(new_n624));
  OAI211_X1 g423(.A(new_n555), .B(new_n582), .C1(new_n598), .C2(new_n599), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n625), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(KEYINPUT10), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G230gat), .A2(G233gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n623), .A2(new_n625), .ZN(new_n632));
  INV_X1    g431(.A(new_n630), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G120gat), .B(G148gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(G176gat), .B(G204gat), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n635), .B(new_n636), .Z(new_n637));
  NAND3_X1  g436(.A1(new_n631), .A2(new_n634), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n630), .B(KEYINPUT98), .Z(new_n640));
  AOI21_X1  g439(.A(new_n640), .B1(new_n626), .B2(new_n628), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n637), .B1(new_n642), .B2(new_n634), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n622), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n546), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n445), .A2(new_n446), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g449(.A1(new_n647), .A2(new_n388), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT16), .B(G8gat), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(KEYINPUT99), .B1(new_n653), .B2(KEYINPUT42), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT99), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT42), .ZN(new_n656));
  OAI211_X1 g455(.A(new_n655), .B(new_n656), .C1(new_n651), .C2(new_n652), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  AOI22_X1  g457(.A1(new_n653), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n651), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(G1325gat));
  NAND2_X1  g459(.A1(new_n482), .A2(new_n485), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n647), .A2(G15gat), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n546), .A2(new_n480), .A3(new_n646), .ZN(new_n663));
  INV_X1    g462(.A(G15gat), .ZN(new_n664));
  AND3_X1   g463(.A1(new_n663), .A2(KEYINPUT100), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(KEYINPUT100), .B1(new_n663), .B2(new_n664), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n662), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT101), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1326gat));
  NAND3_X1  g468(.A1(new_n546), .A2(new_n365), .A3(new_n646), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT43), .B(G22gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(G1327gat));
  NAND2_X1  g471(.A1(new_n620), .A2(new_n621), .ZN(new_n673));
  INV_X1    g472(.A(new_n575), .ZN(new_n674));
  INV_X1    g473(.A(new_n644), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n546), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n648), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n677), .A2(G29gat), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n679), .B(KEYINPUT45), .Z(new_n680));
  NAND2_X1  g479(.A1(new_n490), .A2(new_n575), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n682), .A2(KEYINPUT44), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n490), .A2(new_n575), .A3(new_n685), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n620), .A2(KEYINPUT102), .A3(new_n621), .ZN(new_n688));
  AOI21_X1  g487(.A(KEYINPUT102), .B1(new_n620), .B2(new_n621), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n545), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n691), .A2(new_n692), .A3(new_n675), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n687), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(KEYINPUT104), .B1(new_n694), .B2(new_n678), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(G29gat), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n694), .A2(KEYINPUT104), .A3(new_n678), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n680), .B1(new_n696), .B2(new_n697), .ZN(G1328gat));
  INV_X1    g497(.A(new_n388), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n677), .A2(G36gat), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT46), .ZN(new_n701));
  OAI21_X1  g500(.A(G36gat), .B1(new_n694), .B2(new_n699), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(G1329gat));
  INV_X1    g502(.A(new_n480), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n677), .A2(G43gat), .A3(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n687), .A2(new_n661), .A3(new_n693), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n705), .B1(new_n706), .B2(G43gat), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g507(.A1(new_n684), .A2(new_n365), .A3(new_n686), .A4(new_n693), .ZN(new_n709));
  AOI21_X1  g508(.A(KEYINPUT105), .B1(new_n709), .B2(G50gat), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT48), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(G50gat), .ZN(new_n713));
  AND4_X1   g512(.A1(new_n713), .A2(new_n546), .A3(new_n365), .A4(new_n676), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n714), .B1(G50gat), .B2(new_n709), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n712), .B(new_n715), .ZN(G1331gat));
  NOR2_X1   g515(.A1(new_n545), .A2(new_n644), .ZN(new_n717));
  AND3_X1   g516(.A1(new_n490), .A2(new_n622), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n648), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n388), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n721), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n722));
  XOR2_X1   g521(.A(KEYINPUT49), .B(G64gat), .Z(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(new_n721), .B2(new_n723), .ZN(G1333gat));
  NAND2_X1  g523(.A1(new_n718), .A2(new_n480), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT106), .ZN(new_n726));
  AOI21_X1  g525(.A(G71gat), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n727), .B1(new_n726), .B2(new_n725), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n718), .A2(G71gat), .A3(new_n661), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n728), .A2(new_n729), .A3(new_n731), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(G1334gat));
  NAND2_X1  g534(.A1(new_n718), .A2(new_n365), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g536(.A1(new_n673), .A2(new_n545), .A3(new_n644), .ZN(new_n738));
  AND3_X1   g537(.A1(new_n684), .A2(new_n686), .A3(new_n738), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n739), .A2(new_n648), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n673), .A2(new_n545), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n490), .A2(new_n575), .A3(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT51), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n490), .A2(KEYINPUT51), .A3(new_n575), .A4(new_n741), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n648), .A2(new_n550), .A3(new_n675), .ZN(new_n748));
  OAI22_X1  g547(.A1(new_n740), .A2(new_n550), .B1(new_n747), .B2(new_n748), .ZN(G1336gat));
  NAND4_X1  g548(.A1(new_n684), .A2(new_n388), .A3(new_n686), .A4(new_n738), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n750), .A2(G92gat), .ZN(new_n751));
  AND3_X1   g550(.A1(new_n742), .A2(KEYINPUT108), .A3(KEYINPUT51), .ZN(new_n752));
  AOI21_X1  g551(.A(KEYINPUT51), .B1(new_n742), .B2(KEYINPUT108), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n699), .A2(G92gat), .A3(new_n644), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n752), .A2(new_n753), .A3(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(KEYINPUT52), .B1(new_n751), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT110), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n750), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n750), .A2(new_n758), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n759), .A2(new_n760), .A3(new_n551), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n755), .B1(new_n744), .B2(new_n745), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT109), .ZN(new_n763));
  AOI21_X1  g562(.A(KEYINPUT52), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(new_n763), .B2(new_n762), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n757), .B1(new_n761), .B2(new_n765), .ZN(G1337gat));
  NAND2_X1  g565(.A1(new_n739), .A2(new_n661), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(G99gat), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n704), .A2(G99gat), .A3(new_n644), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n746), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT111), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n768), .A2(KEYINPUT111), .A3(new_n770), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(G1338gat));
  NAND4_X1  g574(.A1(new_n684), .A2(new_n365), .A3(new_n686), .A4(new_n738), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(G106gat), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT53), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n442), .A2(G106gat), .A3(new_n644), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n746), .A2(new_n779), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n777), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n742), .A2(KEYINPUT108), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n743), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n742), .A2(KEYINPUT108), .A3(KEYINPUT51), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n783), .A2(new_n784), .A3(new_n779), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n778), .B1(new_n785), .B2(new_n777), .ZN(new_n786));
  OAI21_X1  g585(.A(KEYINPUT112), .B1(new_n781), .B2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT112), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n777), .A2(new_n778), .A3(new_n780), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n752), .A2(new_n753), .ZN(new_n790));
  AOI22_X1  g589(.A1(new_n790), .A2(new_n779), .B1(G106gat), .B2(new_n776), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n788), .B(new_n789), .C1(new_n791), .C2(new_n778), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n787), .A2(new_n792), .ZN(G1339gat));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT54), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n637), .B1(new_n641), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n633), .B1(new_n626), .B2(new_n628), .ZN(new_n797));
  AND3_X1   g596(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n640), .B1(new_n625), .B2(new_n624), .ZN(new_n799));
  OAI21_X1  g598(.A(KEYINPUT54), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n796), .B1(new_n797), .B2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT55), .B1(new_n800), .B2(new_n797), .ZN(new_n804));
  INV_X1    g603(.A(new_n640), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n629), .A2(new_n795), .A3(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n637), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n804), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n799), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n795), .B1(new_n811), .B2(new_n626), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n802), .B1(new_n631), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT113), .B1(new_n813), .B2(new_n796), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n638), .B(new_n803), .C1(new_n810), .C2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n809), .B1(new_n804), .B2(new_n808), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n813), .A2(KEYINPUT113), .A3(new_n796), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n639), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n820), .A2(KEYINPUT114), .A3(new_n803), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n817), .A2(new_n545), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n526), .B1(new_n525), .B2(new_n527), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n533), .A2(new_n534), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n540), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n544), .A2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n675), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n575), .B1(new_n822), .B2(new_n828), .ZN(new_n829));
  AND4_X1   g628(.A1(new_n575), .A2(new_n817), .A3(new_n827), .A4(new_n821), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n690), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n622), .A2(new_n692), .A3(new_n644), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n794), .B1(new_n833), .B2(new_n442), .ZN(new_n834));
  AOI211_X1 g633(.A(KEYINPUT115), .B(new_n365), .C1(new_n831), .C2(new_n832), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n678), .A2(new_n388), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n838), .A2(new_n704), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(G113gat), .B1(new_n840), .B2(new_n692), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n842));
  AND4_X1   g641(.A1(new_n842), .A2(new_n833), .A3(new_n648), .A4(new_n366), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n678), .B1(new_n831), .B2(new_n832), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n842), .B1(new_n844), .B2(new_n366), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n699), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n692), .A2(new_n243), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(KEYINPUT117), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n841), .B1(new_n846), .B2(new_n848), .ZN(G1340gat));
  OAI21_X1  g648(.A(G120gat), .B1(new_n840), .B2(new_n644), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n644), .A2(G120gat), .ZN(new_n851));
  XOR2_X1   g650(.A(new_n851), .B(KEYINPUT118), .Z(new_n852));
  OAI21_X1  g651(.A(new_n850), .B1(new_n846), .B2(new_n852), .ZN(G1341gat));
  OAI21_X1  g652(.A(G127gat), .B1(new_n840), .B2(new_n690), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n673), .A2(new_n610), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n854), .B1(new_n846), .B2(new_n855), .ZN(G1342gat));
  NOR3_X1   g655(.A1(new_n388), .A2(new_n674), .A3(G134gat), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n857), .B1(new_n843), .B2(new_n845), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT56), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT56), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n860), .B(new_n857), .C1(new_n843), .C2(new_n845), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n575), .B(new_n839), .C1(new_n834), .C2(new_n835), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(G134gat), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n859), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(KEYINPUT119), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n859), .A2(new_n866), .A3(new_n861), .A4(new_n863), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(G1343gat));
  NOR2_X1   g667(.A1(new_n661), .A2(new_n838), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT57), .B1(new_n833), .B2(new_n365), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n442), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n673), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT120), .ZN(new_n875));
  AOI22_X1  g674(.A1(new_n543), .A2(new_n544), .B1(new_n801), .B2(new_n802), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n638), .B1(new_n810), .B2(new_n814), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n875), .B(new_n828), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n674), .ZN(new_n880));
  AOI22_X1  g679(.A1(new_n820), .A2(new_n876), .B1(new_n675), .B2(new_n827), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n881), .A2(new_n875), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n874), .B1(new_n883), .B2(new_n830), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n873), .B1(new_n884), .B2(new_n832), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n545), .B(new_n869), .C1(new_n870), .C2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(G141gat), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n661), .A2(new_n388), .A3(new_n442), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n844), .A2(new_n304), .A3(new_n545), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n890), .B(KEYINPUT58), .ZN(G1344gat));
  AOI21_X1  g690(.A(new_n575), .B1(new_n881), .B2(new_n875), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n828), .B1(new_n877), .B2(new_n878), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(KEYINPUT120), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n820), .A2(new_n575), .A3(new_n803), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n826), .B1(new_n895), .B2(KEYINPUT121), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n820), .A2(new_n897), .A3(new_n575), .A4(new_n803), .ZN(new_n898));
  AOI22_X1  g697(.A1(new_n892), .A2(new_n894), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n832), .B1(new_n899), .B2(new_n673), .ZN(new_n900));
  AOI21_X1  g699(.A(KEYINPUT57), .B1(new_n900), .B2(new_n365), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n873), .B1(new_n831), .B2(new_n832), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n869), .A2(new_n675), .ZN(new_n904));
  OAI211_X1 g703(.A(KEYINPUT59), .B(G148gat), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n844), .A2(new_n675), .A3(new_n888), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n906), .A2(KEYINPUT59), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n869), .B1(new_n870), .B2(new_n885), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n644), .A2(KEYINPUT59), .ZN(new_n909));
  OAI221_X1 g708(.A(new_n905), .B1(G148gat), .B2(new_n907), .C1(new_n908), .C2(new_n909), .ZN(G1345gat));
  OAI21_X1  g709(.A(G155gat), .B1(new_n908), .B2(new_n690), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n844), .A2(new_n309), .A3(new_n673), .A4(new_n888), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1346gat));
  OAI21_X1  g712(.A(G162gat), .B1(new_n908), .B2(new_n674), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n844), .A2(new_n310), .A3(new_n575), .A4(new_n888), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1347gat));
  NOR3_X1   g715(.A1(new_n704), .A2(new_n648), .A3(new_n699), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n545), .B(new_n917), .C1(new_n834), .C2(new_n835), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(G169gat), .ZN(new_n919));
  AND4_X1   g718(.A1(new_n678), .A2(new_n833), .A3(new_n388), .A4(new_n366), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n920), .A2(new_n545), .A3(new_n213), .A4(new_n214), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT122), .ZN(G1348gat));
  OAI211_X1 g722(.A(new_n675), .B(new_n917), .C1(new_n834), .C2(new_n835), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(G176gat), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n920), .A2(new_n207), .A3(new_n675), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n927), .B(new_n928), .ZN(G1349gat));
  OAI211_X1 g728(.A(new_n691), .B(new_n917), .C1(new_n834), .C2(new_n835), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n233), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n920), .A2(new_n264), .A3(new_n673), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g733(.A1(new_n920), .A2(new_n218), .A3(new_n575), .ZN(new_n935));
  XOR2_X1   g734(.A(new_n935), .B(KEYINPUT124), .Z(new_n936));
  OAI211_X1 g735(.A(new_n575), .B(new_n917), .C1(new_n834), .C2(new_n835), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n937), .A2(KEYINPUT61), .A3(G190gat), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n939));
  INV_X1    g738(.A(new_n937), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n940), .B2(new_n218), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n936), .A2(new_n938), .A3(new_n941), .ZN(G1351gat));
  XNOR2_X1  g741(.A(KEYINPUT125), .B(G197gat), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n648), .A2(new_n699), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n482), .A2(new_n485), .A3(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(new_n832), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n895), .A2(KEYINPUT121), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n947), .A2(new_n827), .A3(new_n898), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n948), .B1(new_n880), .B2(new_n882), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n946), .B1(new_n949), .B2(new_n874), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n871), .B1(new_n950), .B2(new_n442), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n833), .A2(new_n872), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n945), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n943), .B1(new_n953), .B2(new_n545), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n648), .B1(new_n831), .B2(new_n832), .ZN(new_n955));
  NOR3_X1   g754(.A1(new_n661), .A2(new_n699), .A3(new_n442), .ZN(new_n956));
  AND4_X1   g755(.A1(new_n545), .A2(new_n955), .A3(new_n943), .A4(new_n956), .ZN(new_n957));
  OR2_X1    g756(.A1(new_n954), .A2(new_n957), .ZN(G1352gat));
  INV_X1    g757(.A(new_n953), .ZN(new_n959));
  OAI21_X1  g758(.A(G204gat), .B1(new_n959), .B2(new_n644), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n644), .A2(G204gat), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n955), .A2(new_n956), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(KEYINPUT62), .ZN(new_n963));
  OR2_X1    g762(.A1(new_n962), .A2(KEYINPUT62), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n960), .A2(new_n963), .A3(new_n964), .ZN(G1353gat));
  INV_X1    g764(.A(KEYINPUT63), .ZN(new_n966));
  INV_X1    g765(.A(new_n945), .ZN(new_n967));
  OAI211_X1 g766(.A(new_n673), .B(new_n967), .C1(new_n901), .C2(new_n902), .ZN(new_n968));
  OAI21_X1  g767(.A(G211gat), .B1(new_n968), .B2(KEYINPUT126), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT126), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n970), .B1(new_n953), .B2(new_n673), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n966), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n968), .A2(KEYINPUT126), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n953), .A2(new_n970), .A3(new_n673), .ZN(new_n974));
  NAND4_X1  g773(.A1(new_n973), .A2(new_n974), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n874), .A2(G211gat), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n955), .A2(new_n956), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n976), .A2(new_n978), .ZN(G1354gat));
  NAND2_X1  g778(.A1(new_n953), .A2(KEYINPUT127), .ZN(new_n980));
  INV_X1    g779(.A(new_n980), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n575), .B1(new_n953), .B2(KEYINPUT127), .ZN(new_n982));
  OAI21_X1  g781(.A(G218gat), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n674), .A2(G218gat), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n955), .A2(new_n956), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n983), .A2(new_n985), .ZN(G1355gat));
endmodule


