

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U323 ( .A(n410), .B(n409), .ZN(n564) );
  XNOR2_X1 U324 ( .A(KEYINPUT111), .B(KEYINPUT46), .ZN(n384) );
  XNOR2_X1 U325 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U326 ( .A(n389), .B(KEYINPUT47), .ZN(n390) );
  XNOR2_X1 U327 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U328 ( .A(KEYINPUT54), .B(KEYINPUT123), .ZN(n409) );
  XNOR2_X1 U329 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U330 ( .A(n303), .B(n302), .ZN(n364) );
  XOR2_X1 U331 ( .A(n395), .B(n322), .Z(n525) );
  XNOR2_X1 U332 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U333 ( .A(n456), .B(n455), .ZN(G1349GAT) );
  XOR2_X1 U334 ( .A(KEYINPUT32), .B(KEYINPUT70), .Z(n292) );
  NAND2_X1 U335 ( .A1(G230GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U336 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U337 ( .A(n293), .B(KEYINPUT33), .Z(n298) );
  XOR2_X1 U338 ( .A(G64GAT), .B(G92GAT), .Z(n295) );
  XNOR2_X1 U339 ( .A(G176GAT), .B(G204GAT), .ZN(n294) );
  XNOR2_X1 U340 ( .A(n295), .B(n294), .ZN(n396) );
  XNOR2_X1 U341 ( .A(G106GAT), .B(G78GAT), .ZN(n296) );
  XNOR2_X1 U342 ( .A(n296), .B(G148GAT), .ZN(n446) );
  XNOR2_X1 U343 ( .A(n396), .B(n446), .ZN(n297) );
  XNOR2_X1 U344 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U345 ( .A(KEYINPUT31), .B(n299), .Z(n303) );
  XOR2_X1 U346 ( .A(G120GAT), .B(G71GAT), .Z(n310) );
  XOR2_X1 U347 ( .A(G99GAT), .B(G85GAT), .Z(n353) );
  XNOR2_X1 U348 ( .A(n310), .B(n353), .ZN(n301) );
  XOR2_X1 U349 ( .A(KEYINPUT13), .B(G57GAT), .Z(n329) );
  XNOR2_X1 U350 ( .A(n329), .B(KEYINPUT71), .ZN(n300) );
  INV_X1 U351 ( .A(n364), .ZN(n574) );
  XNOR2_X1 U352 ( .A(KEYINPUT41), .B(n574), .ZN(n548) );
  XOR2_X1 U353 ( .A(n548), .B(KEYINPUT103), .Z(n529) );
  XOR2_X1 U354 ( .A(KEYINPUT83), .B(G183GAT), .Z(n305) );
  XNOR2_X1 U355 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n304) );
  XNOR2_X1 U356 ( .A(n305), .B(n304), .ZN(n307) );
  XOR2_X1 U357 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n306) );
  XNOR2_X1 U358 ( .A(n307), .B(n306), .ZN(n395) );
  XOR2_X1 U359 ( .A(KEYINPUT20), .B(KEYINPUT85), .Z(n309) );
  XNOR2_X1 U360 ( .A(KEYINPUT84), .B(KEYINPUT82), .ZN(n308) );
  XNOR2_X1 U361 ( .A(n309), .B(n308), .ZN(n321) );
  XOR2_X1 U362 ( .A(G190GAT), .B(G99GAT), .Z(n312) );
  XOR2_X1 U363 ( .A(G15GAT), .B(G127GAT), .Z(n330) );
  XNOR2_X1 U364 ( .A(n330), .B(n310), .ZN(n311) );
  XNOR2_X1 U365 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U366 ( .A(n313), .B(KEYINPUT81), .Z(n319) );
  XNOR2_X1 U367 ( .A(G113GAT), .B(G134GAT), .ZN(n314) );
  XNOR2_X1 U368 ( .A(n314), .B(KEYINPUT0), .ZN(n429) );
  XOR2_X1 U369 ( .A(n429), .B(G176GAT), .Z(n316) );
  NAND2_X1 U370 ( .A1(G227GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U371 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U372 ( .A(G43GAT), .B(n317), .ZN(n318) );
  XNOR2_X1 U373 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U374 ( .A(n321), .B(n320), .Z(n322) );
  INV_X1 U375 ( .A(n525), .ZN(n466) );
  XOR2_X1 U376 ( .A(KEYINPUT15), .B(KEYINPUT79), .Z(n324) );
  XNOR2_X1 U377 ( .A(G64GAT), .B(KEYINPUT80), .ZN(n323) );
  XNOR2_X1 U378 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U379 ( .A(KEYINPUT78), .B(KEYINPUT77), .Z(n326) );
  XNOR2_X1 U380 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n325) );
  XNOR2_X1 U381 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U382 ( .A(n328), .B(n327), .ZN(n342) );
  XOR2_X1 U383 ( .A(n329), .B(G78GAT), .Z(n332) );
  XNOR2_X1 U384 ( .A(n330), .B(G211GAT), .ZN(n331) );
  XNOR2_X1 U385 ( .A(n332), .B(n331), .ZN(n338) );
  XOR2_X1 U386 ( .A(G22GAT), .B(G155GAT), .Z(n435) );
  XOR2_X1 U387 ( .A(G1GAT), .B(KEYINPUT68), .Z(n334) );
  XNOR2_X1 U388 ( .A(G8GAT), .B(KEYINPUT69), .ZN(n333) );
  XNOR2_X1 U389 ( .A(n334), .B(n333), .ZN(n371) );
  XOR2_X1 U390 ( .A(n435), .B(n371), .Z(n336) );
  NAND2_X1 U391 ( .A1(G231GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U392 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U393 ( .A(n338), .B(n337), .Z(n340) );
  XNOR2_X1 U394 ( .A(G183GAT), .B(G71GAT), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U396 ( .A(n342), .B(n341), .ZN(n577) );
  XOR2_X1 U397 ( .A(KEYINPUT9), .B(G92GAT), .Z(n344) );
  XNOR2_X1 U398 ( .A(G134GAT), .B(G106GAT), .ZN(n343) );
  XNOR2_X1 U399 ( .A(n344), .B(n343), .ZN(n361) );
  XOR2_X1 U400 ( .A(KEYINPUT73), .B(KEYINPUT76), .Z(n346) );
  NAND2_X1 U401 ( .A1(G232GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U402 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U403 ( .A(n347), .B(KEYINPUT11), .Z(n352) );
  XOR2_X1 U404 ( .A(G29GAT), .B(G43GAT), .Z(n349) );
  XNOR2_X1 U405 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n348) );
  XNOR2_X1 U406 ( .A(n349), .B(n348), .ZN(n372) );
  XNOR2_X1 U407 ( .A(G50GAT), .B(KEYINPUT72), .ZN(n350) );
  XNOR2_X1 U408 ( .A(n350), .B(G162GAT), .ZN(n439) );
  XNOR2_X1 U409 ( .A(n372), .B(n439), .ZN(n351) );
  XNOR2_X1 U410 ( .A(n352), .B(n351), .ZN(n357) );
  XOR2_X1 U411 ( .A(KEYINPUT75), .B(KEYINPUT10), .Z(n355) );
  XOR2_X1 U412 ( .A(G36GAT), .B(G190GAT), .Z(n403) );
  XNOR2_X1 U413 ( .A(n353), .B(n403), .ZN(n354) );
  XNOR2_X1 U414 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U415 ( .A(n357), .B(n356), .Z(n359) );
  XNOR2_X1 U416 ( .A(G218GAT), .B(KEYINPUT74), .ZN(n358) );
  XNOR2_X1 U417 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U418 ( .A(n361), .B(n360), .Z(n537) );
  XNOR2_X1 U419 ( .A(KEYINPUT36), .B(n537), .ZN(n580) );
  NOR2_X1 U420 ( .A1(n577), .A2(n580), .ZN(n362) );
  XOR2_X1 U421 ( .A(KEYINPUT45), .B(n362), .Z(n363) );
  NOR2_X1 U422 ( .A1(n364), .A2(n363), .ZN(n383) );
  XOR2_X1 U423 ( .A(KEYINPUT66), .B(KEYINPUT67), .Z(n366) );
  XNOR2_X1 U424 ( .A(G169GAT), .B(G15GAT), .ZN(n365) );
  XNOR2_X1 U425 ( .A(n366), .B(n365), .ZN(n382) );
  XOR2_X1 U426 ( .A(G113GAT), .B(G141GAT), .Z(n368) );
  XNOR2_X1 U427 ( .A(G197GAT), .B(G22GAT), .ZN(n367) );
  XNOR2_X1 U428 ( .A(n368), .B(n367), .ZN(n370) );
  XOR2_X1 U429 ( .A(G36GAT), .B(G50GAT), .Z(n369) );
  XNOR2_X1 U430 ( .A(n370), .B(n369), .ZN(n378) );
  XNOR2_X1 U431 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U432 ( .A(KEYINPUT64), .B(KEYINPUT65), .Z(n374) );
  XNOR2_X1 U433 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n373) );
  XNOR2_X1 U434 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U435 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U436 ( .A(n378), .B(n377), .ZN(n380) );
  NAND2_X1 U437 ( .A1(G229GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U438 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U439 ( .A(n382), .B(n381), .Z(n568) );
  NAND2_X1 U440 ( .A1(n383), .A2(n568), .ZN(n393) );
  INV_X1 U441 ( .A(n577), .ZN(n558) );
  INV_X1 U442 ( .A(n568), .ZN(n556) );
  NAND2_X1 U443 ( .A1(n556), .A2(n548), .ZN(n385) );
  NOR2_X1 U444 ( .A1(n558), .A2(n386), .ZN(n387) );
  XNOR2_X1 U445 ( .A(n387), .B(KEYINPUT112), .ZN(n388) );
  NAND2_X1 U446 ( .A1(n388), .A2(n537), .ZN(n391) );
  XNOR2_X1 U447 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n389) );
  NAND2_X1 U448 ( .A1(n393), .A2(n392), .ZN(n394) );
  XNOR2_X1 U449 ( .A(n394), .B(KEYINPUT48), .ZN(n522) );
  INV_X1 U450 ( .A(n395), .ZN(n397) );
  XNOR2_X1 U451 ( .A(n397), .B(n396), .ZN(n407) );
  XOR2_X1 U452 ( .A(G211GAT), .B(KEYINPUT21), .Z(n399) );
  XNOR2_X1 U453 ( .A(G197GAT), .B(G218GAT), .ZN(n398) );
  XNOR2_X1 U454 ( .A(n399), .B(n398), .ZN(n447) );
  XOR2_X1 U455 ( .A(n447), .B(KEYINPUT94), .Z(n401) );
  NAND2_X1 U456 ( .A1(G226GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U457 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U458 ( .A(n402), .B(KEYINPUT95), .Z(n405) );
  XNOR2_X1 U459 ( .A(G8GAT), .B(n403), .ZN(n404) );
  XNOR2_X1 U460 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U461 ( .A(n407), .B(n406), .ZN(n514) );
  XNOR2_X1 U462 ( .A(KEYINPUT122), .B(n514), .ZN(n408) );
  NAND2_X1 U463 ( .A1(n522), .A2(n408), .ZN(n410) );
  XOR2_X1 U464 ( .A(KEYINPUT91), .B(KEYINPUT1), .Z(n412) );
  XNOR2_X1 U465 ( .A(G57GAT), .B(KEYINPUT90), .ZN(n411) );
  XNOR2_X1 U466 ( .A(n412), .B(n411), .ZN(n416) );
  XOR2_X1 U467 ( .A(KEYINPUT5), .B(KEYINPUT88), .Z(n414) );
  XNOR2_X1 U468 ( .A(KEYINPUT89), .B(KEYINPUT6), .ZN(n413) );
  XNOR2_X1 U469 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U470 ( .A(n416), .B(n415), .Z(n421) );
  XOR2_X1 U471 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n418) );
  NAND2_X1 U472 ( .A1(G225GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U473 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U474 ( .A(KEYINPUT4), .B(n419), .ZN(n420) );
  XNOR2_X1 U475 ( .A(n421), .B(n420), .ZN(n433) );
  XOR2_X1 U476 ( .A(G85GAT), .B(G155GAT), .Z(n423) );
  XNOR2_X1 U477 ( .A(G29GAT), .B(G162GAT), .ZN(n422) );
  XNOR2_X1 U478 ( .A(n423), .B(n422), .ZN(n427) );
  XOR2_X1 U479 ( .A(G148GAT), .B(G120GAT), .Z(n425) );
  XNOR2_X1 U480 ( .A(G1GAT), .B(G127GAT), .ZN(n424) );
  XNOR2_X1 U481 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U482 ( .A(n427), .B(n426), .Z(n431) );
  XNOR2_X1 U483 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n428) );
  XNOR2_X1 U484 ( .A(n428), .B(KEYINPUT2), .ZN(n434) );
  XNOR2_X1 U485 ( .A(n429), .B(n434), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U487 ( .A(n433), .B(n432), .ZN(n543) );
  INV_X1 U488 ( .A(n543), .ZN(n565) );
  XOR2_X1 U489 ( .A(n435), .B(n434), .Z(n437) );
  NAND2_X1 U490 ( .A1(G228GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U492 ( .A(n438), .B(G204GAT), .Z(n441) );
  XNOR2_X1 U493 ( .A(n439), .B(KEYINPUT22), .ZN(n440) );
  XNOR2_X1 U494 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U495 ( .A(KEYINPUT86), .B(KEYINPUT24), .Z(n443) );
  XNOR2_X1 U496 ( .A(KEYINPUT23), .B(KEYINPUT87), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U498 ( .A(n445), .B(n444), .Z(n449) );
  XNOR2_X1 U499 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U500 ( .A(n449), .B(n448), .ZN(n465) );
  AND2_X1 U501 ( .A1(n565), .A2(n465), .ZN(n450) );
  AND2_X1 U502 ( .A1(n564), .A2(n450), .ZN(n451) );
  XNOR2_X1 U503 ( .A(n451), .B(KEYINPUT55), .ZN(n452) );
  NOR2_X1 U504 ( .A1(n466), .A2(n452), .ZN(n561) );
  NAND2_X1 U505 ( .A1(n529), .A2(n561), .ZN(n456) );
  XOR2_X1 U506 ( .A(G176GAT), .B(KEYINPUT56), .Z(n454) );
  XNOR2_X1 U507 ( .A(KEYINPUT124), .B(KEYINPUT57), .ZN(n453) );
  XNOR2_X1 U508 ( .A(KEYINPUT100), .B(KEYINPUT101), .ZN(n477) );
  XOR2_X1 U509 ( .A(G1GAT), .B(KEYINPUT34), .Z(n475) );
  NAND2_X1 U510 ( .A1(n514), .A2(n525), .ZN(n457) );
  NAND2_X1 U511 ( .A1(n465), .A2(n457), .ZN(n458) );
  XOR2_X1 U512 ( .A(KEYINPUT25), .B(n458), .Z(n462) );
  XNOR2_X1 U513 ( .A(n514), .B(KEYINPUT96), .ZN(n459) );
  XNOR2_X1 U514 ( .A(n459), .B(KEYINPUT27), .ZN(n523) );
  NOR2_X1 U515 ( .A1(n525), .A2(n465), .ZN(n460) );
  XNOR2_X1 U516 ( .A(n460), .B(KEYINPUT26), .ZN(n566) );
  NAND2_X1 U517 ( .A1(n523), .A2(n566), .ZN(n461) );
  NAND2_X1 U518 ( .A1(n462), .A2(n461), .ZN(n463) );
  XNOR2_X1 U519 ( .A(KEYINPUT97), .B(n463), .ZN(n464) );
  NOR2_X1 U520 ( .A1(n543), .A2(n464), .ZN(n469) );
  XNOR2_X1 U521 ( .A(n465), .B(KEYINPUT28), .ZN(n481) );
  NAND2_X1 U522 ( .A1(n543), .A2(n481), .ZN(n524) );
  NAND2_X1 U523 ( .A1(n523), .A2(n466), .ZN(n467) );
  NOR2_X1 U524 ( .A1(n524), .A2(n467), .ZN(n468) );
  NOR2_X1 U525 ( .A1(n469), .A2(n468), .ZN(n484) );
  INV_X1 U526 ( .A(n537), .ZN(n560) );
  NOR2_X1 U527 ( .A1(n577), .A2(n560), .ZN(n470) );
  XOR2_X1 U528 ( .A(KEYINPUT16), .B(n470), .Z(n471) );
  NOR2_X1 U529 ( .A1(n484), .A2(n471), .ZN(n472) );
  XOR2_X1 U530 ( .A(KEYINPUT98), .B(n472), .Z(n497) );
  NAND2_X1 U531 ( .A1(n556), .A2(n574), .ZN(n487) );
  NOR2_X1 U532 ( .A1(n497), .A2(n487), .ZN(n473) );
  XOR2_X1 U533 ( .A(KEYINPUT99), .B(n473), .Z(n482) );
  NAND2_X1 U534 ( .A1(n482), .A2(n543), .ZN(n474) );
  XNOR2_X1 U535 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n477), .B(n476), .ZN(G1324GAT) );
  NAND2_X1 U537 ( .A1(n482), .A2(n514), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n478), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U539 ( .A(G15GAT), .B(KEYINPUT35), .Z(n480) );
  NAND2_X1 U540 ( .A1(n482), .A2(n525), .ZN(n479) );
  XNOR2_X1 U541 ( .A(n480), .B(n479), .ZN(G1326GAT) );
  INV_X1 U542 ( .A(n481), .ZN(n518) );
  NAND2_X1 U543 ( .A1(n482), .A2(n518), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n483), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U545 ( .A(KEYINPUT102), .B(KEYINPUT39), .Z(n490) );
  NOR2_X1 U546 ( .A1(n484), .A2(n580), .ZN(n485) );
  NAND2_X1 U547 ( .A1(n485), .A2(n577), .ZN(n486) );
  XOR2_X1 U548 ( .A(KEYINPUT37), .B(n486), .Z(n510) );
  NOR2_X1 U549 ( .A1(n510), .A2(n487), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n488), .B(KEYINPUT38), .ZN(n495) );
  NAND2_X1 U551 ( .A1(n495), .A2(n543), .ZN(n489) );
  XNOR2_X1 U552 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U553 ( .A(G29GAT), .B(n491), .ZN(G1328GAT) );
  NAND2_X1 U554 ( .A1(n495), .A2(n514), .ZN(n492) );
  XNOR2_X1 U555 ( .A(n492), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U556 ( .A1(n495), .A2(n525), .ZN(n493) );
  XNOR2_X1 U557 ( .A(n493), .B(KEYINPUT40), .ZN(n494) );
  XNOR2_X1 U558 ( .A(G43GAT), .B(n494), .ZN(G1330GAT) );
  NAND2_X1 U559 ( .A1(n495), .A2(n518), .ZN(n496) );
  XNOR2_X1 U560 ( .A(n496), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U561 ( .A(KEYINPUT42), .B(KEYINPUT104), .Z(n499) );
  NAND2_X1 U562 ( .A1(n568), .A2(n529), .ZN(n509) );
  NOR2_X1 U563 ( .A1(n497), .A2(n509), .ZN(n505) );
  NAND2_X1 U564 ( .A1(n505), .A2(n543), .ZN(n498) );
  XNOR2_X1 U565 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U566 ( .A(G57GAT), .B(n500), .Z(G1332GAT) );
  NAND2_X1 U567 ( .A1(n505), .A2(n514), .ZN(n501) );
  XNOR2_X1 U568 ( .A(n501), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U569 ( .A1(n525), .A2(n505), .ZN(n502) );
  XNOR2_X1 U570 ( .A(n502), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT107), .B(KEYINPUT106), .Z(n504) );
  XNOR2_X1 U572 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n503) );
  XNOR2_X1 U573 ( .A(n504), .B(n503), .ZN(n508) );
  NAND2_X1 U574 ( .A1(n505), .A2(n518), .ZN(n506) );
  XNOR2_X1 U575 ( .A(n506), .B(KEYINPUT105), .ZN(n507) );
  XNOR2_X1 U576 ( .A(n508), .B(n507), .ZN(G1335GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n512) );
  NOR2_X1 U578 ( .A1(n510), .A2(n509), .ZN(n519) );
  NAND2_X1 U579 ( .A1(n519), .A2(n543), .ZN(n511) );
  XNOR2_X1 U580 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U581 ( .A(G85GAT), .B(n513), .ZN(G1336GAT) );
  NAND2_X1 U582 ( .A1(n519), .A2(n514), .ZN(n515) );
  XNOR2_X1 U583 ( .A(n515), .B(KEYINPUT110), .ZN(n516) );
  XNOR2_X1 U584 ( .A(G92GAT), .B(n516), .ZN(G1337GAT) );
  NAND2_X1 U585 ( .A1(n525), .A2(n519), .ZN(n517) );
  XNOR2_X1 U586 ( .A(n517), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U587 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n520), .B(KEYINPUT44), .ZN(n521) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n521), .ZN(G1339GAT) );
  NAND2_X1 U590 ( .A1(n522), .A2(n523), .ZN(n545) );
  NOR2_X1 U591 ( .A1(n545), .A2(n524), .ZN(n526) );
  NAND2_X1 U592 ( .A1(n526), .A2(n525), .ZN(n538) );
  NOR2_X1 U593 ( .A1(n568), .A2(n538), .ZN(n528) );
  XNOR2_X1 U594 ( .A(G113GAT), .B(KEYINPUT115), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n528), .B(n527), .ZN(G1340GAT) );
  XOR2_X1 U596 ( .A(G120GAT), .B(KEYINPUT117), .Z(n531) );
  INV_X1 U597 ( .A(n538), .ZN(n534) );
  NAND2_X1 U598 ( .A1(n534), .A2(n529), .ZN(n530) );
  XNOR2_X1 U599 ( .A(n531), .B(n530), .ZN(n533) );
  XOR2_X1 U600 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n532) );
  XNOR2_X1 U601 ( .A(n533), .B(n532), .ZN(G1341GAT) );
  NAND2_X1 U602 ( .A1(n558), .A2(n534), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n535), .B(KEYINPUT50), .ZN(n536) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(n536), .ZN(G1342GAT) );
  NOR2_X1 U605 ( .A1(n538), .A2(n537), .ZN(n542) );
  XOR2_X1 U606 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n540) );
  XNOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT119), .ZN(n539) );
  XNOR2_X1 U608 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n542), .B(n541), .ZN(G1343GAT) );
  NAND2_X1 U610 ( .A1(n543), .A2(n566), .ZN(n544) );
  NOR2_X1 U611 ( .A1(n545), .A2(n544), .ZN(n554) );
  NAND2_X1 U612 ( .A1(n556), .A2(n554), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n546), .B(KEYINPUT120), .ZN(n547) );
  XNOR2_X1 U614 ( .A(G141GAT), .B(n547), .ZN(G1344GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n550) );
  NAND2_X1 U616 ( .A1(n554), .A2(n548), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(n551), .ZN(G1345GAT) );
  XOR2_X1 U619 ( .A(G155GAT), .B(KEYINPUT121), .Z(n553) );
  NAND2_X1 U620 ( .A1(n554), .A2(n558), .ZN(n552) );
  XNOR2_X1 U621 ( .A(n553), .B(n552), .ZN(G1346GAT) );
  NAND2_X1 U622 ( .A1(n560), .A2(n554), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n555), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U624 ( .A1(n556), .A2(n561), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n557), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U626 ( .A1(n558), .A2(n561), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n559), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U628 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n563) );
  NAND2_X1 U629 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(G1351GAT) );
  AND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n567) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n579) );
  NOR2_X1 U633 ( .A1(n568), .A2(n579), .ZN(n573) );
  XOR2_X1 U634 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n570) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(KEYINPUT60), .B(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  NOR2_X1 U639 ( .A1(n574), .A2(n579), .ZN(n576) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1353GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n579), .ZN(n578) );
  XOR2_X1 U643 ( .A(G211GAT), .B(n578), .Z(G1354GAT) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n582) );
  XNOR2_X1 U645 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

