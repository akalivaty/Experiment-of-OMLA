

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U557 ( .A1(n939), .A2(n614), .ZN(n629) );
  NOR2_X1 U558 ( .A1(G2105), .A2(G2104), .ZN(n526) );
  NOR2_X2 U559 ( .A1(G2104), .A2(n529), .ZN(n873) );
  XNOR2_X2 U560 ( .A(n610), .B(KEYINPUT64), .ZN(n623) );
  AND2_X1 U561 ( .A1(n525), .A2(n935), .ZN(n675) );
  NOR2_X1 U562 ( .A1(n533), .A2(n532), .ZN(n535) );
  AND2_X1 U563 ( .A1(n741), .A2(n740), .ZN(n757) );
  XOR2_X1 U564 ( .A(KEYINPUT64), .B(n610), .Z(n666) );
  XNOR2_X1 U565 ( .A(n674), .B(n673), .ZN(n693) );
  XNOR2_X1 U566 ( .A(KEYINPUT96), .B(KEYINPUT32), .ZN(n673) );
  NOR2_X1 U567 ( .A1(n757), .A2(n756), .ZN(n759) );
  OR2_X1 U568 ( .A1(n659), .A2(n649), .ZN(n524) );
  AND2_X1 U569 ( .A1(n663), .A2(n684), .ZN(n525) );
  INV_X1 U570 ( .A(G8), .ZN(n649) );
  OR2_X1 U571 ( .A1(n658), .A2(n524), .ZN(n650) );
  NOR2_X1 U572 ( .A1(G1966), .A2(n699), .ZN(n658) );
  NOR2_X1 U573 ( .A1(n658), .A2(n664), .ZN(n661) );
  NOR2_X1 U574 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U575 ( .A1(G651), .A2(G543), .ZN(n785) );
  AND2_X2 U576 ( .A1(G2105), .A2(G2104), .ZN(n874) );
  NOR2_X1 U577 ( .A1(G651), .A2(n577), .ZN(n789) );
  INV_X1 U578 ( .A(KEYINPUT40), .ZN(n758) );
  XOR2_X1 U579 ( .A(KEYINPUT17), .B(n526), .Z(n536) );
  AND2_X1 U580 ( .A1(n536), .A2(G138), .ZN(n533) );
  INV_X2 U581 ( .A(G2105), .ZN(n529) );
  AND2_X4 U582 ( .A1(n529), .A2(G2104), .ZN(n878) );
  NAND2_X1 U583 ( .A1(G102), .A2(n878), .ZN(n528) );
  NAND2_X1 U584 ( .A1(G114), .A2(n874), .ZN(n527) );
  AND2_X1 U585 ( .A1(n528), .A2(n527), .ZN(n531) );
  NAND2_X1 U586 ( .A1(G126), .A2(n873), .ZN(n530) );
  NAND2_X1 U587 ( .A1(n531), .A2(n530), .ZN(n532) );
  INV_X1 U588 ( .A(KEYINPUT85), .ZN(n534) );
  XNOR2_X2 U589 ( .A(n535), .B(n534), .ZN(G164) );
  BUF_X1 U590 ( .A(n536), .Z(n877) );
  NAND2_X1 U591 ( .A1(n877), .A2(G137), .ZN(n539) );
  NAND2_X1 U592 ( .A1(G101), .A2(n878), .ZN(n537) );
  XOR2_X1 U593 ( .A(KEYINPUT23), .B(n537), .Z(n538) );
  NAND2_X1 U594 ( .A1(n539), .A2(n538), .ZN(n543) );
  NAND2_X1 U595 ( .A1(G125), .A2(n873), .ZN(n541) );
  NAND2_X1 U596 ( .A1(G113), .A2(n874), .ZN(n540) );
  NAND2_X1 U597 ( .A1(n541), .A2(n540), .ZN(n542) );
  NOR2_X1 U598 ( .A1(n543), .A2(n542), .ZN(G160) );
  INV_X1 U599 ( .A(G651), .ZN(n548) );
  NOR2_X1 U600 ( .A1(G543), .A2(n548), .ZN(n544) );
  XOR2_X1 U601 ( .A(KEYINPUT1), .B(n544), .Z(n784) );
  NAND2_X1 U602 ( .A1(G65), .A2(n784), .ZN(n546) );
  XOR2_X1 U603 ( .A(KEYINPUT0), .B(G543), .Z(n577) );
  NAND2_X1 U604 ( .A1(G53), .A2(n789), .ZN(n545) );
  NAND2_X1 U605 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U606 ( .A(KEYINPUT70), .B(n547), .Z(n552) );
  NAND2_X1 U607 ( .A1(G91), .A2(n785), .ZN(n550) );
  NOR2_X1 U608 ( .A1(n577), .A2(n548), .ZN(n788) );
  NAND2_X1 U609 ( .A1(G78), .A2(n788), .ZN(n549) );
  AND2_X1 U610 ( .A1(n550), .A2(n549), .ZN(n551) );
  NAND2_X1 U611 ( .A1(n552), .A2(n551), .ZN(G299) );
  XNOR2_X1 U612 ( .A(KEYINPUT67), .B(KEYINPUT68), .ZN(n557) );
  NAND2_X1 U613 ( .A1(G90), .A2(n785), .ZN(n554) );
  NAND2_X1 U614 ( .A1(G77), .A2(n788), .ZN(n553) );
  NAND2_X1 U615 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U616 ( .A(n555), .B(KEYINPUT9), .ZN(n556) );
  XNOR2_X1 U617 ( .A(n557), .B(n556), .ZN(n562) );
  NAND2_X1 U618 ( .A1(n784), .A2(G64), .ZN(n558) );
  XNOR2_X1 U619 ( .A(n558), .B(KEYINPUT66), .ZN(n560) );
  NAND2_X1 U620 ( .A1(G52), .A2(n789), .ZN(n559) );
  NAND2_X1 U621 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U622 ( .A1(n562), .A2(n561), .ZN(G171) );
  NAND2_X1 U623 ( .A1(n785), .A2(G89), .ZN(n563) );
  XNOR2_X1 U624 ( .A(n563), .B(KEYINPUT4), .ZN(n565) );
  NAND2_X1 U625 ( .A1(G76), .A2(n788), .ZN(n564) );
  NAND2_X1 U626 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U627 ( .A(KEYINPUT5), .B(n566), .ZN(n572) );
  NAND2_X1 U628 ( .A1(G63), .A2(n784), .ZN(n568) );
  NAND2_X1 U629 ( .A1(G51), .A2(n789), .ZN(n567) );
  NAND2_X1 U630 ( .A1(n568), .A2(n567), .ZN(n570) );
  XOR2_X1 U631 ( .A(KEYINPUT6), .B(KEYINPUT72), .Z(n569) );
  XNOR2_X1 U632 ( .A(n570), .B(n569), .ZN(n571) );
  NAND2_X1 U633 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U634 ( .A(KEYINPUT7), .B(n573), .ZN(G168) );
  NAND2_X1 U635 ( .A1(G49), .A2(n789), .ZN(n575) );
  NAND2_X1 U636 ( .A1(G74), .A2(G651), .ZN(n574) );
  NAND2_X1 U637 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U638 ( .A1(n784), .A2(n576), .ZN(n579) );
  NAND2_X1 U639 ( .A1(n577), .A2(G87), .ZN(n578) );
  NAND2_X1 U640 ( .A1(n579), .A2(n578), .ZN(G288) );
  XOR2_X1 U641 ( .A(KEYINPUT78), .B(KEYINPUT2), .Z(n581) );
  NAND2_X1 U642 ( .A1(G73), .A2(n788), .ZN(n580) );
  XNOR2_X1 U643 ( .A(n581), .B(n580), .ZN(n585) );
  NAND2_X1 U644 ( .A1(G61), .A2(n784), .ZN(n583) );
  NAND2_X1 U645 ( .A1(G86), .A2(n785), .ZN(n582) );
  NAND2_X1 U646 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U647 ( .A1(n585), .A2(n584), .ZN(n587) );
  NAND2_X1 U648 ( .A1(n789), .A2(G48), .ZN(n586) );
  NAND2_X1 U649 ( .A1(n587), .A2(n586), .ZN(G305) );
  XOR2_X1 U650 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U651 ( .A1(G88), .A2(n785), .ZN(n589) );
  NAND2_X1 U652 ( .A1(G75), .A2(n788), .ZN(n588) );
  NAND2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n593) );
  NAND2_X1 U654 ( .A1(G62), .A2(n784), .ZN(n591) );
  NAND2_X1 U655 ( .A1(G50), .A2(n789), .ZN(n590) );
  NAND2_X1 U656 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U657 ( .A1(n593), .A2(n592), .ZN(G166) );
  INV_X1 U658 ( .A(G166), .ZN(G303) );
  NAND2_X1 U659 ( .A1(G85), .A2(n785), .ZN(n595) );
  NAND2_X1 U660 ( .A1(G72), .A2(n788), .ZN(n594) );
  NAND2_X1 U661 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U662 ( .A1(G60), .A2(n784), .ZN(n597) );
  NAND2_X1 U663 ( .A1(G47), .A2(n789), .ZN(n596) );
  NAND2_X1 U664 ( .A1(n597), .A2(n596), .ZN(n598) );
  OR2_X1 U665 ( .A1(n599), .A2(n598), .ZN(G290) );
  NOR2_X1 U666 ( .A1(G164), .A2(G1384), .ZN(n600) );
  XNOR2_X1 U667 ( .A(n600), .B(KEYINPUT65), .ZN(n705) );
  NAND2_X1 U668 ( .A1(G160), .A2(G40), .ZN(n706) );
  NOR2_X2 U669 ( .A1(n705), .A2(n706), .ZN(n610) );
  NAND2_X1 U670 ( .A1(n666), .A2(G8), .ZN(n699) );
  NAND2_X1 U671 ( .A1(G56), .A2(n784), .ZN(n601) );
  XOR2_X1 U672 ( .A(KEYINPUT14), .B(n601), .Z(n607) );
  NAND2_X1 U673 ( .A1(n785), .A2(G81), .ZN(n602) );
  XNOR2_X1 U674 ( .A(n602), .B(KEYINPUT12), .ZN(n604) );
  NAND2_X1 U675 ( .A1(G68), .A2(n788), .ZN(n603) );
  NAND2_X1 U676 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X1 U677 ( .A(KEYINPUT13), .B(n605), .Z(n606) );
  NOR2_X1 U678 ( .A1(n607), .A2(n606), .ZN(n609) );
  NAND2_X1 U679 ( .A1(n789), .A2(G43), .ZN(n608) );
  NAND2_X1 U680 ( .A1(n609), .A2(n608), .ZN(n939) );
  NAND2_X1 U681 ( .A1(n623), .A2(G1996), .ZN(n611) );
  XNOR2_X1 U682 ( .A(n611), .B(KEYINPUT26), .ZN(n613) );
  NAND2_X1 U683 ( .A1(n666), .A2(G1341), .ZN(n612) );
  NAND2_X1 U684 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U685 ( .A1(G66), .A2(n784), .ZN(n616) );
  NAND2_X1 U686 ( .A1(G92), .A2(n785), .ZN(n615) );
  NAND2_X1 U687 ( .A1(n616), .A2(n615), .ZN(n621) );
  NAND2_X1 U688 ( .A1(G79), .A2(n788), .ZN(n618) );
  NAND2_X1 U689 ( .A1(G54), .A2(n789), .ZN(n617) );
  NAND2_X1 U690 ( .A1(n618), .A2(n617), .ZN(n619) );
  XOR2_X1 U691 ( .A(KEYINPUT71), .B(n619), .Z(n620) );
  NOR2_X1 U692 ( .A1(n621), .A2(n620), .ZN(n622) );
  XOR2_X1 U693 ( .A(KEYINPUT15), .B(n622), .Z(n897) );
  NAND2_X1 U694 ( .A1(n629), .A2(n897), .ZN(n627) );
  NOR2_X1 U695 ( .A1(G1348), .A2(n623), .ZN(n625) );
  NOR2_X1 U696 ( .A1(G2067), .A2(n666), .ZN(n624) );
  NOR2_X1 U697 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U698 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U699 ( .A(n628), .B(KEYINPUT94), .ZN(n631) );
  OR2_X1 U700 ( .A1(n629), .A2(n897), .ZN(n630) );
  NAND2_X1 U701 ( .A1(n631), .A2(n630), .ZN(n636) );
  INV_X1 U702 ( .A(G299), .ZN(n924) );
  NAND2_X1 U703 ( .A1(G2072), .A2(n623), .ZN(n632) );
  XNOR2_X1 U704 ( .A(n632), .B(KEYINPUT27), .ZN(n634) );
  INV_X1 U705 ( .A(G1956), .ZN(n951) );
  NOR2_X1 U706 ( .A1(n623), .A2(n951), .ZN(n633) );
  NOR2_X1 U707 ( .A1(n634), .A2(n633), .ZN(n637) );
  NAND2_X1 U708 ( .A1(n924), .A2(n637), .ZN(n635) );
  NAND2_X1 U709 ( .A1(n636), .A2(n635), .ZN(n641) );
  NOR2_X1 U710 ( .A1(n924), .A2(n637), .ZN(n639) );
  XNOR2_X1 U711 ( .A(KEYINPUT93), .B(KEYINPUT28), .ZN(n638) );
  XNOR2_X1 U712 ( .A(n639), .B(n638), .ZN(n640) );
  NAND2_X1 U713 ( .A1(n641), .A2(n640), .ZN(n643) );
  XOR2_X1 U714 ( .A(KEYINPUT95), .B(KEYINPUT29), .Z(n642) );
  XNOR2_X1 U715 ( .A(n643), .B(n642), .ZN(n648) );
  XOR2_X1 U716 ( .A(G2078), .B(KEYINPUT25), .Z(n1011) );
  NAND2_X1 U717 ( .A1(n623), .A2(n1011), .ZN(n645) );
  NAND2_X1 U718 ( .A1(n666), .A2(G1961), .ZN(n644) );
  NAND2_X1 U719 ( .A1(n645), .A2(n644), .ZN(n646) );
  XOR2_X1 U720 ( .A(n646), .B(KEYINPUT92), .Z(n652) );
  AND2_X1 U721 ( .A1(n652), .A2(G171), .ZN(n647) );
  NOR2_X1 U722 ( .A1(n648), .A2(n647), .ZN(n657) );
  NOR2_X1 U723 ( .A1(n666), .A2(G2084), .ZN(n659) );
  XNOR2_X1 U724 ( .A(KEYINPUT30), .B(n650), .ZN(n651) );
  NOR2_X1 U725 ( .A1(G168), .A2(n651), .ZN(n654) );
  NOR2_X1 U726 ( .A1(G171), .A2(n652), .ZN(n653) );
  NOR2_X1 U727 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U728 ( .A(n655), .B(KEYINPUT31), .ZN(n656) );
  NOR2_X1 U729 ( .A1(n657), .A2(n656), .ZN(n664) );
  NAND2_X1 U730 ( .A1(n659), .A2(G8), .ZN(n660) );
  NAND2_X1 U731 ( .A1(n661), .A2(n660), .ZN(n694) );
  NAND2_X1 U732 ( .A1(G1976), .A2(G288), .ZN(n922) );
  AND2_X1 U733 ( .A1(n694), .A2(n922), .ZN(n663) );
  NOR2_X1 U734 ( .A1(G1976), .A2(G288), .ZN(n920) );
  NAND2_X1 U735 ( .A1(n920), .A2(KEYINPUT33), .ZN(n662) );
  OR2_X1 U736 ( .A1(n662), .A2(n699), .ZN(n684) );
  XOR2_X1 U737 ( .A(G1981), .B(G305), .Z(n935) );
  INV_X1 U738 ( .A(n664), .ZN(n665) );
  NAND2_X1 U739 ( .A1(n665), .A2(G286), .ZN(n672) );
  NOR2_X1 U740 ( .A1(n666), .A2(G2090), .ZN(n668) );
  NOR2_X1 U741 ( .A1(G1971), .A2(n699), .ZN(n667) );
  NOR2_X1 U742 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U743 ( .A1(n669), .A2(G303), .ZN(n670) );
  OR2_X1 U744 ( .A1(n649), .A2(n670), .ZN(n671) );
  AND2_X1 U745 ( .A1(n672), .A2(n671), .ZN(n674) );
  NAND2_X1 U746 ( .A1(n675), .A2(n693), .ZN(n688) );
  INV_X1 U747 ( .A(n935), .ZN(n686) );
  INV_X1 U748 ( .A(n922), .ZN(n679) );
  NOR2_X1 U749 ( .A1(G1971), .A2(G303), .ZN(n676) );
  NOR2_X1 U750 ( .A1(n920), .A2(n676), .ZN(n677) );
  XOR2_X1 U751 ( .A(KEYINPUT97), .B(n677), .Z(n678) );
  OR2_X1 U752 ( .A1(n679), .A2(n678), .ZN(n680) );
  OR2_X1 U753 ( .A1(n699), .A2(n680), .ZN(n682) );
  INV_X1 U754 ( .A(KEYINPUT33), .ZN(n681) );
  NAND2_X1 U755 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U756 ( .A1(n684), .A2(n683), .ZN(n685) );
  OR2_X1 U757 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U758 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U759 ( .A(n689), .B(KEYINPUT98), .ZN(n703) );
  NOR2_X1 U760 ( .A1(G1981), .A2(G305), .ZN(n690) );
  XNOR2_X1 U761 ( .A(KEYINPUT24), .B(n690), .ZN(n692) );
  INV_X1 U762 ( .A(n699), .ZN(n691) );
  NAND2_X1 U763 ( .A1(n692), .A2(n691), .ZN(n701) );
  NAND2_X1 U764 ( .A1(n694), .A2(n693), .ZN(n697) );
  NOR2_X1 U765 ( .A1(G2090), .A2(G303), .ZN(n695) );
  NAND2_X1 U766 ( .A1(G8), .A2(n695), .ZN(n696) );
  NAND2_X1 U767 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U768 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U769 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U770 ( .A(n704), .B(KEYINPUT99), .ZN(n741) );
  INV_X1 U771 ( .A(n705), .ZN(n707) );
  NOR2_X1 U772 ( .A1(n707), .A2(n706), .ZN(n754) );
  XNOR2_X1 U773 ( .A(G1986), .B(G290), .ZN(n931) );
  AND2_X1 U774 ( .A1(n754), .A2(n931), .ZN(n739) );
  NAND2_X1 U775 ( .A1(n878), .A2(G105), .ZN(n709) );
  XNOR2_X1 U776 ( .A(KEYINPUT88), .B(KEYINPUT38), .ZN(n708) );
  XNOR2_X1 U777 ( .A(n709), .B(n708), .ZN(n716) );
  NAND2_X1 U778 ( .A1(G129), .A2(n873), .ZN(n711) );
  NAND2_X1 U779 ( .A1(G117), .A2(n874), .ZN(n710) );
  NAND2_X1 U780 ( .A1(n711), .A2(n710), .ZN(n714) );
  NAND2_X1 U781 ( .A1(G141), .A2(n877), .ZN(n712) );
  XNOR2_X1 U782 ( .A(KEYINPUT89), .B(n712), .ZN(n713) );
  NOR2_X1 U783 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U784 ( .A1(n716), .A2(n715), .ZN(n872) );
  NAND2_X1 U785 ( .A1(n872), .A2(G1996), .ZN(n725) );
  NAND2_X1 U786 ( .A1(G119), .A2(n873), .ZN(n718) );
  NAND2_X1 U787 ( .A1(G131), .A2(n877), .ZN(n717) );
  NAND2_X1 U788 ( .A1(n718), .A2(n717), .ZN(n722) );
  NAND2_X1 U789 ( .A1(G107), .A2(n874), .ZN(n720) );
  NAND2_X1 U790 ( .A1(G95), .A2(n878), .ZN(n719) );
  NAND2_X1 U791 ( .A1(n720), .A2(n719), .ZN(n721) );
  OR2_X1 U792 ( .A1(n722), .A2(n721), .ZN(n860) );
  NAND2_X1 U793 ( .A1(G1991), .A2(n860), .ZN(n723) );
  XOR2_X1 U794 ( .A(KEYINPUT87), .B(n723), .Z(n724) );
  NAND2_X1 U795 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U796 ( .A(n726), .B(KEYINPUT90), .ZN(n998) );
  NAND2_X1 U797 ( .A1(n754), .A2(n998), .ZN(n742) );
  NAND2_X1 U798 ( .A1(n877), .A2(G140), .ZN(n727) );
  XNOR2_X1 U799 ( .A(n727), .B(KEYINPUT86), .ZN(n729) );
  NAND2_X1 U800 ( .A1(G104), .A2(n878), .ZN(n728) );
  NAND2_X1 U801 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U802 ( .A(KEYINPUT34), .B(n730), .ZN(n735) );
  NAND2_X1 U803 ( .A1(G128), .A2(n873), .ZN(n732) );
  NAND2_X1 U804 ( .A1(G116), .A2(n874), .ZN(n731) );
  NAND2_X1 U805 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U806 ( .A(KEYINPUT35), .B(n733), .Z(n734) );
  NOR2_X1 U807 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U808 ( .A(KEYINPUT36), .B(n736), .ZN(n890) );
  XNOR2_X1 U809 ( .A(KEYINPUT37), .B(G2067), .ZN(n751) );
  NOR2_X1 U810 ( .A1(n890), .A2(n751), .ZN(n1002) );
  NAND2_X1 U811 ( .A1(n754), .A2(n1002), .ZN(n749) );
  NAND2_X1 U812 ( .A1(n742), .A2(n749), .ZN(n737) );
  XOR2_X1 U813 ( .A(KEYINPUT91), .B(n737), .Z(n738) );
  NOR2_X1 U814 ( .A1(n739), .A2(n738), .ZN(n740) );
  INV_X1 U815 ( .A(n742), .ZN(n745) );
  NOR2_X1 U816 ( .A1(G1986), .A2(G290), .ZN(n743) );
  NOR2_X1 U817 ( .A1(G1991), .A2(n860), .ZN(n988) );
  NOR2_X1 U818 ( .A1(n743), .A2(n988), .ZN(n744) );
  NOR2_X1 U819 ( .A1(n745), .A2(n744), .ZN(n747) );
  NOR2_X1 U820 ( .A1(n872), .A2(G1996), .ZN(n746) );
  XNOR2_X1 U821 ( .A(n746), .B(KEYINPUT100), .ZN(n983) );
  NOR2_X1 U822 ( .A1(n747), .A2(n983), .ZN(n748) );
  XNOR2_X1 U823 ( .A(n748), .B(KEYINPUT39), .ZN(n750) );
  NAND2_X1 U824 ( .A1(n750), .A2(n749), .ZN(n752) );
  NAND2_X1 U825 ( .A1(n890), .A2(n751), .ZN(n1003) );
  NAND2_X1 U826 ( .A1(n752), .A2(n1003), .ZN(n753) );
  NAND2_X1 U827 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U828 ( .A(KEYINPUT101), .B(n755), .ZN(n756) );
  XNOR2_X1 U829 ( .A(n759), .B(n758), .ZN(G329) );
  INV_X1 U830 ( .A(G108), .ZN(G238) );
  INV_X1 U831 ( .A(G120), .ZN(G236) );
  INV_X1 U832 ( .A(G69), .ZN(G235) );
  INV_X1 U833 ( .A(G132), .ZN(G219) );
  INV_X1 U834 ( .A(G82), .ZN(G220) );
  NAND2_X1 U835 ( .A1(G94), .A2(G452), .ZN(n760) );
  XNOR2_X1 U836 ( .A(n760), .B(KEYINPUT69), .ZN(G173) );
  NAND2_X1 U837 ( .A1(G7), .A2(G661), .ZN(n761) );
  XNOR2_X1 U838 ( .A(n761), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U839 ( .A(G223), .ZN(n827) );
  NAND2_X1 U840 ( .A1(n827), .A2(G567), .ZN(n762) );
  XOR2_X1 U841 ( .A(KEYINPUT11), .B(n762), .Z(G234) );
  INV_X1 U842 ( .A(G860), .ZN(n768) );
  OR2_X1 U843 ( .A1(n939), .A2(n768), .ZN(G153) );
  INV_X1 U844 ( .A(G171), .ZN(G301) );
  NAND2_X1 U845 ( .A1(G868), .A2(G301), .ZN(n764) );
  INV_X1 U846 ( .A(n897), .ZN(n944) );
  INV_X1 U847 ( .A(G868), .ZN(n806) );
  NAND2_X1 U848 ( .A1(n944), .A2(n806), .ZN(n763) );
  NAND2_X1 U849 ( .A1(n764), .A2(n763), .ZN(G284) );
  XNOR2_X1 U850 ( .A(KEYINPUT73), .B(G868), .ZN(n765) );
  NOR2_X1 U851 ( .A1(G286), .A2(n765), .ZN(n767) );
  NOR2_X1 U852 ( .A1(G868), .A2(G299), .ZN(n766) );
  NOR2_X1 U853 ( .A1(n767), .A2(n766), .ZN(G297) );
  NAND2_X1 U854 ( .A1(n768), .A2(G559), .ZN(n769) );
  NAND2_X1 U855 ( .A1(n769), .A2(n897), .ZN(n770) );
  XNOR2_X1 U856 ( .A(n770), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U857 ( .A1(G868), .A2(n939), .ZN(n773) );
  NAND2_X1 U858 ( .A1(n897), .A2(G868), .ZN(n771) );
  NOR2_X1 U859 ( .A1(G559), .A2(n771), .ZN(n772) );
  NOR2_X1 U860 ( .A1(n773), .A2(n772), .ZN(G282) );
  XNOR2_X1 U861 ( .A(G2100), .B(KEYINPUT75), .ZN(n783) );
  NAND2_X1 U862 ( .A1(n873), .A2(G123), .ZN(n774) );
  XNOR2_X1 U863 ( .A(n774), .B(KEYINPUT18), .ZN(n776) );
  NAND2_X1 U864 ( .A1(G135), .A2(n877), .ZN(n775) );
  NAND2_X1 U865 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U866 ( .A(KEYINPUT74), .B(n777), .ZN(n781) );
  NAND2_X1 U867 ( .A1(G111), .A2(n874), .ZN(n779) );
  NAND2_X1 U868 ( .A1(G99), .A2(n878), .ZN(n778) );
  NAND2_X1 U869 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U870 ( .A1(n781), .A2(n780), .ZN(n994) );
  XNOR2_X1 U871 ( .A(n994), .B(G2096), .ZN(n782) );
  NAND2_X1 U872 ( .A1(n783), .A2(n782), .ZN(G156) );
  NAND2_X1 U873 ( .A1(G67), .A2(n784), .ZN(n787) );
  NAND2_X1 U874 ( .A1(G93), .A2(n785), .ZN(n786) );
  NAND2_X1 U875 ( .A1(n787), .A2(n786), .ZN(n793) );
  NAND2_X1 U876 ( .A1(G80), .A2(n788), .ZN(n791) );
  NAND2_X1 U877 ( .A1(G55), .A2(n789), .ZN(n790) );
  NAND2_X1 U878 ( .A1(n791), .A2(n790), .ZN(n792) );
  OR2_X1 U879 ( .A1(n793), .A2(n792), .ZN(n807) );
  XNOR2_X1 U880 ( .A(n939), .B(KEYINPUT76), .ZN(n795) );
  NAND2_X1 U881 ( .A1(n897), .A2(G559), .ZN(n794) );
  XNOR2_X1 U882 ( .A(n795), .B(n794), .ZN(n804) );
  XOR2_X1 U883 ( .A(n804), .B(KEYINPUT77), .Z(n796) );
  NOR2_X1 U884 ( .A1(G860), .A2(n796), .ZN(n797) );
  XOR2_X1 U885 ( .A(n807), .B(n797), .Z(G145) );
  XOR2_X1 U886 ( .A(KEYINPUT19), .B(KEYINPUT79), .Z(n799) );
  XNOR2_X1 U887 ( .A(G166), .B(n924), .ZN(n798) );
  XNOR2_X1 U888 ( .A(n799), .B(n798), .ZN(n800) );
  XNOR2_X1 U889 ( .A(n807), .B(n800), .ZN(n801) );
  XNOR2_X1 U890 ( .A(G305), .B(n801), .ZN(n802) );
  XNOR2_X1 U891 ( .A(n802), .B(G290), .ZN(n803) );
  XNOR2_X1 U892 ( .A(n803), .B(G288), .ZN(n893) );
  XOR2_X1 U893 ( .A(n893), .B(n804), .Z(n805) );
  NOR2_X1 U894 ( .A1(n806), .A2(n805), .ZN(n809) );
  NOR2_X1 U895 ( .A1(G868), .A2(n807), .ZN(n808) );
  NOR2_X1 U896 ( .A1(n809), .A2(n808), .ZN(G295) );
  NAND2_X1 U897 ( .A1(G2078), .A2(G2084), .ZN(n810) );
  XOR2_X1 U898 ( .A(KEYINPUT20), .B(n810), .Z(n811) );
  NAND2_X1 U899 ( .A1(n811), .A2(G2090), .ZN(n812) );
  XNOR2_X1 U900 ( .A(n812), .B(KEYINPUT80), .ZN(n813) );
  XNOR2_X1 U901 ( .A(KEYINPUT21), .B(n813), .ZN(n814) );
  NAND2_X1 U902 ( .A1(G2072), .A2(n814), .ZN(G158) );
  XNOR2_X1 U903 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U904 ( .A1(G220), .A2(G219), .ZN(n815) );
  XOR2_X1 U905 ( .A(KEYINPUT22), .B(n815), .Z(n816) );
  NOR2_X1 U906 ( .A1(G218), .A2(n816), .ZN(n817) );
  XOR2_X1 U907 ( .A(KEYINPUT81), .B(n817), .Z(n818) );
  NAND2_X1 U908 ( .A1(G96), .A2(n818), .ZN(n832) );
  NAND2_X1 U909 ( .A1(n832), .A2(G2106), .ZN(n824) );
  NOR2_X1 U910 ( .A1(G235), .A2(G236), .ZN(n819) );
  XNOR2_X1 U911 ( .A(KEYINPUT82), .B(n819), .ZN(n820) );
  NAND2_X1 U912 ( .A1(n820), .A2(G57), .ZN(n821) );
  NOR2_X1 U913 ( .A1(n821), .A2(G238), .ZN(n822) );
  XNOR2_X1 U914 ( .A(n822), .B(KEYINPUT83), .ZN(n833) );
  NAND2_X1 U915 ( .A1(n833), .A2(G567), .ZN(n823) );
  NAND2_X1 U916 ( .A1(n824), .A2(n823), .ZN(n834) );
  NAND2_X1 U917 ( .A1(G483), .A2(G661), .ZN(n825) );
  NOR2_X1 U918 ( .A1(n834), .A2(n825), .ZN(n829) );
  NAND2_X1 U919 ( .A1(n829), .A2(G36), .ZN(n826) );
  XNOR2_X1 U920 ( .A(KEYINPUT84), .B(n826), .ZN(G176) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n827), .ZN(G217) );
  AND2_X1 U922 ( .A1(G15), .A2(G2), .ZN(n828) );
  NAND2_X1 U923 ( .A1(G661), .A2(n828), .ZN(G259) );
  NAND2_X1 U924 ( .A1(G3), .A2(G1), .ZN(n830) );
  NAND2_X1 U925 ( .A1(n830), .A2(n829), .ZN(n831) );
  XNOR2_X1 U926 ( .A(n831), .B(KEYINPUT104), .ZN(G188) );
  INV_X1 U928 ( .A(G96), .ZN(G221) );
  INV_X1 U929 ( .A(G57), .ZN(G237) );
  NOR2_X1 U930 ( .A1(n833), .A2(n832), .ZN(G325) );
  INV_X1 U931 ( .A(G325), .ZN(G261) );
  INV_X1 U932 ( .A(n834), .ZN(G319) );
  XOR2_X1 U933 ( .A(KEYINPUT105), .B(G2084), .Z(n836) );
  XNOR2_X1 U934 ( .A(G2072), .B(G2078), .ZN(n835) );
  XNOR2_X1 U935 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U936 ( .A(n837), .B(G2096), .Z(n839) );
  XNOR2_X1 U937 ( .A(G2067), .B(G2090), .ZN(n838) );
  XNOR2_X1 U938 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U939 ( .A(G2100), .B(KEYINPUT43), .Z(n841) );
  XNOR2_X1 U940 ( .A(G2678), .B(KEYINPUT42), .ZN(n840) );
  XNOR2_X1 U941 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U942 ( .A(n843), .B(n842), .Z(G227) );
  XOR2_X1 U943 ( .A(G1981), .B(G1966), .Z(n845) );
  XNOR2_X1 U944 ( .A(G1986), .B(G1956), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U946 ( .A(n846), .B(KEYINPUT41), .Z(n848) );
  XNOR2_X1 U947 ( .A(G1971), .B(G1976), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U949 ( .A(G2474), .B(G1961), .Z(n850) );
  XNOR2_X1 U950 ( .A(G1996), .B(G1991), .ZN(n849) );
  XNOR2_X1 U951 ( .A(n850), .B(n849), .ZN(n851) );
  XNOR2_X1 U952 ( .A(n852), .B(n851), .ZN(G229) );
  NAND2_X1 U953 ( .A1(n873), .A2(G124), .ZN(n853) );
  XNOR2_X1 U954 ( .A(n853), .B(KEYINPUT44), .ZN(n855) );
  NAND2_X1 U955 ( .A1(G112), .A2(n874), .ZN(n854) );
  NAND2_X1 U956 ( .A1(n855), .A2(n854), .ZN(n859) );
  NAND2_X1 U957 ( .A1(G136), .A2(n877), .ZN(n857) );
  NAND2_X1 U958 ( .A1(G100), .A2(n878), .ZN(n856) );
  NAND2_X1 U959 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U960 ( .A1(n859), .A2(n858), .ZN(G162) );
  XNOR2_X1 U961 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n860), .B(KEYINPUT106), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n862), .B(n861), .ZN(n863) );
  XNOR2_X1 U964 ( .A(G164), .B(n863), .ZN(n889) );
  NAND2_X1 U965 ( .A1(G139), .A2(n877), .ZN(n865) );
  NAND2_X1 U966 ( .A1(G103), .A2(n878), .ZN(n864) );
  NAND2_X1 U967 ( .A1(n865), .A2(n864), .ZN(n870) );
  NAND2_X1 U968 ( .A1(G127), .A2(n873), .ZN(n867) );
  NAND2_X1 U969 ( .A1(G115), .A2(n874), .ZN(n866) );
  NAND2_X1 U970 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U971 ( .A(KEYINPUT47), .B(n868), .Z(n869) );
  NOR2_X1 U972 ( .A1(n870), .A2(n869), .ZN(n989) );
  XOR2_X1 U973 ( .A(n994), .B(n989), .Z(n871) );
  XNOR2_X1 U974 ( .A(n872), .B(n871), .ZN(n885) );
  NAND2_X1 U975 ( .A1(G130), .A2(n873), .ZN(n876) );
  NAND2_X1 U976 ( .A1(G118), .A2(n874), .ZN(n875) );
  NAND2_X1 U977 ( .A1(n876), .A2(n875), .ZN(n883) );
  NAND2_X1 U978 ( .A1(G142), .A2(n877), .ZN(n880) );
  NAND2_X1 U979 ( .A1(G106), .A2(n878), .ZN(n879) );
  NAND2_X1 U980 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U981 ( .A(KEYINPUT45), .B(n881), .Z(n882) );
  NOR2_X1 U982 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U983 ( .A(n885), .B(n884), .Z(n887) );
  XNOR2_X1 U984 ( .A(G160), .B(G162), .ZN(n886) );
  XNOR2_X1 U985 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U986 ( .A(n889), .B(n888), .ZN(n891) );
  XNOR2_X1 U987 ( .A(n891), .B(n890), .ZN(n892) );
  NOR2_X1 U988 ( .A1(G37), .A2(n892), .ZN(G395) );
  XOR2_X1 U989 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n895) );
  XNOR2_X1 U990 ( .A(G171), .B(n893), .ZN(n894) );
  XNOR2_X1 U991 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U992 ( .A(n939), .B(n896), .ZN(n899) );
  XNOR2_X1 U993 ( .A(G286), .B(n897), .ZN(n898) );
  XNOR2_X1 U994 ( .A(n899), .B(n898), .ZN(n900) );
  NOR2_X1 U995 ( .A1(G37), .A2(n900), .ZN(n901) );
  XOR2_X1 U996 ( .A(KEYINPUT109), .B(n901), .Z(G397) );
  XNOR2_X1 U997 ( .A(G2443), .B(G2427), .ZN(n911) );
  XOR2_X1 U998 ( .A(G2430), .B(KEYINPUT103), .Z(n903) );
  XNOR2_X1 U999 ( .A(G2454), .B(G2435), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n907) );
  XOR2_X1 U1001 ( .A(G2438), .B(KEYINPUT102), .Z(n905) );
  XNOR2_X1 U1002 ( .A(G1341), .B(G1348), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1004 ( .A(n907), .B(n906), .Z(n909) );
  XNOR2_X1 U1005 ( .A(G2451), .B(G2446), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(n911), .B(n910), .ZN(n912) );
  NAND2_X1 U1008 ( .A1(n912), .A2(G14), .ZN(n918) );
  NAND2_X1 U1009 ( .A1(G319), .A2(n918), .ZN(n915) );
  NOR2_X1 U1010 ( .A1(G227), .A2(G229), .ZN(n913) );
  XNOR2_X1 U1011 ( .A(KEYINPUT49), .B(n913), .ZN(n914) );
  NOR2_X1 U1012 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1014 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(n918), .ZN(G401) );
  INV_X1 U1017 ( .A(G16), .ZN(n979) );
  XNOR2_X1 U1018 ( .A(KEYINPUT56), .B(KEYINPUT115), .ZN(n919) );
  XNOR2_X1 U1019 ( .A(n979), .B(n919), .ZN(n950) );
  INV_X1 U1020 ( .A(n920), .ZN(n921) );
  NAND2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n923) );
  XOR2_X1 U1022 ( .A(KEYINPUT119), .B(n923), .Z(n928) );
  XNOR2_X1 U1023 ( .A(n924), .B(G1956), .ZN(n926) );
  XNOR2_X1 U1024 ( .A(G166), .B(G1971), .ZN(n925) );
  NAND2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1027 ( .A(KEYINPUT120), .B(n929), .Z(n930) );
  NOR2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1029 ( .A(KEYINPUT121), .B(n932), .Z(n948) );
  XNOR2_X1 U1030 ( .A(G168), .B(G1966), .ZN(n933) );
  XNOR2_X1 U1031 ( .A(n933), .B(KEYINPUT116), .ZN(n934) );
  NAND2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n938) );
  XOR2_X1 U1033 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n936) );
  XNOR2_X1 U1034 ( .A(KEYINPUT57), .B(n936), .ZN(n937) );
  XNOR2_X1 U1035 ( .A(n938), .B(n937), .ZN(n943) );
  XNOR2_X1 U1036 ( .A(n939), .B(G1341), .ZN(n941) );
  XNOR2_X1 U1037 ( .A(G301), .B(G1961), .ZN(n940) );
  NOR2_X1 U1038 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1039 ( .A1(n943), .A2(n942), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(G1348), .B(n944), .ZN(n945) );
  NOR2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1043 ( .A1(n950), .A2(n949), .ZN(n981) );
  XNOR2_X1 U1044 ( .A(n951), .B(G20), .ZN(n959) );
  XOR2_X1 U1045 ( .A(G1341), .B(G19), .Z(n954) );
  XOR2_X1 U1046 ( .A(G6), .B(KEYINPUT122), .Z(n952) );
  XNOR2_X1 U1047 ( .A(G1981), .B(n952), .ZN(n953) );
  NAND2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n957) );
  XOR2_X1 U1049 ( .A(KEYINPUT59), .B(G1348), .Z(n955) );
  XNOR2_X1 U1050 ( .A(G4), .B(n955), .ZN(n956) );
  NOR2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(n960), .B(KEYINPUT60), .ZN(n975) );
  XOR2_X1 U1054 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n969) );
  XOR2_X1 U1055 ( .A(G1976), .B(G23), .Z(n963) );
  XOR2_X1 U1056 ( .A(G24), .B(KEYINPUT124), .Z(n961) );
  XNOR2_X1 U1057 ( .A(n961), .B(G1986), .ZN(n962) );
  NAND2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n966) );
  XOR2_X1 U1059 ( .A(KEYINPUT123), .B(G1971), .Z(n964) );
  XNOR2_X1 U1060 ( .A(G22), .B(n964), .ZN(n965) );
  NOR2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1062 ( .A(n967), .B(KEYINPUT58), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(n969), .B(n968), .ZN(n973) );
  XNOR2_X1 U1064 ( .A(G1961), .B(G5), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(G1966), .B(G21), .ZN(n970) );
  NOR2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1069 ( .A(KEYINPUT127), .B(n976), .Z(n977) );
  XNOR2_X1 U1070 ( .A(KEYINPUT61), .B(n977), .ZN(n978) );
  NAND2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n1035) );
  INV_X1 U1073 ( .A(KEYINPUT55), .ZN(n1007) );
  XOR2_X1 U1074 ( .A(G2090), .B(G162), .Z(n982) );
  NOR2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1076 ( .A(KEYINPUT111), .B(n984), .ZN(n985) );
  XNOR2_X1 U1077 ( .A(n985), .B(KEYINPUT51), .ZN(n1000) );
  XOR2_X1 U1078 ( .A(G160), .B(G2084), .Z(n986) );
  XNOR2_X1 U1079 ( .A(KEYINPUT110), .B(n986), .ZN(n987) );
  NOR2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n996) );
  XOR2_X1 U1081 ( .A(G2072), .B(n989), .Z(n991) );
  XOR2_X1 U1082 ( .A(G164), .B(G2078), .Z(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n992) );
  XOR2_X1 U1084 ( .A(KEYINPUT50), .B(n992), .Z(n993) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  NAND2_X1 U1090 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1091 ( .A(KEYINPUT52), .B(n1005), .Z(n1006) );
  NAND2_X1 U1092 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1093 ( .A1(n1008), .A2(G29), .ZN(n1033) );
  XNOR2_X1 U1094 ( .A(G1996), .B(G32), .ZN(n1010) );
  XNOR2_X1 U1095 ( .A(G2067), .B(G26), .ZN(n1009) );
  NOR2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1015) );
  XNOR2_X1 U1097 ( .A(G2072), .B(G33), .ZN(n1013) );
  XNOR2_X1 U1098 ( .A(G27), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1100 ( .A1(n1015), .A2(n1014), .ZN(n1019) );
  XOR2_X1 U1101 ( .A(G1991), .B(G25), .Z(n1016) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(G28), .ZN(n1017) );
  XNOR2_X1 U1103 ( .A(KEYINPUT112), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1105 ( .A(KEYINPUT53), .B(n1020), .Z(n1024) );
  XNOR2_X1 U1106 ( .A(KEYINPUT54), .B(G34), .ZN(n1021) );
  XNOR2_X1 U1107 ( .A(n1021), .B(KEYINPUT113), .ZN(n1022) );
  XNOR2_X1 U1108 ( .A(G2084), .B(n1022), .ZN(n1023) );
  NAND2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1026) );
  XNOR2_X1 U1110 ( .A(G35), .B(G2090), .ZN(n1025) );
  NOR2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1112 ( .A(KEYINPUT55), .B(n1027), .ZN(n1029) );
  INV_X1 U1113 ( .A(G29), .ZN(n1028) );
  NAND2_X1 U1114 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1115 ( .A1(n1030), .A2(G11), .ZN(n1031) );
  XOR2_X1 U1116 ( .A(KEYINPUT114), .B(n1031), .Z(n1032) );
  NAND2_X1 U1117 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NOR2_X1 U1118 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XNOR2_X1 U1119 ( .A(n1036), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1120 ( .A(G311), .ZN(G150) );
endmodule

