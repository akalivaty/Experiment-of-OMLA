//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 1 0 1 0 0 1 0 1 0 0 1 1 0 0 1 1 0 1 0 0 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1285,
    new_n1286, new_n1287, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  XOR2_X1   g0008(.A(KEYINPUT67), .B(G244), .Z(new_n209));
  AND2_X1   g0009(.A1(new_n209), .A2(G77), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G107), .A2(G264), .ZN(new_n214));
  NAND4_X1  g0014(.A1(new_n211), .A2(new_n212), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n208), .B1(new_n210), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(KEYINPUT1), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT68), .Z(new_n218));
  NAND2_X1  g0018(.A1(new_n202), .A2(G50), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT66), .Z(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n221), .A2(new_n206), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT64), .ZN(new_n224));
  OR3_X1    g0024(.A1(new_n208), .A2(new_n224), .A3(G13), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n224), .B1(new_n208), .B2(G13), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT0), .ZN(new_n229));
  INV_X1    g0029(.A(KEYINPUT65), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n223), .B1(KEYINPUT1), .B2(new_n216), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n218), .B(new_n231), .C1(new_n230), .C2(new_n229), .ZN(G361));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT69), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G226), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT70), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  INV_X1    g0041(.A(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n238), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n244), .B(new_n245), .Z(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  AOI21_X1  g0050(.A(new_n221), .B1(G33), .B2(G41), .ZN(new_n251));
  INV_X1    g0051(.A(G41), .ZN(new_n252));
  INV_X1    g0052(.A(G45), .ZN(new_n253));
  AOI21_X1  g0053(.A(G1), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G274), .ZN(new_n256));
  AND2_X1   g0056(.A1(G1), .A2(G13), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n255), .A2(G232), .B1(new_n259), .B2(new_n254), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  INV_X1    g0061(.A(G87), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G1698), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT71), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT71), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G1698), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n265), .A2(new_n267), .A3(G223), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G226), .A2(G1698), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT80), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n271), .B1(new_n261), .B2(KEYINPUT3), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT3), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(KEYINPUT80), .A3(G33), .ZN(new_n275));
  AND3_X1   g0075(.A1(new_n272), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n263), .B1(new_n270), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n257), .A2(new_n258), .ZN(new_n278));
  OAI211_X1 g0078(.A(G179), .B(new_n260), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n259), .A2(new_n254), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G232), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n280), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n263), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT71), .B(G1698), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n286), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n272), .A2(new_n273), .A3(new_n275), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n285), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n284), .B1(new_n289), .B2(new_n251), .ZN(new_n290));
  INV_X1    g0090(.A(G169), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n279), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT81), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G58), .ZN(new_n295));
  INV_X1    g0095(.A(G68), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(G20), .B1(new_n297), .B2(new_n201), .ZN(new_n298));
  NOR2_X1   g0098(.A1(G20), .A2(G33), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G159), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT7), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n275), .A2(new_n273), .ZN(new_n304));
  AOI21_X1  g0104(.A(KEYINPUT80), .B1(new_n274), .B2(G33), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n303), .B(new_n206), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G68), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n303), .B1(new_n288), .B2(new_n206), .ZN(new_n308));
  OAI211_X1 g0108(.A(KEYINPUT16), .B(new_n302), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n221), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT16), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT3), .B(G33), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n303), .B1(new_n313), .B2(G20), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n274), .A2(G33), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n273), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n316), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n296), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n312), .B1(new_n318), .B2(new_n301), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n309), .A2(new_n311), .A3(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT72), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT72), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n323), .A2(new_n205), .A3(G13), .A4(G20), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n311), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n205), .A2(G20), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT8), .B(G58), .ZN(new_n330));
  NOR3_X1   g0130(.A1(new_n327), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n322), .A2(new_n324), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n331), .B1(new_n332), .B2(new_n330), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n320), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n260), .B1(new_n277), .B2(new_n278), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G169), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(KEYINPUT81), .A3(new_n279), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n294), .A2(new_n334), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT18), .ZN(new_n339));
  INV_X1    g0139(.A(G190), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n340), .B(new_n260), .C1(new_n277), .C2(new_n278), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(new_n290), .B2(G200), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(new_n320), .A3(new_n333), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT17), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n342), .A2(new_n320), .A3(new_n333), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT17), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT18), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n294), .A2(new_n334), .A3(new_n348), .A4(new_n337), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n339), .A2(new_n345), .A3(new_n347), .A4(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT73), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT10), .ZN(new_n353));
  OR2_X1    g0153(.A1(new_n352), .A2(KEYINPUT10), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n206), .A2(G33), .ZN(new_n355));
  INV_X1    g0155(.A(G150), .ZN(new_n356));
  INV_X1    g0156(.A(new_n299), .ZN(new_n357));
  OAI22_X1  g0157(.A1(new_n330), .A2(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G50), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n206), .B1(new_n201), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n311), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n328), .A2(G50), .ZN(new_n362));
  OAI221_X1 g0162(.A(new_n361), .B1(G50), .B2(new_n325), .C1(new_n327), .C2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT9), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n363), .B(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(G226), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n280), .B1(new_n282), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n313), .A2(G223), .A3(G1698), .ZN(new_n368));
  INV_X1    g0168(.A(G77), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n313), .A2(new_n286), .ZN(new_n370));
  INV_X1    g0170(.A(G222), .ZN(new_n371));
  OAI221_X1 g0171(.A(new_n368), .B1(new_n369), .B2(new_n313), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n367), .B1(new_n372), .B2(new_n251), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(G190), .ZN(new_n374));
  INV_X1    g0174(.A(G200), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n374), .B1(new_n375), .B2(new_n373), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n353), .B(new_n354), .C1(new_n365), .C2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n376), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n363), .B(KEYINPUT9), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n378), .A2(new_n379), .A3(new_n352), .A4(KEYINPUT10), .ZN(new_n380));
  AND2_X1   g0180(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n363), .B1(new_n373), .B2(G169), .ZN(new_n382));
  INV_X1    g0182(.A(G179), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n373), .A2(new_n383), .ZN(new_n384));
  OR2_X1    g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(G238), .A2(G1698), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n265), .A2(new_n267), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n313), .B(new_n386), .C1(new_n387), .C2(new_n283), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n388), .B(new_n251), .C1(G107), .C2(new_n313), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n255), .A2(new_n209), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n389), .A2(new_n280), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(G200), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(new_n340), .B2(new_n391), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n328), .A2(G77), .ZN(new_n394));
  OR2_X1    g0194(.A1(new_n327), .A2(new_n394), .ZN(new_n395));
  OAI22_X1  g0195(.A1(new_n330), .A2(new_n357), .B1(new_n206), .B2(new_n369), .ZN(new_n396));
  XNOR2_X1  g0196(.A(KEYINPUT15), .B(G87), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n397), .A2(new_n355), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n311), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n332), .A2(new_n369), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n395), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n393), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n391), .A2(new_n291), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n403), .B(new_n401), .C1(G179), .C2(new_n391), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n351), .A2(new_n381), .A3(new_n385), .A4(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n265), .A2(new_n267), .A3(G226), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G232), .A2(G1698), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n316), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G33), .A2(G97), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n251), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT13), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n255), .A2(G238), .B1(new_n259), .B2(new_n254), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT74), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT74), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n413), .A2(new_n418), .A3(new_n414), .A4(new_n415), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n413), .A2(new_n415), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT13), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n417), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(G200), .ZN(new_n423));
  XNOR2_X1  g0223(.A(new_n423), .B(KEYINPUT75), .ZN(new_n424));
  OAI22_X1  g0224(.A1(new_n355), .A2(new_n369), .B1(new_n206), .B2(G68), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT77), .ZN(new_n426));
  OAI22_X1  g0226(.A1(new_n425), .A2(new_n426), .B1(new_n359), .B2(new_n357), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n425), .A2(new_n426), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n311), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n429), .B(KEYINPUT11), .ZN(new_n430));
  NOR3_X1   g0230(.A1(new_n325), .A2(KEYINPUT12), .A3(G68), .ZN(new_n431));
  OR2_X1    g0231(.A1(new_n431), .A2(KEYINPUT78), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(KEYINPUT78), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT12), .B1(new_n325), .B2(G68), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n327), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n436), .A2(G68), .A3(new_n328), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n430), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n421), .A2(new_n416), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n440), .A2(KEYINPUT76), .A3(G190), .ZN(new_n441));
  AOI21_X1  g0241(.A(KEYINPUT76), .B1(new_n440), .B2(G190), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n439), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n424), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT79), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT14), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n422), .A2(new_n446), .A3(G169), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n421), .A2(G179), .A3(new_n416), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n446), .B1(new_n422), .B2(G169), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n445), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n422), .A2(G169), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT14), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n454), .A2(KEYINPUT79), .A3(new_n449), .A4(new_n447), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n439), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n407), .A2(new_n444), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT19), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n206), .B1(new_n411), .B2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(G97), .ZN(new_n460));
  INV_X1    g0260(.A(G107), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n262), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n206), .A2(G33), .A3(G97), .ZN(new_n463));
  AOI22_X1  g0263(.A1(new_n459), .A2(new_n462), .B1(new_n458), .B2(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n272), .A2(new_n275), .A3(new_n206), .A4(new_n273), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n464), .B1(new_n296), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n311), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n332), .A2(new_n397), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n205), .A2(G33), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n325), .A2(G87), .A3(new_n326), .A4(new_n469), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n467), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(G33), .A2(G116), .ZN(new_n472));
  INV_X1    g0272(.A(G244), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(new_n264), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n474), .B1(new_n286), .B2(G238), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n472), .B1(new_n475), .B2(new_n288), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n251), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n253), .A2(G1), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n259), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n205), .A2(G45), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n278), .A2(G250), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(KEYINPUT84), .B1(new_n477), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT84), .ZN(new_n485));
  AOI211_X1 g0285(.A(new_n485), .B(new_n482), .C1(new_n476), .C2(new_n251), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(KEYINPUT85), .B(new_n471), .C1(new_n487), .C2(new_n375), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT85), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n265), .A2(new_n267), .A3(G238), .ZN(new_n490));
  INV_X1    g0290(.A(new_n474), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n276), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n278), .B1(new_n493), .B2(new_n472), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n485), .B1(new_n494), .B2(new_n482), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n477), .A2(KEYINPUT84), .A3(new_n483), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n375), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n467), .A2(new_n468), .A3(new_n470), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n489), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n495), .A2(new_n496), .A3(G190), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n488), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n387), .A2(new_n473), .ZN(new_n502));
  AOI21_X1  g0302(.A(KEYINPUT4), .B1(new_n502), .B2(new_n276), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n315), .A2(new_n273), .A3(G250), .A4(G1698), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G283), .ZN(new_n505));
  NAND2_X1  g0305(.A1(KEYINPUT4), .A2(G244), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n504), .B(new_n505), .C1(new_n370), .C2(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n251), .B1(new_n503), .B2(new_n507), .ZN(new_n508));
  AND2_X1   g0308(.A1(KEYINPUT5), .A2(G41), .ZN(new_n509));
  NOR2_X1   g0309(.A1(KEYINPUT5), .A2(G41), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n478), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n511), .A2(G257), .A3(new_n278), .ZN(new_n512));
  XNOR2_X1  g0312(.A(KEYINPUT5), .B(G41), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n259), .A2(new_n478), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT82), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n512), .A2(new_n514), .A3(KEYINPUT82), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n517), .A2(KEYINPUT83), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT83), .B1(new_n517), .B2(new_n518), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n508), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G200), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n332), .A2(new_n460), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n325), .A2(G97), .A3(new_n326), .A4(new_n469), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n461), .B1(new_n314), .B2(new_n317), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  XNOR2_X1  g0327(.A(G97), .B(G107), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT6), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NOR3_X1   g0330(.A1(new_n529), .A2(new_n460), .A3(G107), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n533), .A2(G20), .B1(G77), .B2(new_n299), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n527), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n525), .B1(new_n535), .B2(new_n311), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n508), .A2(G190), .A3(new_n517), .A4(new_n518), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n383), .B(new_n508), .C1(new_n519), .C2(new_n520), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n508), .A2(new_n517), .A3(new_n518), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n531), .B1(new_n529), .B2(new_n528), .ZN(new_n541));
  OAI22_X1  g0341(.A1(new_n541), .A2(new_n206), .B1(new_n369), .B2(new_n357), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n311), .B1(new_n542), .B2(new_n526), .ZN(new_n543));
  INV_X1    g0343(.A(new_n525), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n540), .A2(new_n291), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n522), .A2(new_n538), .B1(new_n539), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n495), .A2(new_n496), .A3(new_n383), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n436), .A2(new_n469), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n468), .B(new_n467), .C1(new_n548), .C2(new_n397), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n547), .B(new_n549), .C1(new_n487), .C2(G169), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n501), .A2(new_n546), .A3(new_n550), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n286), .A2(G250), .B1(G257), .B2(G1698), .ZN(new_n552));
  OR2_X1    g0352(.A1(KEYINPUT90), .A2(G294), .ZN(new_n553));
  NAND2_X1  g0353(.A1(KEYINPUT90), .A2(G294), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI22_X1  g0355(.A1(new_n552), .A2(new_n288), .B1(new_n261), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n278), .B1(new_n556), .B2(KEYINPUT91), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT91), .ZN(new_n558));
  OAI221_X1 g0358(.A(new_n558), .B1(new_n261), .B2(new_n555), .C1(new_n552), .C2(new_n288), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n251), .B1(new_n478), .B2(new_n513), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n557), .A2(new_n559), .B1(G264), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n561), .A2(new_n340), .A3(new_n514), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(G264), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n261), .B1(new_n553), .B2(new_n554), .ZN(new_n564));
  NAND2_X1  g0364(.A1(G257), .A2(G1698), .ZN(new_n565));
  INV_X1    g0365(.A(G250), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n565), .B1(new_n387), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n564), .B1(new_n567), .B2(new_n276), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n251), .B1(new_n568), .B2(new_n558), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n556), .A2(KEYINPUT91), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n514), .B(new_n563), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n375), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n562), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g0373(.A(KEYINPUT88), .B(KEYINPUT24), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT22), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n206), .A2(G87), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n576), .B1(new_n316), .B2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT23), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(new_n206), .B2(G107), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n461), .A2(KEYINPUT23), .A3(G20), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n261), .A2(G20), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n580), .A2(new_n581), .B1(new_n582), .B2(G116), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(KEYINPUT22), .A2(G87), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n465), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n575), .B1(new_n584), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n578), .A2(new_n583), .ZN(new_n589));
  NOR3_X1   g0389(.A1(new_n589), .A2(new_n586), .A3(new_n574), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n311), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n436), .A2(G107), .A3(new_n469), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n332), .A2(new_n461), .ZN(new_n593));
  XNOR2_X1  g0393(.A(KEYINPUT89), .B(KEYINPUT25), .ZN(new_n594));
  XNOR2_X1  g0394(.A(new_n593), .B(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n591), .A2(new_n592), .A3(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n573), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n571), .A2(new_n291), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n286), .A2(G250), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n288), .B1(new_n600), .B2(new_n565), .ZN(new_n601));
  OAI21_X1  g0401(.A(KEYINPUT91), .B1(new_n601), .B2(new_n564), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n602), .A2(new_n559), .A3(new_n251), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n603), .A2(new_n383), .A3(new_n514), .A4(new_n563), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n599), .A2(new_n596), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n598), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n560), .A2(G270), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n514), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n316), .A2(G303), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n286), .A2(G257), .B1(G264), .B2(G1698), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n609), .B1(new_n610), .B2(new_n288), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n278), .B1(new_n611), .B2(KEYINPUT86), .ZN(new_n612));
  NAND2_X1  g0412(.A1(G264), .A2(G1698), .ZN(new_n613));
  INV_X1    g0413(.A(G257), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n613), .B1(new_n387), .B2(new_n614), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n615), .A2(new_n276), .B1(G303), .B2(new_n316), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT86), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n608), .B1(new_n612), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(G190), .ZN(new_n620));
  INV_X1    g0420(.A(G116), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n332), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n325), .A2(G116), .A3(new_n326), .A4(new_n469), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n310), .A2(new_n221), .B1(G20), .B2(new_n621), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n505), .B(new_n206), .C1(G33), .C2(new_n460), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n625), .A2(KEYINPUT20), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(KEYINPUT20), .B1(new_n625), .B2(new_n626), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n620), .B(new_n630), .C1(new_n375), .C2(new_n619), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT87), .ZN(new_n632));
  OAI21_X1  g0432(.A(G169), .B1(new_n624), .B2(new_n629), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n632), .B1(new_n619), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(KEYINPUT21), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT21), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n632), .B(new_n636), .C1(new_n619), .C2(new_n633), .ZN(new_n637));
  INV_X1    g0437(.A(new_n608), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n251), .B1(new_n616), .B2(new_n617), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n611), .A2(KEYINPUT86), .ZN(new_n640));
  OAI211_X1 g0440(.A(G179), .B(new_n638), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n641), .A2(new_n630), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n631), .A2(new_n635), .A3(new_n637), .A4(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n606), .A2(new_n643), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n457), .A2(new_n551), .A3(new_n644), .ZN(G372));
  NAND2_X1  g0445(.A1(new_n545), .A2(new_n539), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n501), .A2(new_n550), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(KEYINPUT26), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n605), .A2(new_n635), .A3(new_n637), .A4(new_n642), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT92), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n375), .B1(new_n477), .B2(new_n483), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n651), .B1(new_n652), .B2(new_n498), .ZN(new_n653));
  OAI21_X1  g0453(.A(G200), .B1(new_n494), .B2(new_n482), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n471), .A2(KEYINPUT92), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n653), .A2(new_n655), .A3(new_n500), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n291), .B1(new_n494), .B2(new_n482), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n547), .A2(new_n549), .A3(new_n657), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n650), .A2(new_n546), .A3(new_n598), .A4(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n656), .A2(new_n658), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(new_n646), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT26), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n649), .A2(new_n660), .A3(new_n658), .A4(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n457), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n381), .ZN(new_n667));
  AOI22_X1  g0467(.A1(new_n320), .A2(new_n333), .B1(new_n336), .B2(new_n279), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n668), .B(KEYINPUT18), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n414), .B1(new_n413), .B2(new_n415), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n671), .B1(KEYINPUT74), .B2(new_n416), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n291), .B1(new_n672), .B2(new_n419), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n448), .B1(new_n673), .B2(new_n446), .ZN(new_n674));
  AOI21_X1  g0474(.A(KEYINPUT79), .B1(new_n674), .B2(new_n454), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n450), .A2(new_n445), .A3(new_n451), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n438), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n405), .B1(new_n424), .B2(new_n443), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n343), .B(KEYINPUT17), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n670), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n666), .B(new_n385), .C1(new_n667), .C2(new_n681), .ZN(G369));
  INV_X1    g0482(.A(new_n606), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(G213), .A3(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(G343), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n683), .B1(new_n597), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n605), .B2(new_n690), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n635), .A2(new_n637), .A3(new_n642), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n630), .A2(new_n690), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n643), .B2(new_n694), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n692), .A2(new_n698), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n693), .A2(new_n690), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n683), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n605), .B2(new_n689), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n699), .A2(new_n703), .ZN(G399));
  INV_X1    g0504(.A(new_n227), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G41), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n462), .A2(G116), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n706), .A2(new_n205), .A3(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n219), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n709), .B1(new_n710), .B2(new_n706), .ZN(new_n711));
  XOR2_X1   g0511(.A(new_n711), .B(KEYINPUT28), .Z(new_n712));
  NAND2_X1  g0512(.A1(new_n648), .A2(new_n663), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n661), .A2(new_n646), .A3(new_n663), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n716), .A2(new_n658), .A3(new_n660), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT95), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n717), .A2(new_n718), .A3(KEYINPUT29), .A4(new_n690), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n714), .B1(new_n648), .B2(new_n663), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n659), .A2(new_n546), .A3(new_n598), .ZN(new_n721));
  AND4_X1   g0521(.A1(new_n605), .A2(new_n635), .A3(new_n637), .A4(new_n642), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n658), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OAI211_X1 g0523(.A(KEYINPUT29), .B(new_n690), .C1(new_n720), .C2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(KEYINPUT95), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT29), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n665), .A2(new_n690), .ZN(new_n727));
  AOI22_X1  g0527(.A1(new_n719), .A2(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(G330), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT31), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n690), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n619), .ZN(new_n733));
  AOI21_X1  g0533(.A(G179), .B1(new_n477), .B2(new_n483), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n521), .A2(new_n733), .A3(new_n571), .A4(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT30), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n540), .A2(new_n737), .ZN(new_n738));
  AOI211_X1 g0538(.A(new_n383), .B(new_n608), .C1(new_n612), .C2(new_n618), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n738), .A2(new_n739), .A3(new_n487), .A4(new_n561), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(KEYINPUT93), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n495), .A2(new_n603), .A3(new_n496), .A4(new_n563), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(new_n641), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT93), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n743), .A2(new_n744), .A3(new_n738), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n736), .B1(new_n741), .B2(new_n745), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n742), .A2(new_n641), .A3(new_n540), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(KEYINPUT30), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n732), .B1(new_n746), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n740), .A2(KEYINPUT93), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n744), .B1(new_n743), .B2(new_n738), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n735), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(KEYINPUT94), .B1(new_n747), .B2(KEYINPUT30), .ZN(new_n754));
  INV_X1    g0554(.A(new_n540), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n739), .A2(new_n487), .A3(new_n755), .A4(new_n561), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT94), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n756), .A2(new_n757), .A3(new_n737), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n689), .B1(new_n753), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n750), .B1(new_n760), .B2(new_n730), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n644), .A2(new_n551), .A3(new_n690), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n729), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n728), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n712), .B1(new_n764), .B2(G1), .ZN(G364));
  NAND2_X1  g0565(.A1(new_n206), .A2(G13), .ZN(new_n766));
  XOR2_X1   g0566(.A(new_n766), .B(KEYINPUT96), .Z(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n205), .B1(new_n768), .B2(G45), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n706), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n698), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(G330), .B2(new_n696), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n221), .B1(G20), .B2(new_n291), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n206), .A2(new_n383), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G200), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G190), .ZN(new_n777));
  NOR2_X1   g0577(.A1(KEYINPUT33), .A2(G317), .ZN(new_n778));
  AND2_X1   g0578(.A1(KEYINPUT33), .A2(G317), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n340), .A2(G179), .A3(G200), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n206), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n780), .B1(new_n555), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n206), .A2(G190), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n784), .A2(new_n383), .A3(new_n375), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(G190), .A2(G200), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n775), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI22_X1  g0589(.A1(G329), .A2(new_n786), .B1(new_n789), .B2(G311), .ZN(new_n790));
  OR3_X1    g0590(.A1(new_n375), .A2(KEYINPUT99), .A3(G179), .ZN(new_n791));
  OAI21_X1  g0591(.A(KEYINPUT99), .B1(new_n375), .B2(G179), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n206), .A2(new_n340), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G303), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n791), .A2(new_n792), .A3(new_n784), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G283), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n775), .A2(G190), .A3(new_n375), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n313), .B1(new_n801), .B2(G322), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n790), .A2(new_n796), .A3(new_n799), .A4(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n776), .A2(new_n340), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n783), .B(new_n803), .C1(G326), .C2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G159), .ZN(new_n806));
  OAI21_X1  g0606(.A(KEYINPUT32), .B1(new_n785), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n804), .ZN(new_n808));
  INV_X1    g0608(.A(new_n777), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n807), .B1(new_n808), .B2(new_n359), .C1(new_n296), .C2(new_n809), .ZN(new_n810));
  NOR3_X1   g0610(.A1(new_n785), .A2(KEYINPUT32), .A3(new_n806), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n782), .A2(new_n460), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n316), .B1(new_n789), .B2(G77), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n813), .B(new_n814), .C1(new_n295), .C2(new_n800), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n797), .A2(new_n461), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n794), .A2(new_n262), .ZN(new_n817));
  NOR4_X1   g0617(.A1(new_n810), .A2(new_n815), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n774), .B1(new_n805), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(new_n771), .ZN(new_n820));
  NOR2_X1   g0620(.A1(G13), .A2(G33), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(G20), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(new_n774), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n705), .A2(new_n316), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n825), .A2(G355), .B1(new_n621), .B2(new_n705), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n246), .A2(new_n253), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  OR2_X1    g0628(.A1(new_n828), .A2(KEYINPUT97), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n220), .A2(new_n253), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n828), .A2(KEYINPUT97), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n227), .A2(new_n288), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT98), .Z(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n826), .B1(new_n832), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n820), .B1(new_n824), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n823), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n837), .B1(new_n696), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n773), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(G396));
  AOI21_X1  g0641(.A(new_n402), .B1(new_n401), .B2(new_n689), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n842), .A2(new_n405), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n404), .A2(new_n689), .ZN(new_n844));
  OAI21_X1  g0644(.A(KEYINPUT101), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OR3_X1    g0645(.A1(new_n843), .A2(KEYINPUT101), .A3(new_n844), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n727), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT102), .ZN(new_n848));
  NOR3_X1   g0648(.A1(new_n402), .A2(new_n405), .A3(new_n689), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n665), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n763), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n851), .A2(new_n771), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n848), .A2(new_n763), .A3(new_n850), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n774), .A2(new_n821), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n771), .B1(G77), .B2(new_n856), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n801), .A2(G143), .B1(new_n789), .B2(G159), .ZN(new_n858));
  INV_X1    g0658(.A(G137), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n858), .B1(new_n808), .B2(new_n859), .C1(new_n356), .C2(new_n809), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT34), .ZN(new_n861));
  OR2_X1    g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n860), .A2(new_n861), .ZN(new_n863));
  INV_X1    g0663(.A(G132), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n276), .B1(new_n864), .B2(new_n785), .ZN(new_n865));
  INV_X1    g0665(.A(new_n782), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n865), .B1(G58), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n797), .A2(new_n296), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n868), .B1(G50), .B2(new_n795), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n862), .A2(new_n863), .A3(new_n867), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n798), .A2(G87), .ZN(new_n871));
  INV_X1    g0671(.A(G311), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n871), .B1(new_n872), .B2(new_n785), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n873), .B(KEYINPUT100), .ZN(new_n874));
  INV_X1    g0674(.A(G283), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n809), .A2(new_n875), .ZN(new_n876));
  AOI211_X1 g0676(.A(new_n812), .B(new_n876), .C1(G303), .C2(new_n804), .ZN(new_n877));
  INV_X1    g0677(.A(G294), .ZN(new_n878));
  OAI221_X1 g0678(.A(new_n316), .B1(new_n788), .B2(new_n621), .C1(new_n878), .C2(new_n800), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(G107), .B2(new_n795), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n874), .A2(new_n877), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n870), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n857), .B1(new_n882), .B2(new_n774), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n843), .A2(new_n844), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n883), .B1(new_n884), .B2(new_n822), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n854), .A2(new_n885), .ZN(G384));
  OAI211_X1 g0686(.A(G116), .B(new_n222), .C1(new_n533), .C2(KEYINPUT35), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n887), .A2(KEYINPUT103), .B1(KEYINPUT35), .B2(new_n533), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(KEYINPUT103), .B2(new_n887), .ZN(new_n889));
  XOR2_X1   g0689(.A(new_n889), .B(KEYINPUT36), .Z(new_n890));
  OR3_X1    g0690(.A1(new_n219), .A2(new_n369), .A3(new_n297), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n359), .A2(G68), .ZN(new_n892));
  AOI211_X1 g0692(.A(new_n205), .B(G13), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n844), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n850), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n309), .A2(new_n311), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT7), .B1(new_n276), .B2(G20), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n898), .A2(G68), .A3(new_n306), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT16), .B1(new_n899), .B2(new_n302), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n333), .B1(new_n897), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n687), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n350), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n901), .A2(new_n292), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n903), .A2(new_n906), .A3(new_n343), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(KEYINPUT37), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n687), .B1(new_n320), .B2(new_n333), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n346), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT37), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n910), .A2(new_n911), .A3(new_n338), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n905), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT38), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n905), .A2(new_n913), .A3(KEYINPUT38), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n444), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n438), .A2(new_n689), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n677), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n920), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n456), .B2(new_n444), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n896), .A2(new_n918), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n670), .A2(new_n687), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT104), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT39), .ZN(new_n930));
  NOR3_X1   g0730(.A1(new_n346), .A2(new_n668), .A3(new_n909), .ZN(new_n931));
  OAI21_X1  g0731(.A(KEYINPUT106), .B1(new_n931), .B2(new_n911), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT106), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n334), .A2(new_n902), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n343), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n933), .B(KEYINPUT37), .C1(new_n935), .C2(new_n668), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n932), .A2(new_n912), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n669), .A2(new_n680), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n909), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT38), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  AND3_X1   g0740(.A1(new_n905), .A2(KEYINPUT38), .A3(new_n913), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n930), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n438), .B(new_n690), .C1(new_n675), .C2(new_n676), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT105), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n456), .A2(KEYINPUT105), .A3(new_n690), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n916), .A2(KEYINPUT39), .A3(new_n917), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n942), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n925), .A2(KEYINPUT104), .A3(new_n926), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n929), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n385), .B1(new_n681), .B2(new_n667), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(new_n728), .B2(new_n457), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n951), .B(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n731), .B1(new_n753), .B2(new_n759), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n756), .A2(new_n757), .A3(new_n737), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n757), .B1(new_n756), .B2(new_n737), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n690), .B1(new_n958), .B2(new_n746), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n762), .B(new_n955), .C1(new_n959), .C2(KEYINPUT31), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n924), .A2(new_n918), .A3(new_n960), .A4(new_n884), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT40), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n937), .A2(new_n939), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n915), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n962), .B1(new_n965), .B2(new_n917), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n966), .A2(new_n884), .A3(new_n924), .A4(new_n960), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n963), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n457), .A2(new_n960), .ZN(new_n969));
  OAI21_X1  g0769(.A(G330), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(new_n968), .B2(new_n969), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n954), .A2(new_n971), .B1(new_n205), .B2(new_n768), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n954), .A2(new_n971), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n894), .B1(new_n972), .B2(new_n973), .ZN(G367));
  NAND2_X1  g0774(.A1(new_n498), .A2(new_n689), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n659), .A2(new_n975), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n976), .A2(KEYINPUT107), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(KEYINPUT107), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n977), .B(new_n978), .C1(new_n658), .C2(new_n975), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n823), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n835), .A2(new_n242), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n824), .B1(new_n227), .B2(new_n397), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n771), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(G317), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n985), .A2(new_n785), .B1(new_n788), .B2(new_n875), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(G303), .B2(new_n801), .ZN(new_n987));
  INV_X1    g0787(.A(new_n555), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n276), .B1(new_n777), .B2(new_n988), .ZN(new_n989));
  AOI22_X1  g0789(.A1(G107), .A2(new_n866), .B1(new_n804), .B2(G311), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n798), .A2(G97), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n987), .A2(new_n989), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n794), .A2(new_n621), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT46), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n866), .A2(G68), .ZN(new_n995));
  INV_X1    g0795(.A(G143), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n995), .B1(new_n808), .B2(new_n996), .C1(new_n806), .C2(new_n809), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n801), .A2(G150), .B1(new_n789), .B2(G50), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n795), .A2(G58), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n798), .A2(G77), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n316), .B1(new_n786), .B2(G137), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n992), .A2(new_n994), .B1(new_n997), .B2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT47), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n984), .B1(new_n1004), .B2(new_n774), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n981), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n546), .B1(new_n536), .B2(new_n690), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n647), .A2(new_n689), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n702), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT45), .ZN(new_n1011));
  XOR2_X1   g0811(.A(KEYINPUT110), .B(KEYINPUT44), .Z(new_n1012));
  NAND3_X1  g0812(.A1(new_n702), .A2(new_n1009), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1012), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1009), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1014), .B1(new_n703), .B2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1011), .A2(new_n1013), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n699), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1011), .A2(new_n699), .A3(new_n1013), .A4(new_n1016), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n701), .B1(new_n692), .B2(new_n700), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(new_n698), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n764), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1025));
  XOR2_X1   g0825(.A(KEYINPUT109), .B(KEYINPUT41), .Z(new_n1026));
  XNOR2_X1  g0826(.A(new_n706), .B(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n770), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1009), .A2(new_n701), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT42), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n605), .B1(new_n522), .B2(new_n538), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n690), .B1(new_n1032), .B2(new_n647), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  XOR2_X1   g0834(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n1035));
  NAND2_X1  g0835(.A1(new_n980), .A2(new_n1035), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1034), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT43), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1036), .B1(new_n1039), .B2(new_n980), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1037), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n699), .A2(new_n1009), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1041), .B(new_n1042), .Z(new_n1043));
  OAI21_X1  g0843(.A(new_n1006), .B1(new_n1029), .B2(new_n1043), .ZN(G387));
  OAI21_X1  g0844(.A(new_n1024), .B1(new_n728), .B2(new_n763), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n764), .A2(new_n1023), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1045), .A2(new_n706), .A3(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n692), .A2(new_n838), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n237), .A2(G45), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT111), .Z(new_n1050));
  NOR2_X1   g0850(.A1(new_n330), .A2(G50), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT50), .ZN(new_n1052));
  AOI211_X1 g0852(.A(G45), .B(new_n708), .C1(G68), .C2(G77), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n835), .B(new_n1050), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n825), .A2(new_n708), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(G107), .B2(new_n227), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n824), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n276), .B1(G326), .B2(new_n786), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n794), .A2(new_n555), .B1(new_n875), .B2(new_n782), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n801), .A2(G317), .B1(new_n789), .B2(G303), .ZN(new_n1060));
  INV_X1    g0860(.A(G322), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1060), .B1(new_n808), .B2(new_n1061), .C1(new_n872), .C2(new_n809), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT48), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1059), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n1063), .B2(new_n1062), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT49), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1058), .B1(new_n621), .B2(new_n797), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n1066), .B2(new_n1065), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n801), .A2(G50), .B1(new_n789), .B2(G68), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1069), .B(new_n991), .C1(new_n356), .C2(new_n785), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n276), .B1(new_n808), .B2(new_n806), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n782), .A2(new_n397), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n809), .B2(new_n330), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n794), .A2(new_n369), .ZN(new_n1074));
  NOR4_X1   g0874(.A1(new_n1070), .A2(new_n1071), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n774), .B1(new_n1068), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1057), .A2(new_n771), .A3(new_n1076), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1047), .B1(new_n769), .B2(new_n1024), .C1(new_n1048), .C2(new_n1077), .ZN(G393));
  OR2_X1    g0878(.A1(new_n1021), .A2(new_n1046), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1021), .A2(new_n1046), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1079), .A2(new_n706), .A3(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1019), .A2(new_n770), .A3(new_n1020), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n835), .A2(new_n249), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n824), .B1(new_n227), .B2(new_n460), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n771), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n316), .B1(new_n788), .B2(new_n878), .C1(new_n782), .C2(new_n621), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n816), .B(new_n1086), .C1(G303), .C2(new_n777), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(G317), .A2(new_n804), .B1(new_n801), .B2(G311), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1088), .B(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n794), .A2(new_n875), .B1(new_n1061), .B2(new_n785), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT114), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(G77), .A2(new_n866), .B1(new_n777), .B2(G50), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n996), .A2(new_n785), .B1(new_n788), .B2(new_n330), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1095), .A2(new_n288), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n795), .A2(G68), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1094), .A2(new_n1096), .A3(new_n871), .A4(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(G150), .A2(new_n804), .B1(new_n801), .B2(G159), .ZN(new_n1099));
  XOR2_X1   g0899(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n1100));
  XNOR2_X1  g0900(.A(new_n1099), .B(new_n1100), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n1091), .A2(new_n1093), .B1(new_n1098), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1085), .B1(new_n1102), .B2(new_n774), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n1015), .B2(new_n838), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1081), .A2(new_n1082), .A3(new_n1104), .ZN(G390));
  INV_X1    g0905(.A(new_n843), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n690), .B(new_n1106), .C1(new_n720), .C2(new_n723), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n895), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n924), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT115), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n947), .A2(new_n1110), .B1(new_n965), .B2(new_n917), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n945), .A2(KEYINPUT115), .A3(new_n946), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1109), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n942), .A2(new_n948), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n850), .A2(new_n895), .B1(new_n921), .B2(new_n923), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1114), .B1(new_n1115), .B2(new_n947), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n731), .B1(new_n753), .B2(new_n748), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n762), .B(new_n1117), .C1(new_n959), .C2(KEYINPUT31), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n924), .A2(new_n1118), .A3(G330), .A4(new_n884), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1113), .A2(new_n1116), .A3(new_n1119), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n456), .A2(KEYINPUT105), .A3(new_n690), .ZN(new_n1121));
  AOI21_X1  g0921(.A(KEYINPUT105), .B1(new_n456), .B2(new_n690), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1110), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(KEYINPUT37), .B1(new_n935), .B2(new_n668), .ZN(new_n1124));
  AND2_X1   g0924(.A1(new_n338), .A2(new_n911), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n1124), .A2(KEYINPUT106), .B1(new_n1125), .B2(new_n910), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1126), .A2(new_n936), .B1(new_n909), .B2(new_n938), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n917), .B1(new_n1127), .B2(KEYINPUT38), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n1123), .A2(new_n1128), .A3(new_n1112), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n947), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n921), .A2(new_n923), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n844), .B1(new_n665), .B2(new_n849), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1130), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1129), .A2(new_n1109), .B1(new_n1133), .B2(new_n1114), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n924), .A2(new_n960), .A3(G330), .A4(new_n884), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1120), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1114), .A2(new_n821), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n855), .A2(new_n330), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n771), .A2(new_n1139), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n1140), .B(KEYINPUT117), .Z(new_n1141));
  INV_X1    g0941(.A(new_n774), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(G159), .A2(new_n866), .B1(new_n777), .B2(G137), .ZN(new_n1143));
  INV_X1    g0943(.A(G128), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1143), .B1(new_n1144), .B2(new_n808), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(KEYINPUT54), .B(G143), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n800), .A2(new_n864), .B1(new_n788), .B2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n797), .A2(new_n359), .ZN(new_n1148));
  INV_X1    g0948(.A(G125), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n313), .B1(new_n785), .B2(new_n1149), .ZN(new_n1150));
  NOR4_X1   g0950(.A1(new_n1145), .A2(new_n1147), .A3(new_n1148), .A4(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n794), .A2(new_n356), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT53), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n809), .A2(new_n461), .B1(new_n808), .B2(new_n875), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n316), .B1(new_n788), .B2(new_n460), .C1(new_n878), .C2(new_n785), .ZN(new_n1155));
  NOR4_X1   g0955(.A1(new_n1154), .A2(new_n817), .A3(new_n868), .A4(new_n1155), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n782), .A2(new_n369), .B1(new_n800), .B2(new_n621), .ZN(new_n1157));
  XOR2_X1   g0957(.A(new_n1157), .B(KEYINPUT118), .Z(new_n1158));
  AOI22_X1  g0958(.A1(new_n1151), .A2(new_n1153), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1141), .B1(new_n1142), .B2(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT119), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n1137), .A2(new_n770), .B1(new_n1138), .B2(new_n1161), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n457), .A2(new_n960), .A3(G330), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n846), .A2(new_n845), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n960), .A2(G330), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n1131), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1108), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n1167), .A2(new_n1119), .A3(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1118), .A2(G330), .A3(new_n884), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n1131), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1132), .B1(new_n1171), .B2(new_n1135), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n953), .B(new_n1164), .C1(new_n1169), .C2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n1136), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n924), .B1(new_n763), .B2(new_n884), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1135), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n896), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1167), .A2(new_n1119), .A3(new_n1168), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n952), .B(new_n1163), .C1(new_n728), .C2(new_n457), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n896), .A2(new_n924), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n1181), .A2(new_n1130), .B1(new_n942), .B2(new_n948), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1123), .A2(new_n1128), .A3(new_n1112), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n1107), .A2(new_n895), .B1(new_n921), .B2(new_n923), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1176), .B1(new_n1182), .B2(new_n1185), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1179), .A2(new_n1180), .A3(new_n1186), .A4(new_n1120), .ZN(new_n1187));
  AND4_X1   g0987(.A1(KEYINPUT116), .A2(new_n1174), .A3(new_n706), .A4(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n706), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n1173), .B2(new_n1136), .ZN(new_n1190));
  AOI21_X1  g0990(.A(KEYINPUT116), .B1(new_n1190), .B2(new_n1187), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1162), .B1(new_n1188), .B2(new_n1191), .ZN(G378));
  INV_X1    g0992(.A(KEYINPUT57), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n1187), .B2(new_n1180), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT122), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n963), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1128), .A2(KEYINPUT40), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n924), .A2(new_n960), .A3(new_n884), .ZN(new_n1198));
  OAI21_X1  g0998(.A(G330), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1195), .B1(new_n1196), .B2(new_n1199), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n963), .A2(new_n967), .A3(KEYINPUT122), .A4(G330), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n381), .A2(new_n385), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n363), .A2(new_n902), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT121), .Z(new_n1204));
  XNOR2_X1  g1004(.A(new_n1202), .B(new_n1204), .ZN(new_n1205));
  XOR2_X1   g1005(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1206));
  XNOR2_X1  g1006(.A(new_n1205), .B(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1200), .A2(new_n1201), .A3(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1207), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1209), .B(new_n1195), .C1(new_n1196), .C2(new_n1199), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n951), .B1(new_n1208), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1201), .A2(new_n1207), .ZN(new_n1212));
  AND3_X1   g1012(.A1(new_n924), .A2(new_n960), .A3(new_n884), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n729), .B1(new_n1213), .B2(new_n966), .ZN(new_n1214));
  AOI21_X1  g1014(.A(KEYINPUT122), .B1(new_n1214), .B2(new_n963), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n951), .B(new_n1210), .C1(new_n1212), .C2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1194), .B1(new_n1211), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n706), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1210), .B1(new_n1212), .B2(new_n1215), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n951), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n1216), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1187), .A2(new_n1180), .ZN(new_n1224));
  AOI21_X1  g1024(.A(KEYINPUT57), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  OR2_X1    g1025(.A1(new_n1219), .A2(new_n1225), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1209), .A2(new_n822), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n800), .A2(new_n1144), .B1(new_n788), .B2(new_n859), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(G132), .B2(new_n777), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(G150), .A2(new_n866), .B1(new_n804), .B2(G125), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1229), .B(new_n1230), .C1(new_n794), .C2(new_n1146), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1231), .A2(KEYINPUT59), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(KEYINPUT59), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n798), .A2(G159), .ZN(new_n1234));
  AOI211_X1 g1034(.A(G33), .B(G41), .C1(new_n786), .C2(G124), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1232), .A2(new_n1233), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n798), .A2(G58), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(new_n1237), .B(KEYINPUT120), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n800), .A2(new_n461), .B1(new_n785), .B2(new_n875), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n252), .B1(new_n788), .B2(new_n397), .ZN(new_n1241));
  NOR3_X1   g1041(.A1(new_n1074), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(G97), .A2(new_n777), .B1(new_n804), .B2(G116), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1242), .A2(new_n288), .A3(new_n995), .A4(new_n1243), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1239), .A2(new_n1244), .ZN(new_n1245));
  OR2_X1    g1045(.A1(new_n1245), .A2(KEYINPUT58), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(KEYINPUT58), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n252), .B1(new_n288), .B2(new_n261), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n359), .ZN(new_n1249));
  AND4_X1   g1049(.A1(new_n1236), .A2(new_n1246), .A3(new_n1247), .A4(new_n1249), .ZN(new_n1250));
  OAI221_X1 g1050(.A(new_n771), .B1(G50), .B2(new_n856), .C1(new_n1250), .C2(new_n1142), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1227), .A2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n1223), .B2(new_n770), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1226), .A2(new_n1253), .ZN(G375));
  NAND2_X1  g1054(.A1(new_n953), .A2(new_n1164), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1255), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1256), .A2(new_n1028), .A3(new_n1173), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1131), .A2(new_n821), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n771), .B1(G68), .B2(new_n856), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n800), .A2(new_n859), .B1(new_n785), .B2(new_n1144), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(G150), .B2(new_n789), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n288), .B1(new_n804), .B2(G132), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1146), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(G50), .A2(new_n866), .B1(new_n777), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n795), .A2(G159), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1261), .A2(new_n1262), .A3(new_n1264), .A4(new_n1265), .ZN(new_n1266));
  OAI221_X1 g1066(.A(new_n1072), .B1(new_n808), .B2(new_n878), .C1(new_n621), .C2(new_n809), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(G303), .A2(new_n786), .B1(new_n789), .B2(G107), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n795), .A2(G97), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n313), .B1(new_n801), .B2(G283), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1268), .A2(new_n1269), .A3(new_n1000), .A4(new_n1270), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n1239), .A2(new_n1266), .B1(new_n1267), .B2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1259), .B1(new_n1272), .B2(new_n774), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n1179), .A2(new_n770), .B1(new_n1258), .B2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1257), .A2(new_n1274), .ZN(G381));
  AND3_X1   g1075(.A1(new_n1081), .A2(new_n1082), .A3(new_n1104), .ZN(new_n1276));
  INV_X1    g1076(.A(G384), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  NOR4_X1   g1078(.A1(new_n1278), .A2(G396), .A3(G393), .A4(G381), .ZN(new_n1279));
  INV_X1    g1079(.A(G375), .ZN(new_n1280));
  INV_X1    g1080(.A(G387), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1190), .A2(new_n1187), .ZN(new_n1282));
  AND2_X1   g1082(.A1(new_n1282), .A2(new_n1162), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1279), .A2(new_n1280), .A3(new_n1281), .A4(new_n1283), .ZN(G407));
  NAND4_X1  g1084(.A1(new_n1280), .A2(G213), .A3(new_n688), .A4(new_n1283), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(G407), .A2(new_n1285), .A3(G213), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT123), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(new_n1286), .B(new_n1287), .ZN(G409));
  AND2_X1   g1088(.A1(new_n1276), .A2(G387), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1276), .A2(G387), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(G393), .A2(G396), .ZN(new_n1291));
  AND2_X1   g1091(.A1(G393), .A2(G396), .ZN(new_n1292));
  OAI22_X1  g1092(.A1(new_n1289), .A2(new_n1290), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1281), .A2(G390), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1292), .A2(new_n1291), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1276), .A2(G387), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1294), .A2(new_n1295), .A3(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT61), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1293), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1256), .A2(KEYINPUT125), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT60), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1256), .A2(KEYINPUT125), .A3(KEYINPUT60), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1173), .A2(new_n706), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1304), .A2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1307), .A2(G384), .A3(new_n1274), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1305), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1274), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1277), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT63), .ZN(new_n1314));
  NOR3_X1   g1114(.A1(new_n1309), .A2(new_n1313), .A3(new_n1314), .ZN(new_n1315));
  OAI211_X1 g1115(.A(G378), .B(new_n1253), .C1(new_n1219), .C2(new_n1225), .ZN(new_n1316));
  OAI211_X1 g1116(.A(new_n1028), .B(new_n1224), .C1(new_n1217), .C2(new_n1211), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n770), .B1(new_n1217), .B2(new_n1211), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1252), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1317), .A2(new_n1318), .A3(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n1283), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1316), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n688), .A2(G213), .ZN(new_n1323));
  AND2_X1   g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1299), .B1(new_n1315), .B2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT124), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1322), .A2(new_n1326), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1316), .A2(KEYINPUT124), .A3(new_n1321), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1327), .A2(new_n1323), .A3(new_n1328), .ZN(new_n1329));
  AND3_X1   g1129(.A1(new_n688), .A2(G213), .A3(G2897), .ZN(new_n1330));
  AND3_X1   g1130(.A1(new_n1308), .A2(new_n1312), .A3(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1330), .B1(new_n1308), .B2(new_n1312), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1329), .B1(new_n1331), .B2(new_n1332), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1309), .A2(new_n1313), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1327), .A2(new_n1323), .A3(new_n1334), .A4(new_n1328), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1335), .A2(new_n1314), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1325), .A2(new_n1333), .A3(new_n1336), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1298), .B1(new_n1324), .B2(new_n1338), .ZN(new_n1339));
  XNOR2_X1  g1139(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1335), .A2(new_n1340), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1324), .A2(KEYINPUT62), .A3(new_n1334), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1339), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1343));
  AND2_X1   g1143(.A1(new_n1293), .A2(new_n1297), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1337), .B1(new_n1343), .B2(new_n1344), .ZN(G405));
  NAND2_X1  g1145(.A1(G375), .A2(new_n1283), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1346), .A2(new_n1316), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1334), .A2(KEYINPUT127), .ZN(new_n1348));
  INV_X1    g1148(.A(KEYINPUT127), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1349), .B1(new_n1309), .B2(new_n1313), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1347), .A2(new_n1348), .A3(new_n1350), .ZN(new_n1351));
  NAND4_X1  g1151(.A1(new_n1346), .A2(KEYINPUT127), .A3(new_n1334), .A4(new_n1316), .ZN(new_n1352));
  AND3_X1   g1152(.A1(new_n1351), .A2(new_n1344), .A3(new_n1352), .ZN(new_n1353));
  AOI21_X1  g1153(.A(new_n1344), .B1(new_n1351), .B2(new_n1352), .ZN(new_n1354));
  NOR2_X1   g1154(.A1(new_n1353), .A2(new_n1354), .ZN(G402));
endmodule


