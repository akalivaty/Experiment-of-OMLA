//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 1 1 0 0 0 1 1 0 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 0 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n846, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n202));
  INV_X1    g001(.A(G127gat), .ZN(new_n203));
  INV_X1    g002(.A(G134gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT70), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT70), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G134gat), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n203), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n203), .A2(KEYINPUT71), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT71), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G127gat), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n204), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n202), .B1(new_n208), .B2(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n206), .A2(G134gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n204), .A2(KEYINPUT70), .ZN(new_n215));
  OAI21_X1  g014(.A(G127gat), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n210), .A2(G127gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n203), .A2(KEYINPUT71), .ZN(new_n218));
  OAI21_X1  g017(.A(G134gat), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n216), .A2(new_n219), .A3(KEYINPUT72), .ZN(new_n220));
  XOR2_X1   g019(.A(G113gat), .B(G120gat), .Z(new_n221));
  INV_X1    g020(.A(KEYINPUT1), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n213), .A2(new_n220), .A3(new_n223), .ZN(new_n224));
  XOR2_X1   g023(.A(G127gat), .B(G134gat), .Z(new_n225));
  NAND3_X1  g024(.A1(new_n221), .A2(new_n225), .A3(new_n222), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  AND2_X1   g026(.A1(G155gat), .A2(G162gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(G155gat), .A2(G162gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G141gat), .B(G148gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(G155gat), .A2(G162gat), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n232), .A2(KEYINPUT2), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n230), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(G141gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(G148gat), .ZN(new_n236));
  INV_X1    g035(.A(G148gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(G141gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(G155gat), .B(G162gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n232), .A2(KEYINPUT2), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n234), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT4), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(G225gat), .A2(G233gat), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n243), .B1(new_n224), .B2(new_n226), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT4), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n234), .A2(new_n242), .A3(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT76), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n234), .A2(new_n242), .A3(KEYINPUT76), .A4(new_n251), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n243), .A2(KEYINPUT3), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n256), .A2(new_n226), .A3(new_n224), .A4(new_n257), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n247), .A2(new_n248), .A3(new_n250), .A4(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n248), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n224), .A2(new_n243), .A3(new_n226), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n260), .B1(new_n261), .B2(new_n249), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT77), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT78), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n265), .B1(new_n259), .B2(KEYINPUT5), .ZN(new_n266));
  OAI21_X1  g065(.A(KEYINPUT5), .B1(new_n262), .B2(KEYINPUT77), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n264), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n249), .B(new_n246), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT5), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n270), .A2(new_n271), .A3(new_n248), .A4(new_n258), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n259), .A2(new_n263), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n272), .B(new_n265), .C1(new_n273), .C2(new_n267), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(KEYINPUT0), .B(G57gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(G85gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(G1gat), .B(G29gat), .ZN(new_n278));
  XOR2_X1   g077(.A(new_n277), .B(new_n278), .Z(new_n279));
  NAND2_X1  g078(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n281));
  INV_X1    g080(.A(new_n279), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n269), .A2(new_n274), .A3(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n280), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n269), .A2(new_n274), .A3(KEYINPUT6), .A4(new_n282), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OR2_X1    g085(.A1(G197gat), .A2(G204gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(G197gat), .A2(G204gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT75), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n287), .A2(KEYINPUT75), .A3(new_n288), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT22), .ZN(new_n294));
  XOR2_X1   g093(.A(G211gat), .B(G218gat), .Z(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n295), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT22), .ZN(new_n298));
  INV_X1    g097(.A(G211gat), .ZN(new_n299));
  INV_X1    g098(.A(G218gat), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n293), .A2(new_n297), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n296), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G226gat), .A2(G233gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT67), .ZN(new_n307));
  NOR2_X1   g106(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n310));
  OR2_X1    g109(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n312));
  AOI22_X1  g111(.A1(new_n309), .A2(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G183gat), .A2(G190gat), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT24), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n314), .B(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n307), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(G169gat), .A2(G176gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT23), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n318), .A2(KEYINPUT64), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT64), .ZN(new_n321));
  OAI22_X1  g120(.A1(new_n321), .A2(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n321), .A2(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n310), .ZN(new_n326));
  INV_X1    g125(.A(new_n312), .ZN(new_n327));
  NOR2_X1   g126(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n328));
  OAI22_X1  g127(.A1(new_n308), .A2(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n314), .B(KEYINPUT24), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n329), .A2(new_n330), .A3(KEYINPUT67), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n317), .A2(new_n325), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT25), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n334), .B(KEYINPUT68), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT26), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n318), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT69), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n337), .A2(new_n338), .B1(G169gat), .B2(G176gat), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n335), .B(new_n339), .C1(new_n338), .C2(new_n337), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n326), .A2(new_n308), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT28), .ZN(new_n343));
  AND3_X1   g142(.A1(new_n311), .A2(KEYINPUT27), .A3(new_n312), .ZN(new_n344));
  NOR2_X1   g143(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n342), .B(new_n343), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  XOR2_X1   g145(.A(KEYINPUT27), .B(G183gat), .Z(new_n347));
  OAI21_X1  g146(.A(KEYINPUT28), .B1(new_n347), .B2(new_n341), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n340), .A2(new_n346), .A3(new_n348), .A4(new_n314), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT25), .ZN(new_n350));
  NOR2_X1   g149(.A1(G183gat), .A2(G190gat), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n350), .B1(new_n316), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n323), .A2(new_n324), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n333), .A2(new_n349), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT29), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n306), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n354), .B1(new_n332), .B2(KEYINPUT25), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n305), .B1(new_n359), .B2(new_n349), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n304), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(G8gat), .B(G36gat), .ZN(new_n362));
  INV_X1    g161(.A(G64gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n362), .B(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(G92gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n356), .A2(new_n306), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT29), .B1(new_n359), .B2(new_n349), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n368), .B(new_n303), .C1(new_n369), .C2(new_n306), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n361), .A2(new_n367), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n367), .B1(new_n361), .B2(new_n370), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT30), .ZN(new_n373));
  NOR3_X1   g172(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n361), .A2(new_n370), .ZN(new_n375));
  NOR3_X1   g174(.A1(new_n375), .A2(KEYINPUT30), .A3(new_n366), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n286), .A2(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(G78gat), .B(G106gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n380), .B(KEYINPUT31), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(G50gat), .ZN(new_n382));
  XOR2_X1   g181(.A(new_n382), .B(KEYINPUT79), .Z(new_n383));
  NAND2_X1  g182(.A1(new_n302), .A2(KEYINPUT80), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT80), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n293), .A2(new_n385), .A3(new_n297), .A4(new_n301), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n384), .A2(new_n296), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n357), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n244), .B1(new_n388), .B2(new_n251), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n303), .B1(new_n357), .B2(new_n256), .ZN(new_n390));
  INV_X1    g189(.A(G228gat), .ZN(new_n391));
  INV_X1    g190(.A(G233gat), .ZN(new_n392));
  OAI22_X1  g191(.A1(new_n389), .A2(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT81), .ZN(new_n394));
  INV_X1    g193(.A(new_n302), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n297), .B1(new_n293), .B2(KEYINPUT22), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n394), .B(new_n357), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n251), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n394), .B1(new_n303), .B2(new_n357), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n243), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n391), .A2(new_n392), .ZN(new_n401));
  INV_X1    g200(.A(new_n390), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(G22gat), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n393), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT82), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n404), .B1(new_n393), .B2(new_n403), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  AOI211_X1 g209(.A(KEYINPUT82), .B(new_n404), .C1(new_n393), .C2(new_n403), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n383), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n409), .A2(new_n382), .A3(new_n405), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(G227gat), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n416), .A2(new_n392), .ZN(new_n417));
  AND4_X1   g216(.A1(new_n227), .A2(new_n333), .A3(new_n349), .A4(new_n355), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n227), .B1(new_n359), .B2(new_n349), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(G15gat), .B(G43gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(G71gat), .ZN(new_n422));
  INV_X1    g221(.A(G99gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT33), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n420), .A2(KEYINPUT32), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT73), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n420), .A2(KEYINPUT73), .A3(KEYINPUT32), .A4(new_n425), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT33), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n420), .B1(KEYINPUT32), .B2(new_n430), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n428), .A2(new_n429), .B1(new_n424), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT74), .ZN(new_n433));
  INV_X1    g232(.A(new_n227), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n356), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n359), .A2(new_n227), .A3(new_n349), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n435), .B(new_n436), .C1(new_n416), .C2(new_n392), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n437), .B(KEYINPUT34), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n432), .A2(new_n433), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n438), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n431), .A2(new_n424), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT32), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n435), .A2(new_n436), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n442), .B1(new_n443), .B2(new_n417), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT73), .B1(new_n444), .B2(new_n425), .ZN(new_n445));
  INV_X1    g244(.A(new_n429), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n441), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n440), .B1(new_n447), .B2(KEYINPUT74), .ZN(new_n448));
  OAI22_X1  g247(.A1(new_n413), .A2(new_n415), .B1(new_n439), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT35), .B1(new_n379), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n377), .B1(new_n284), .B2(new_n285), .ZN(new_n451));
  INV_X1    g250(.A(new_n383), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n408), .B1(new_n406), .B2(new_n405), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n452), .B1(new_n453), .B2(new_n411), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n414), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n432), .A2(new_n440), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n432), .A2(new_n440), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(KEYINPUT85), .B(KEYINPUT35), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n451), .A2(new_n455), .A3(new_n459), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n450), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n413), .A2(new_n415), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT36), .B1(new_n439), .B2(new_n448), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT36), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n465), .B1(new_n457), .B2(new_n458), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n379), .A2(new_n463), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n375), .A2(KEYINPUT37), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT38), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT37), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n361), .A2(new_n370), .A3(new_n470), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n468), .A2(new_n469), .A3(new_n366), .A4(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n468), .A2(new_n366), .A3(new_n471), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n473), .B1(KEYINPUT38), .B2(new_n371), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n284), .A2(new_n285), .A3(new_n472), .A4(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT83), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n247), .A2(new_n250), .A3(new_n258), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT39), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(new_n478), .A3(new_n260), .ZN(new_n479));
  AND2_X1   g278(.A1(new_n479), .A2(new_n279), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n477), .A2(new_n260), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n261), .A2(new_n249), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n248), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n481), .A2(KEYINPUT39), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n476), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT84), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n486), .B1(new_n480), .B2(new_n484), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT40), .ZN(new_n488));
  OAI22_X1  g287(.A1(KEYINPUT84), .A2(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n484), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n479), .A2(new_n279), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT83), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n492), .A2(new_n486), .A3(KEYINPUT40), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n489), .A2(new_n377), .A3(new_n283), .A4(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n475), .A2(new_n494), .A3(new_n455), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n467), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n462), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(G15gat), .B(G22gat), .ZN(new_n498));
  INV_X1    g297(.A(G1gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT16), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n501), .B1(G1gat), .B2(new_n498), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(G8gat), .ZN(new_n503));
  INV_X1    g302(.A(G8gat), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n501), .B(new_n504), .C1(G1gat), .C2(new_n498), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G71gat), .B(G78gat), .ZN(new_n507));
  OR2_X1    g306(.A1(new_n507), .A2(KEYINPUT94), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(KEYINPUT94), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(G57gat), .B(G64gat), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n508), .B(new_n509), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT95), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n510), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n514), .B(new_n507), .C1(new_n513), .C2(new_n511), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n506), .B1(new_n517), .B2(KEYINPUT21), .ZN(new_n518));
  XOR2_X1   g317(.A(new_n518), .B(G183gat), .Z(new_n519));
  NAND2_X1  g318(.A1(G231gat), .A2(G233gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n518), .B(G183gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n522), .A2(G231gat), .A3(G233gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G127gat), .B(G155gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(new_n299), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n517), .A2(KEYINPUT21), .ZN(new_n528));
  XNOR2_X1  g327(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n526), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n532), .B1(new_n521), .B2(new_n523), .ZN(new_n533));
  OR3_X1    g332(.A1(new_n527), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n531), .B1(new_n527), .B2(new_n533), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT96), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT7), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n539), .A2(G85gat), .A3(G92gat), .A4(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(G85gat), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n537), .B(new_n538), .C1(new_n542), .C2(new_n365), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(G99gat), .A2(G106gat), .ZN(new_n545));
  AOI22_X1  g344(.A1(KEYINPUT8), .A2(new_n545), .B1(new_n542), .B2(new_n365), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n546), .A2(KEYINPUT97), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(KEYINPUT97), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n544), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  XOR2_X1   g348(.A(G99gat), .B(G106gat), .Z(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  OR3_X1    g350(.A1(new_n549), .A2(KEYINPUT99), .A3(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT99), .B1(new_n549), .B2(new_n551), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n546), .A2(KEYINPUT97), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n546), .A2(KEYINPUT97), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n541), .B(new_n543), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  NOR3_X1   g356(.A1(new_n557), .A2(KEYINPUT98), .A3(new_n550), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT98), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n559), .B1(new_n549), .B2(new_n551), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n554), .A2(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(KEYINPUT88), .B(G36gat), .Z(new_n563));
  NAND3_X1  g362(.A1(new_n563), .A2(KEYINPUT89), .A3(G29gat), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT89), .ZN(new_n565));
  XNOR2_X1  g364(.A(KEYINPUT88), .B(G36gat), .ZN(new_n566));
  INV_X1    g365(.A(G29gat), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(G43gat), .B(G50gat), .Z(new_n570));
  INV_X1    g369(.A(KEYINPUT15), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g371(.A1(G29gat), .A2(G36gat), .ZN(new_n573));
  XOR2_X1   g372(.A(new_n573), .B(KEYINPUT14), .Z(new_n574));
  NAND3_X1  g373(.A1(new_n569), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n570), .A2(new_n571), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n576), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n569), .A2(new_n578), .A3(new_n572), .A4(new_n574), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n562), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT17), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n577), .A2(KEYINPUT17), .A3(new_n579), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n581), .B(new_n582), .C1(new_n562), .C2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G134gat), .B(G162gat), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G190gat), .B(G218gat), .ZN(new_n591));
  AOI21_X1  g390(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n587), .A2(new_n588), .ZN(new_n594));
  AND3_X1   g393(.A1(new_n590), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n593), .B1(new_n590), .B2(new_n594), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n536), .A2(new_n597), .ZN(new_n598));
  AND3_X1   g397(.A1(new_n503), .A2(new_n505), .A3(KEYINPUT90), .ZN(new_n599));
  AOI21_X1  g398(.A(KEYINPUT90), .B1(new_n503), .B2(new_n505), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n584), .A2(new_n585), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(G229gat), .A2(G233gat), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT91), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n604), .B1(new_n580), .B2(new_n506), .ZN(new_n605));
  AND3_X1   g404(.A1(new_n580), .A2(new_n604), .A3(new_n506), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n602), .B(new_n603), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(KEYINPUT92), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT18), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n606), .A2(new_n605), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n580), .A2(new_n506), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(new_n603), .B(KEYINPUT93), .Z(new_n613));
  XOR2_X1   g412(.A(new_n613), .B(KEYINPUT13), .Z(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT18), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n607), .A2(KEYINPUT92), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n609), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(G113gat), .B(G141gat), .Z(new_n619));
  XNOR2_X1  g418(.A(G169gat), .B(G197gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(KEYINPUT87), .B(KEYINPUT12), .Z(new_n624));
  XOR2_X1   g423(.A(new_n623), .B(new_n624), .Z(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n618), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n609), .A2(new_n615), .A3(new_n625), .A4(new_n617), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G230gat), .A2(G233gat), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  OR2_X1    g430(.A1(new_n557), .A2(KEYINPUT100), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n557), .A2(KEYINPUT100), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n632), .A2(new_n550), .A3(new_n633), .ZN(new_n634));
  OAI211_X1 g433(.A(new_n634), .B(new_n517), .C1(new_n560), .C2(new_n558), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n516), .B1(new_n554), .B2(new_n561), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT10), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n562), .A2(KEYINPUT10), .A3(new_n517), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n631), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n635), .A2(new_n636), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n631), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G176gat), .B(G204gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT101), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(G120gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(new_n237), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n648), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n641), .A2(new_n643), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n598), .A2(new_n629), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n497), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n654), .A2(new_n286), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(new_n499), .ZN(G1324gat));
  NOR2_X1   g455(.A1(new_n654), .A2(new_n378), .ZN(new_n657));
  NAND2_X1  g456(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n658));
  OR2_X1    g457(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n659));
  AND3_X1   g458(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n660), .A2(KEYINPUT42), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(KEYINPUT42), .ZN(new_n662));
  OAI211_X1 g461(.A(new_n661), .B(new_n662), .C1(new_n504), .C2(new_n657), .ZN(G1325gat));
  INV_X1    g462(.A(G15gat), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n464), .A2(new_n466), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n654), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n497), .A2(new_n459), .A3(new_n653), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n666), .B1(new_n664), .B2(new_n667), .ZN(G1326gat));
  NOR2_X1   g467(.A1(new_n654), .A2(new_n455), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT43), .B(G22gat), .Z(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1327gat));
  INV_X1    g470(.A(KEYINPUT104), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT103), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n475), .A2(new_n494), .A3(new_n455), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n438), .B1(new_n432), .B2(new_n433), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n447), .A2(KEYINPUT74), .A3(new_n440), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n465), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n447), .A2(new_n438), .ZN(new_n678));
  AOI21_X1  g477(.A(KEYINPUT36), .B1(new_n678), .B2(new_n456), .ZN(new_n679));
  OAI22_X1  g478(.A1(new_n451), .A2(new_n455), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n673), .B1(new_n674), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n379), .A2(new_n463), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n682), .A2(new_n495), .A3(KEYINPUT103), .A4(new_n665), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n681), .A2(new_n462), .A3(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685));
  INV_X1    g484(.A(new_n597), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  AOI22_X1  g486(.A1(new_n450), .A2(new_n461), .B1(new_n467), .B2(new_n495), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT44), .B1(new_n688), .B2(new_n597), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n536), .A2(new_n629), .A3(new_n652), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT102), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n672), .B1(new_n693), .B2(new_n286), .ZN(new_n694));
  INV_X1    g493(.A(new_n286), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n690), .A2(KEYINPUT104), .A3(new_n695), .A4(new_n692), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n694), .A2(G29gat), .A3(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n497), .A2(new_n686), .A3(new_n691), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n699), .A2(new_n567), .A3(new_n695), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT45), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n697), .A2(new_n701), .ZN(G1328gat));
  NOR3_X1   g501(.A1(new_n698), .A2(new_n378), .A3(new_n563), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT46), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n563), .B1(new_n693), .B2(new_n378), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(G1329gat));
  NOR3_X1   g505(.A1(new_n698), .A2(new_n457), .A3(new_n458), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n707), .A2(G43gat), .ZN(new_n708));
  INV_X1    g507(.A(new_n665), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n690), .A2(G43gat), .A3(new_n709), .A4(new_n692), .ZN(new_n710));
  AOI211_X1 g509(.A(KEYINPUT105), .B(KEYINPUT47), .C1(new_n708), .C2(new_n710), .ZN(new_n711));
  OR2_X1    g510(.A1(KEYINPUT105), .A2(KEYINPUT47), .ZN(new_n712));
  NAND2_X1  g511(.A1(KEYINPUT105), .A2(KEYINPUT47), .ZN(new_n713));
  AND4_X1   g512(.A1(new_n712), .A2(new_n708), .A3(new_n710), .A4(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n711), .A2(new_n714), .ZN(G1330gat));
  NAND2_X1  g514(.A1(new_n699), .A2(KEYINPUT106), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT106), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n698), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n716), .A2(new_n463), .A3(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(G50gat), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n690), .A2(G50gat), .A3(new_n463), .A4(new_n692), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(KEYINPUT48), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT48), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n721), .A2(new_n725), .A3(new_n722), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(G1331gat));
  NAND2_X1  g526(.A1(new_n627), .A2(new_n628), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n598), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n684), .A2(new_n652), .A3(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(new_n286), .ZN(new_n731));
  XOR2_X1   g530(.A(KEYINPUT107), .B(G57gat), .Z(new_n732));
  XNOR2_X1  g531(.A(new_n731), .B(new_n732), .ZN(G1332gat));
  AOI211_X1 g532(.A(new_n378), .B(new_n730), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n734));
  NOR2_X1   g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1333gat));
  XNOR2_X1  g535(.A(new_n459), .B(KEYINPUT108), .ZN(new_n737));
  AND4_X1   g536(.A1(new_n652), .A2(new_n684), .A3(new_n729), .A4(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n709), .A2(G71gat), .ZN(new_n739));
  OAI22_X1  g538(.A1(new_n738), .A2(G71gat), .B1(new_n730), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g540(.A1(new_n730), .A2(new_n455), .ZN(new_n742));
  XOR2_X1   g541(.A(new_n742), .B(G78gat), .Z(G1335gat));
  INV_X1    g542(.A(new_n652), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n536), .A2(new_n728), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  AOI211_X1 g545(.A(new_n744), .B(new_n746), .C1(new_n687), .C2(new_n689), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(G85gat), .B1(new_n748), .B2(new_n286), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n684), .A2(new_n686), .A3(new_n745), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n684), .A2(KEYINPUT51), .A3(new_n686), .A4(new_n745), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT109), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n753), .A2(new_n754), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n752), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n652), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n695), .A2(new_n542), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n749), .B1(new_n758), .B2(new_n759), .ZN(G1336gat));
  NOR2_X1   g559(.A1(new_n378), .A2(G92gat), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(new_n652), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n684), .A2(new_n686), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n763), .A2(KEYINPUT109), .A3(KEYINPUT51), .A4(new_n745), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n753), .A2(new_n754), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n751), .A2(KEYINPUT110), .ZN(new_n767));
  OR2_X1    g566(.A1(new_n751), .A2(KEYINPUT110), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n750), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n762), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n365), .B1(new_n747), .B2(new_n377), .ZN(new_n771));
  OAI21_X1  g570(.A(KEYINPUT52), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n757), .A2(new_n652), .A3(new_n761), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n690), .A2(new_n377), .A3(new_n652), .A4(new_n745), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT52), .B1(new_n774), .B2(G92gat), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n772), .A2(new_n776), .ZN(G1337gat));
  NAND3_X1  g576(.A1(new_n747), .A2(KEYINPUT111), .A3(new_n709), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n690), .A2(new_n709), .A3(new_n652), .A4(new_n745), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT111), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n778), .A2(new_n781), .A3(G99gat), .ZN(new_n782));
  AOI22_X1  g581(.A1(new_n764), .A2(new_n765), .B1(new_n751), .B2(new_n750), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n459), .A2(new_n423), .A3(new_n652), .ZN(new_n784));
  XOR2_X1   g583(.A(new_n784), .B(KEYINPUT112), .Z(new_n785));
  OAI21_X1  g584(.A(new_n782), .B1(new_n783), .B2(new_n785), .ZN(G1338gat));
  NAND4_X1  g585(.A1(new_n690), .A2(new_n463), .A3(new_n652), .A4(new_n745), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(G106gat), .ZN(new_n788));
  XOR2_X1   g587(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n789));
  OR3_X1    g588(.A1(new_n455), .A2(new_n744), .A3(G106gat), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n788), .B(new_n789), .C1(new_n783), .C2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n769), .B1(new_n755), .B2(new_n756), .ZN(new_n792));
  XOR2_X1   g591(.A(new_n790), .B(KEYINPUT113), .Z(new_n793));
  AOI22_X1  g592(.A1(new_n792), .A2(new_n793), .B1(G106gat), .B2(new_n787), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n791), .B1(new_n794), .B2(new_n795), .ZN(G1339gat));
  INV_X1    g595(.A(new_n536), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n638), .A2(new_n631), .A3(new_n639), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT54), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n800), .A2(new_n640), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n638), .A2(new_n639), .ZN(new_n802));
  XNOR2_X1  g601(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n802), .A2(new_n630), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n648), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n798), .B1(new_n801), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n650), .B1(new_n640), .B2(new_n803), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n807), .B(KEYINPUT55), .C1(new_n640), .C2(new_n800), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n728), .A2(new_n651), .A3(new_n806), .A4(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n810), .B1(new_n612), .B2(new_n614), .ZN(new_n811));
  INV_X1    g610(.A(new_n614), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n610), .A2(KEYINPUT116), .A3(new_n611), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n603), .B1(new_n610), .B2(new_n602), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n623), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n652), .A2(new_n816), .A3(new_n628), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n686), .B1(new_n809), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n806), .A2(new_n651), .A3(new_n808), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n816), .A2(new_n628), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n819), .A2(new_n820), .A3(new_n597), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n797), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n729), .A2(new_n744), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR4_X1   g623(.A1(new_n286), .A2(new_n377), .A3(new_n457), .A4(new_n458), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n824), .A2(new_n455), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(KEYINPUT117), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n824), .A2(new_n828), .A3(new_n455), .A4(new_n825), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(G113gat), .B1(new_n830), .B2(new_n629), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n286), .B1(new_n822), .B2(new_n823), .ZN(new_n832));
  INV_X1    g631(.A(new_n449), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n832), .A2(new_n378), .A3(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(G113gat), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n835), .A3(new_n728), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n831), .A2(new_n836), .ZN(G1340gat));
  OAI21_X1  g636(.A(G120gat), .B1(new_n830), .B2(new_n744), .ZN(new_n838));
  INV_X1    g637(.A(G120gat), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n834), .A2(new_n839), .A3(new_n652), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(KEYINPUT118), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT118), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n838), .A2(new_n843), .A3(new_n840), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n844), .ZN(G1341gat));
  NAND2_X1  g644(.A1(new_n209), .A2(new_n211), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n830), .A2(new_n846), .A3(new_n797), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n834), .A2(new_n536), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n847), .B1(new_n846), .B2(new_n848), .ZN(G1342gat));
  OAI211_X1 g648(.A(new_n834), .B(new_n686), .C1(new_n214), .C2(new_n215), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n851));
  OAI21_X1  g650(.A(G134gat), .B1(new_n830), .B2(new_n597), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(G1343gat));
  NAND3_X1  g653(.A1(new_n665), .A2(new_n695), .A3(new_n378), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n455), .B1(new_n822), .B2(new_n823), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT57), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT119), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n819), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n806), .A2(KEYINPUT119), .A3(new_n808), .A4(new_n651), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(new_n728), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n686), .B1(new_n862), .B2(new_n817), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n797), .B1(new_n863), .B2(new_n821), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n455), .B1(new_n864), .B2(new_n823), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n858), .B(new_n728), .C1(new_n865), .C2(new_n857), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(G141gat), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n832), .B(KEYINPUT120), .ZN(new_n868));
  OR3_X1    g667(.A1(new_n709), .A2(KEYINPUT121), .A3(new_n455), .ZN(new_n869));
  OAI21_X1  g668(.A(KEYINPUT121), .B1(new_n709), .B2(new_n455), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n377), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n868), .A2(new_n235), .A3(new_n728), .A4(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n867), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(KEYINPUT58), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT58), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n867), .A2(new_n872), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(new_n876), .ZN(G1344gat));
  INV_X1    g676(.A(KEYINPUT59), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n864), .A2(new_n823), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(new_n857), .A3(new_n463), .ZN(new_n880));
  INV_X1    g679(.A(new_n855), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n856), .A2(new_n857), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n880), .A2(new_n652), .A3(new_n881), .A4(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n878), .B1(new_n883), .B2(G148gat), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n858), .B(new_n652), .C1(new_n865), .C2(new_n857), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n885), .A2(new_n878), .A3(G148gat), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n868), .A2(new_n871), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n652), .A2(new_n237), .ZN(new_n888));
  OAI22_X1  g687(.A1(new_n884), .A2(new_n886), .B1(new_n887), .B2(new_n888), .ZN(G1345gat));
  NOR2_X1   g688(.A1(new_n887), .A2(new_n797), .ZN(new_n890));
  OR2_X1    g689(.A1(new_n865), .A2(new_n857), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n536), .A3(new_n858), .ZN(new_n892));
  MUX2_X1   g691(.A(new_n890), .B(new_n892), .S(G155gat), .Z(G1346gat));
  NOR2_X1   g692(.A1(new_n887), .A2(new_n597), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n891), .A2(new_n686), .A3(new_n858), .ZN(new_n895));
  MUX2_X1   g694(.A(new_n894), .B(new_n895), .S(G162gat), .Z(G1347gat));
  NOR2_X1   g695(.A1(new_n695), .A2(new_n378), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n737), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n817), .B1(new_n819), .B2(new_n629), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n597), .ZN(new_n900));
  OR3_X1    g699(.A1(new_n819), .A2(new_n820), .A3(new_n597), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n536), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n598), .A2(new_n728), .A3(new_n652), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n455), .B(new_n898), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n824), .A2(KEYINPUT122), .A3(new_n455), .A4(new_n898), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n906), .A2(new_n728), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(G169gat), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n824), .A2(new_n833), .A3(new_n897), .ZN(new_n910));
  OR2_X1    g709(.A1(new_n910), .A2(G169gat), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n909), .B1(new_n629), .B2(new_n911), .ZN(G1348gat));
  INV_X1    g711(.A(G176gat), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n913), .B1(new_n910), .B2(new_n744), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n914), .A2(KEYINPUT123), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(KEYINPUT123), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n906), .A2(G176gat), .A3(new_n652), .A4(new_n907), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(G1349gat));
  NAND3_X1  g717(.A1(new_n906), .A2(new_n536), .A3(new_n907), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n311), .A3(new_n312), .ZN(new_n920));
  OR3_X1    g719(.A1(new_n910), .A2(new_n347), .A3(new_n797), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(KEYINPUT60), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT60), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n920), .A2(new_n924), .A3(new_n921), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(G1350gat));
  NAND3_X1  g725(.A1(new_n906), .A2(new_n686), .A3(new_n907), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(G190gat), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n927), .A2(KEYINPUT124), .A3(G190gat), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n930), .A2(KEYINPUT61), .A3(new_n931), .ZN(new_n932));
  OR3_X1    g731(.A1(new_n910), .A2(new_n341), .A3(new_n597), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT61), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n928), .A2(new_n929), .A3(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n932), .A2(new_n933), .A3(new_n935), .ZN(G1351gat));
  AND2_X1   g735(.A1(new_n880), .A2(new_n882), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n897), .A2(new_n665), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT126), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(G197gat), .B1(new_n940), .B2(new_n629), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n856), .A2(new_n938), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(KEYINPUT125), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT125), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n856), .A2(new_n944), .A3(new_n938), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(G197gat), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n946), .A2(new_n947), .A3(new_n728), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n941), .A2(new_n948), .ZN(G1352gat));
  NAND3_X1  g748(.A1(new_n937), .A2(new_n652), .A3(new_n939), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(G204gat), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n942), .A2(G204gat), .A3(new_n744), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT62), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n953), .ZN(G1353gat));
  NAND4_X1  g753(.A1(new_n943), .A2(new_n299), .A3(new_n536), .A4(new_n945), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT127), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n880), .A2(new_n536), .A3(new_n882), .A4(new_n939), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(G211gat), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(KEYINPUT63), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT63), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n957), .A2(new_n960), .A3(G211gat), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n956), .A2(new_n959), .A3(new_n961), .ZN(G1354gat));
  OAI21_X1  g761(.A(G218gat), .B1(new_n940), .B2(new_n597), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n946), .A2(new_n300), .A3(new_n686), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(G1355gat));
endmodule


