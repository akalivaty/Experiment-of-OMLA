

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596;

  XNOR2_X1 U326 ( .A(n476), .B(n475), .ZN(n537) );
  INV_X1 U327 ( .A(KEYINPUT48), .ZN(n473) );
  XNOR2_X1 U328 ( .A(KEYINPUT89), .B(n449), .ZN(n527) );
  INV_X1 U329 ( .A(n348), .ZN(n323) );
  XNOR2_X1 U330 ( .A(n478), .B(KEYINPUT54), .ZN(n479) );
  INV_X1 U331 ( .A(G92GAT), .ZN(n397) );
  XNOR2_X1 U332 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U333 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U334 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U335 ( .A(KEYINPUT55), .B(KEYINPUT117), .ZN(n483) );
  XNOR2_X1 U336 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U337 ( .A(n484), .B(n483), .ZN(n486) );
  NOR2_X1 U338 ( .A1(n525), .A2(n516), .ZN(n522) );
  XOR2_X1 U339 ( .A(n482), .B(KEYINPUT28), .Z(n540) );
  XNOR2_X1 U340 ( .A(n488), .B(G183GAT), .ZN(n489) );
  XNOR2_X1 U341 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U342 ( .A(n490), .B(n489), .ZN(G1350GAT) );
  XNOR2_X1 U343 ( .A(n461), .B(n460), .ZN(G1330GAT) );
  XNOR2_X1 U344 ( .A(G22GAT), .B(G15GAT), .ZN(n294) );
  XNOR2_X1 U345 ( .A(n294), .B(KEYINPUT66), .ZN(n335) );
  XOR2_X1 U346 ( .A(n335), .B(KEYINPUT29), .Z(n296) );
  NAND2_X1 U347 ( .A1(G229GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U348 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U349 ( .A(KEYINPUT65), .B(KEYINPUT30), .Z(n298) );
  XNOR2_X1 U350 ( .A(G197GAT), .B(G1GAT), .ZN(n297) );
  XNOR2_X1 U351 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U352 ( .A(n300), .B(n299), .Z(n302) );
  XOR2_X1 U353 ( .A(G141GAT), .B(G113GAT), .Z(n415) );
  XOR2_X1 U354 ( .A(G169GAT), .B(G8GAT), .Z(n396) );
  XNOR2_X1 U355 ( .A(n415), .B(n396), .ZN(n301) );
  XNOR2_X1 U356 ( .A(n302), .B(n301), .ZN(n307) );
  XNOR2_X1 U357 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n303) );
  XNOR2_X1 U358 ( .A(n303), .B(G29GAT), .ZN(n304) );
  XOR2_X1 U359 ( .A(n304), .B(KEYINPUT8), .Z(n306) );
  XNOR2_X1 U360 ( .A(G43GAT), .B(G50GAT), .ZN(n305) );
  XOR2_X1 U361 ( .A(n306), .B(n305), .Z(n361) );
  XNOR2_X1 U362 ( .A(n307), .B(n361), .ZN(n585) );
  XNOR2_X1 U363 ( .A(n585), .B(KEYINPUT67), .ZN(n565) );
  XOR2_X1 U364 ( .A(KEYINPUT70), .B(KEYINPUT71), .Z(n309) );
  XNOR2_X1 U365 ( .A(G57GAT), .B(KEYINPUT32), .ZN(n308) );
  XOR2_X1 U366 ( .A(n309), .B(n308), .Z(n333) );
  INV_X1 U367 ( .A(KEYINPUT73), .ZN(n310) );
  NAND2_X1 U368 ( .A1(G64GAT), .A2(n310), .ZN(n313) );
  INV_X1 U369 ( .A(G64GAT), .ZN(n311) );
  NAND2_X1 U370 ( .A1(n311), .A2(KEYINPUT73), .ZN(n312) );
  NAND2_X1 U371 ( .A1(n313), .A2(n312), .ZN(n315) );
  XNOR2_X1 U372 ( .A(G176GAT), .B(G204GAT), .ZN(n314) );
  XNOR2_X1 U373 ( .A(n315), .B(n314), .ZN(n389) );
  NAND2_X1 U374 ( .A1(n397), .A2(KEYINPUT72), .ZN(n318) );
  INV_X1 U375 ( .A(KEYINPUT72), .ZN(n316) );
  NAND2_X1 U376 ( .A1(n316), .A2(G92GAT), .ZN(n317) );
  NAND2_X1 U377 ( .A1(n318), .A2(n317), .ZN(n320) );
  XNOR2_X1 U378 ( .A(G99GAT), .B(G85GAT), .ZN(n319) );
  XNOR2_X1 U379 ( .A(n320), .B(n319), .ZN(n351) );
  XNOR2_X1 U380 ( .A(n389), .B(n351), .ZN(n324) );
  XOR2_X1 U381 ( .A(KEYINPUT68), .B(KEYINPUT13), .Z(n322) );
  XNOR2_X1 U382 ( .A(G71GAT), .B(KEYINPUT69), .ZN(n321) );
  XNOR2_X1 U383 ( .A(n322), .B(n321), .ZN(n348) );
  XNOR2_X1 U384 ( .A(n324), .B(n323), .ZN(n329) );
  XNOR2_X1 U385 ( .A(KEYINPUT74), .B(KEYINPUT31), .ZN(n326) );
  AND2_X1 U386 ( .A1(G230GAT), .A2(G233GAT), .ZN(n325) );
  XNOR2_X1 U387 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U388 ( .A(KEYINPUT33), .B(n327), .Z(n328) );
  XNOR2_X1 U389 ( .A(n329), .B(n328), .ZN(n331) );
  XOR2_X1 U390 ( .A(G106GAT), .B(G78GAT), .Z(n368) );
  XOR2_X1 U391 ( .A(G120GAT), .B(G148GAT), .Z(n405) );
  XNOR2_X1 U392 ( .A(n368), .B(n405), .ZN(n330) );
  XNOR2_X1 U393 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U394 ( .A(n333), .B(n332), .ZN(n588) );
  NAND2_X1 U395 ( .A1(n565), .A2(n588), .ZN(n334) );
  XNOR2_X1 U396 ( .A(n334), .B(KEYINPUT75), .ZN(n494) );
  XOR2_X1 U397 ( .A(G183GAT), .B(G211GAT), .Z(n388) );
  XOR2_X1 U398 ( .A(n388), .B(G78GAT), .Z(n337) );
  XNOR2_X1 U399 ( .A(n335), .B(G155GAT), .ZN(n336) );
  XNOR2_X1 U400 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U401 ( .A(KEYINPUT77), .B(KEYINPUT14), .Z(n339) );
  NAND2_X1 U402 ( .A1(G231GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U403 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U404 ( .A(n341), .B(n340), .Z(n346) );
  XOR2_X1 U405 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n343) );
  XNOR2_X1 U406 ( .A(G8GAT), .B(G64GAT), .ZN(n342) );
  XNOR2_X1 U407 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U408 ( .A(n344), .B(KEYINPUT78), .ZN(n345) );
  XNOR2_X1 U409 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U410 ( .A(n348), .B(n347), .ZN(n350) );
  XNOR2_X1 U411 ( .A(G1GAT), .B(G127GAT), .ZN(n349) );
  XOR2_X1 U412 ( .A(n349), .B(G57GAT), .Z(n403) );
  XOR2_X1 U413 ( .A(n350), .B(n403), .Z(n465) );
  XOR2_X1 U414 ( .A(n351), .B(G134GAT), .Z(n353) );
  NAND2_X1 U415 ( .A1(G232GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U416 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U417 ( .A(KEYINPUT10), .B(G106GAT), .Z(n355) );
  XNOR2_X1 U418 ( .A(G190GAT), .B(G162GAT), .ZN(n354) );
  XNOR2_X1 U419 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U420 ( .A(n357), .B(n356), .Z(n363) );
  XOR2_X1 U421 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n359) );
  XNOR2_X1 U422 ( .A(G218GAT), .B(KEYINPUT76), .ZN(n358) );
  XNOR2_X1 U423 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U424 ( .A(n361), .B(n360), .Z(n362) );
  XOR2_X1 U425 ( .A(n363), .B(n362), .Z(n563) );
  XNOR2_X1 U426 ( .A(n563), .B(KEYINPUT102), .ZN(n364) );
  XNOR2_X1 U427 ( .A(KEYINPUT36), .B(n364), .ZN(n592) );
  XOR2_X1 U428 ( .A(KEYINPUT24), .B(KEYINPUT84), .Z(n366) );
  XNOR2_X1 U429 ( .A(G50GAT), .B(G204GAT), .ZN(n365) );
  XNOR2_X1 U430 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U431 ( .A(n368), .B(n367), .Z(n370) );
  NAND2_X1 U432 ( .A1(G228GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U433 ( .A(n370), .B(n369), .ZN(n384) );
  XOR2_X1 U434 ( .A(KEYINPUT83), .B(KEYINPUT86), .Z(n372) );
  XNOR2_X1 U435 ( .A(G22GAT), .B(KEYINPUT23), .ZN(n371) );
  XNOR2_X1 U436 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U437 ( .A(G148GAT), .B(G211GAT), .Z(n374) );
  XNOR2_X1 U438 ( .A(G141GAT), .B(KEYINPUT22), .ZN(n373) );
  XNOR2_X1 U439 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U440 ( .A(n376), .B(n375), .Z(n382) );
  XOR2_X1 U441 ( .A(G155GAT), .B(KEYINPUT2), .Z(n378) );
  XNOR2_X1 U442 ( .A(G162GAT), .B(KEYINPUT3), .ZN(n377) );
  XNOR2_X1 U443 ( .A(n378), .B(n377), .ZN(n404) );
  XOR2_X1 U444 ( .A(KEYINPUT21), .B(KEYINPUT85), .Z(n380) );
  XNOR2_X1 U445 ( .A(G197GAT), .B(G218GAT), .ZN(n379) );
  XNOR2_X1 U446 ( .A(n380), .B(n379), .ZN(n393) );
  XNOR2_X1 U447 ( .A(n404), .B(n393), .ZN(n381) );
  XNOR2_X1 U448 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U449 ( .A(n384), .B(n383), .Z(n482) );
  XOR2_X1 U450 ( .A(KEYINPUT17), .B(G190GAT), .Z(n386) );
  XNOR2_X1 U451 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n385) );
  XNOR2_X1 U452 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U453 ( .A(KEYINPUT80), .B(n387), .Z(n437) );
  INV_X1 U454 ( .A(n437), .ZN(n402) );
  XOR2_X1 U455 ( .A(n389), .B(n388), .Z(n391) );
  NAND2_X1 U456 ( .A1(G226GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U457 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U458 ( .A(n392), .B(KEYINPUT91), .Z(n395) );
  XNOR2_X1 U459 ( .A(n393), .B(KEYINPUT90), .ZN(n394) );
  XNOR2_X1 U460 ( .A(n395), .B(n394), .ZN(n400) );
  XNOR2_X1 U461 ( .A(G36GAT), .B(n396), .ZN(n398) );
  XOR2_X1 U462 ( .A(n402), .B(n401), .Z(n442) );
  XNOR2_X1 U463 ( .A(KEYINPUT27), .B(n442), .ZN(n441) );
  XOR2_X1 U464 ( .A(n404), .B(n403), .Z(n419) );
  XOR2_X1 U465 ( .A(G134GAT), .B(KEYINPUT0), .Z(n428) );
  XOR2_X1 U466 ( .A(n428), .B(n405), .Z(n407) );
  NAND2_X1 U467 ( .A1(G225GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U468 ( .A(n407), .B(n406), .ZN(n411) );
  XOR2_X1 U469 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n409) );
  XNOR2_X1 U470 ( .A(KEYINPUT6), .B(KEYINPUT87), .ZN(n408) );
  XNOR2_X1 U471 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U472 ( .A(n411), .B(n410), .Z(n417) );
  XOR2_X1 U473 ( .A(KEYINPUT1), .B(KEYINPUT88), .Z(n413) );
  XNOR2_X1 U474 ( .A(G29GAT), .B(G85GAT), .ZN(n412) );
  XNOR2_X1 U475 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U476 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U477 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U478 ( .A(n419), .B(n418), .ZN(n449) );
  NAND2_X1 U479 ( .A1(n441), .A2(n527), .ZN(n536) );
  NOR2_X1 U480 ( .A1(n540), .A2(n536), .ZN(n438) );
  XOR2_X1 U481 ( .A(G120GAT), .B(G127GAT), .Z(n421) );
  XNOR2_X1 U482 ( .A(G113GAT), .B(KEYINPUT81), .ZN(n420) );
  XNOR2_X1 U483 ( .A(n421), .B(n420), .ZN(n435) );
  XOR2_X1 U484 ( .A(KEYINPUT79), .B(G183GAT), .Z(n423) );
  XNOR2_X1 U485 ( .A(G43GAT), .B(G99GAT), .ZN(n422) );
  XNOR2_X1 U486 ( .A(n423), .B(n422), .ZN(n427) );
  XOR2_X1 U487 ( .A(KEYINPUT82), .B(G176GAT), .Z(n425) );
  XNOR2_X1 U488 ( .A(G169GAT), .B(KEYINPUT20), .ZN(n424) );
  XNOR2_X1 U489 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U490 ( .A(n427), .B(n426), .Z(n433) );
  XOR2_X1 U491 ( .A(G71GAT), .B(n428), .Z(n430) );
  NAND2_X1 U492 ( .A1(G227GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U493 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U494 ( .A(G15GAT), .B(n431), .ZN(n432) );
  XNOR2_X1 U495 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U496 ( .A(n435), .B(n434), .Z(n436) );
  XOR2_X1 U497 ( .A(n437), .B(n436), .Z(n485) );
  NAND2_X1 U498 ( .A1(n438), .A2(n485), .ZN(n452) );
  INV_X1 U499 ( .A(n485), .ZN(n538) );
  NOR2_X1 U500 ( .A1(n482), .A2(n538), .ZN(n440) );
  XNOR2_X1 U501 ( .A(KEYINPUT26), .B(KEYINPUT92), .ZN(n439) );
  XNOR2_X1 U502 ( .A(n440), .B(n439), .ZN(n582) );
  NAND2_X1 U503 ( .A1(n441), .A2(n582), .ZN(n448) );
  XOR2_X1 U504 ( .A(KEYINPUT25), .B(KEYINPUT94), .Z(n446) );
  NAND2_X1 U505 ( .A1(n538), .A2(n442), .ZN(n443) );
  XOR2_X1 U506 ( .A(KEYINPUT93), .B(n443), .Z(n444) );
  NAND2_X1 U507 ( .A1(n444), .A2(n482), .ZN(n445) );
  XNOR2_X1 U508 ( .A(n446), .B(n445), .ZN(n447) );
  NAND2_X1 U509 ( .A1(n448), .A2(n447), .ZN(n450) );
  NAND2_X1 U510 ( .A1(n450), .A2(n449), .ZN(n451) );
  NAND2_X1 U511 ( .A1(n452), .A2(n451), .ZN(n453) );
  XNOR2_X1 U512 ( .A(KEYINPUT95), .B(n453), .ZN(n493) );
  NOR2_X1 U513 ( .A1(n592), .A2(n493), .ZN(n454) );
  NAND2_X1 U514 ( .A1(n465), .A2(n454), .ZN(n455) );
  XOR2_X1 U515 ( .A(KEYINPUT37), .B(n455), .Z(n526) );
  INV_X1 U516 ( .A(n526), .ZN(n456) );
  NAND2_X1 U517 ( .A1(n494), .A2(n456), .ZN(n457) );
  XOR2_X1 U518 ( .A(KEYINPUT38), .B(n457), .Z(n512) );
  NAND2_X1 U519 ( .A1(n512), .A2(n538), .ZN(n461) );
  XOR2_X1 U520 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n459) );
  INV_X1 U521 ( .A(G43GAT), .ZN(n458) );
  XOR2_X1 U522 ( .A(KEYINPUT41), .B(n588), .Z(n558) );
  OR2_X1 U523 ( .A1(n558), .A2(n585), .ZN(n463) );
  INV_X1 U524 ( .A(KEYINPUT46), .ZN(n462) );
  XNOR2_X1 U525 ( .A(n463), .B(n462), .ZN(n464) );
  INV_X1 U526 ( .A(n563), .ZN(n575) );
  NOR2_X1 U527 ( .A1(n464), .A2(n575), .ZN(n466) );
  XOR2_X1 U528 ( .A(KEYINPUT109), .B(n465), .Z(n546) );
  NAND2_X1 U529 ( .A1(n466), .A2(n546), .ZN(n467) );
  XNOR2_X1 U530 ( .A(n467), .B(KEYINPUT47), .ZN(n472) );
  NOR2_X1 U531 ( .A1(n465), .A2(n592), .ZN(n468) );
  XNOR2_X1 U532 ( .A(KEYINPUT45), .B(n468), .ZN(n469) );
  NAND2_X1 U533 ( .A1(n469), .A2(n588), .ZN(n470) );
  NOR2_X1 U534 ( .A1(n565), .A2(n470), .ZN(n471) );
  NOR2_X1 U535 ( .A1(n472), .A2(n471), .ZN(n476) );
  XOR2_X1 U536 ( .A(KEYINPUT64), .B(KEYINPUT110), .Z(n474) );
  INV_X1 U537 ( .A(n537), .ZN(n477) );
  NAND2_X1 U538 ( .A1(n477), .A2(n442), .ZN(n480) );
  XOR2_X1 U539 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n478) );
  NOR2_X1 U540 ( .A1(n527), .A2(n481), .ZN(n583) );
  NAND2_X1 U541 ( .A1(n583), .A2(n482), .ZN(n484) );
  NOR2_X1 U542 ( .A1(n486), .A2(n485), .ZN(n576) );
  INV_X1 U543 ( .A(n576), .ZN(n487) );
  NOR2_X1 U544 ( .A1(n487), .A2(n546), .ZN(n490) );
  XNOR2_X1 U545 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n488) );
  NOR2_X1 U546 ( .A1(n575), .A2(n465), .ZN(n491) );
  XOR2_X1 U547 ( .A(KEYINPUT16), .B(n491), .Z(n492) );
  NOR2_X1 U548 ( .A1(n493), .A2(n492), .ZN(n515) );
  AND2_X1 U549 ( .A1(n494), .A2(n515), .ZN(n505) );
  NAND2_X1 U550 ( .A1(n527), .A2(n505), .ZN(n498) );
  XOR2_X1 U551 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n496) );
  XNOR2_X1 U552 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n495) );
  XNOR2_X1 U553 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U554 ( .A(n498), .B(n497), .ZN(G1324GAT) );
  NAND2_X1 U555 ( .A1(n442), .A2(n505), .ZN(n499) );
  XNOR2_X1 U556 ( .A(n499), .B(KEYINPUT98), .ZN(n500) );
  XNOR2_X1 U557 ( .A(G8GAT), .B(n500), .ZN(G1325GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT100), .B(KEYINPUT35), .Z(n502) );
  NAND2_X1 U559 ( .A1(n505), .A2(n538), .ZN(n501) );
  XNOR2_X1 U560 ( .A(n502), .B(n501), .ZN(n504) );
  XOR2_X1 U561 ( .A(G15GAT), .B(KEYINPUT99), .Z(n503) );
  XNOR2_X1 U562 ( .A(n504), .B(n503), .ZN(G1326GAT) );
  XOR2_X1 U563 ( .A(G22GAT), .B(KEYINPUT101), .Z(n507) );
  NAND2_X1 U564 ( .A1(n505), .A2(n540), .ZN(n506) );
  XNOR2_X1 U565 ( .A(n507), .B(n506), .ZN(G1327GAT) );
  XOR2_X1 U566 ( .A(G29GAT), .B(KEYINPUT39), .Z(n509) );
  NAND2_X1 U567 ( .A1(n512), .A2(n527), .ZN(n508) );
  XNOR2_X1 U568 ( .A(n509), .B(n508), .ZN(G1328GAT) );
  XOR2_X1 U569 ( .A(G36GAT), .B(KEYINPUT103), .Z(n511) );
  NAND2_X1 U570 ( .A1(n512), .A2(n442), .ZN(n510) );
  XNOR2_X1 U571 ( .A(n511), .B(n510), .ZN(G1329GAT) );
  XOR2_X1 U572 ( .A(G50GAT), .B(KEYINPUT105), .Z(n514) );
  NAND2_X1 U573 ( .A1(n540), .A2(n512), .ZN(n513) );
  XNOR2_X1 U574 ( .A(n514), .B(n513), .ZN(G1331GAT) );
  INV_X1 U575 ( .A(n558), .ZN(n570) );
  NAND2_X1 U576 ( .A1(n585), .A2(n570), .ZN(n525) );
  INV_X1 U577 ( .A(n515), .ZN(n516) );
  NAND2_X1 U578 ( .A1(n527), .A2(n522), .ZN(n519) );
  XNOR2_X1 U579 ( .A(G57GAT), .B(KEYINPUT106), .ZN(n517) );
  XNOR2_X1 U580 ( .A(n517), .B(KEYINPUT42), .ZN(n518) );
  XNOR2_X1 U581 ( .A(n519), .B(n518), .ZN(G1332GAT) );
  NAND2_X1 U582 ( .A1(n442), .A2(n522), .ZN(n520) );
  XNOR2_X1 U583 ( .A(n520), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U584 ( .A1(n538), .A2(n522), .ZN(n521) );
  XNOR2_X1 U585 ( .A(n521), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U586 ( .A(G78GAT), .B(KEYINPUT43), .Z(n524) );
  NAND2_X1 U587 ( .A1(n522), .A2(n540), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n524), .B(n523), .ZN(G1335GAT) );
  NOR2_X1 U589 ( .A1(n526), .A2(n525), .ZN(n533) );
  NAND2_X1 U590 ( .A1(n533), .A2(n527), .ZN(n528) );
  XNOR2_X1 U591 ( .A(G85GAT), .B(n528), .ZN(G1336GAT) );
  XOR2_X1 U592 ( .A(G92GAT), .B(KEYINPUT107), .Z(n530) );
  NAND2_X1 U593 ( .A1(n533), .A2(n442), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n530), .B(n529), .ZN(G1337GAT) );
  NAND2_X1 U595 ( .A1(n538), .A2(n533), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n531), .B(KEYINPUT108), .ZN(n532) );
  XNOR2_X1 U597 ( .A(G99GAT), .B(n532), .ZN(G1338GAT) );
  NAND2_X1 U598 ( .A1(n533), .A2(n540), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n534), .B(KEYINPUT44), .ZN(n535) );
  XNOR2_X1 U600 ( .A(G106GAT), .B(n535), .ZN(G1339GAT) );
  NOR2_X1 U601 ( .A1(n537), .A2(n536), .ZN(n554) );
  NAND2_X1 U602 ( .A1(n554), .A2(n538), .ZN(n539) );
  NOR2_X1 U603 ( .A1(n540), .A2(n539), .ZN(n550) );
  NAND2_X1 U604 ( .A1(n550), .A2(n565), .ZN(n541) );
  XNOR2_X1 U605 ( .A(G113GAT), .B(n541), .ZN(G1340GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT111), .B(KEYINPUT49), .Z(n543) );
  NAND2_X1 U607 ( .A1(n550), .A2(n570), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U609 ( .A(G120GAT), .B(n544), .Z(G1341GAT) );
  INV_X1 U610 ( .A(n550), .ZN(n545) );
  NOR2_X1 U611 ( .A1(n546), .A2(n545), .ZN(n548) );
  XNOR2_X1 U612 ( .A(KEYINPUT112), .B(KEYINPUT50), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(n549) );
  XOR2_X1 U614 ( .A(G127GAT), .B(n549), .Z(G1342GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT113), .B(KEYINPUT51), .Z(n552) );
  NAND2_X1 U616 ( .A1(n550), .A2(n575), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U618 ( .A(G134GAT), .B(n553), .Z(G1343GAT) );
  NAND2_X1 U619 ( .A1(n582), .A2(n554), .ZN(n562) );
  NOR2_X1 U620 ( .A1(n585), .A2(n562), .ZN(n555) );
  XOR2_X1 U621 ( .A(G141GAT), .B(n555), .Z(G1344GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT52), .B(KEYINPUT53), .Z(n557) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(KEYINPUT114), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n560) );
  NOR2_X1 U625 ( .A1(n558), .A2(n562), .ZN(n559) );
  XOR2_X1 U626 ( .A(n560), .B(n559), .Z(G1345GAT) );
  NOR2_X1 U627 ( .A1(n465), .A2(n562), .ZN(n561) );
  XOR2_X1 U628 ( .A(G155GAT), .B(n561), .Z(G1346GAT) );
  NOR2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U630 ( .A(G162GAT), .B(n564), .Z(G1347GAT) );
  NAND2_X1 U631 ( .A1(n565), .A2(n576), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT57), .B(KEYINPUT119), .Z(n568) );
  XNOR2_X1 U634 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n569) );
  XOR2_X1 U636 ( .A(KEYINPUT118), .B(n569), .Z(n572) );
  NAND2_X1 U637 ( .A1(n576), .A2(n570), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(G1349GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n574) );
  XNOR2_X1 U640 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n573) );
  XNOR2_X1 U641 ( .A(n574), .B(n573), .ZN(n579) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n577), .B(KEYINPUT122), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1351GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n581) );
  XNOR2_X1 U646 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n587) );
  NAND2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U649 ( .A(KEYINPUT125), .B(n584), .Z(n593) );
  NOR2_X1 U650 ( .A1(n585), .A2(n593), .ZN(n586) );
  XOR2_X1 U651 ( .A(n587), .B(n586), .Z(G1352GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n593), .ZN(n590) );
  XNOR2_X1 U653 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n590), .B(n589), .ZN(G1353GAT) );
  NOR2_X1 U655 ( .A1(n593), .A2(n465), .ZN(n591) );
  XOR2_X1 U656 ( .A(G211GAT), .B(n591), .Z(G1354GAT) );
  NOR2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n595) );
  XNOR2_X1 U658 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n594) );
  XNOR2_X1 U659 ( .A(n595), .B(n594), .ZN(n596) );
  XNOR2_X1 U660 ( .A(G218GAT), .B(n596), .ZN(G1355GAT) );
endmodule

