//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 0 0 1 1 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1267, new_n1268, new_n1269, new_n1271, new_n1272, new_n1273,
    new_n1274, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(G13), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  OAI21_X1  g0013(.A(G50), .B1(G58), .B2(G68), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n207), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(KEYINPUT64), .B(G77), .ZN(new_n219));
  AND2_X1   g0019(.A1(new_n219), .A2(G244), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G58), .A2(G232), .ZN(new_n224));
  NAND4_X1  g0024(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  OAI22_X1  g0025(.A1(new_n220), .A2(new_n225), .B1(new_n206), .B2(new_n207), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n213), .B(new_n218), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G250), .B(G257), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G264), .B(G270), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT65), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n232), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XOR2_X1   g0038(.A(G107), .B(G116), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  NAND3_X1  g0044(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT12), .ZN(new_n249));
  NOR2_X1   g0049(.A1(G20), .A2(G33), .ZN(new_n250));
  AOI22_X1  g0050(.A1(new_n250), .A2(G50), .B1(G20), .B2(new_n247), .ZN(new_n251));
  INV_X1    g0051(.A(G77), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n207), .A2(G33), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n216), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n254), .A2(KEYINPUT11), .A3(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n246), .A2(new_n256), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n206), .A2(G20), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(G68), .A3(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n249), .A2(new_n257), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(KEYINPUT11), .B1(new_n254), .B2(new_n256), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT74), .ZN(new_n265));
  INV_X1    g0065(.A(G1698), .ZN(new_n266));
  AND2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  OAI211_X1 g0068(.A(G226), .B(new_n266), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT69), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT3), .B(G33), .ZN(new_n272));
  NAND4_X1  g0072(.A1(new_n272), .A2(KEYINPUT69), .A3(G226), .A4(new_n266), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G97), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n272), .A2(G232), .A3(G1698), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n271), .A2(new_n273), .A3(new_n274), .A4(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(G1), .A3(G13), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT13), .ZN(new_n281));
  INV_X1    g0081(.A(G41), .ZN(new_n282));
  INV_X1    g0082(.A(G45), .ZN(new_n283));
  AOI21_X1  g0083(.A(G1), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n284), .A2(new_n278), .A3(G274), .ZN(new_n285));
  INV_X1    g0085(.A(G238), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n278), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n285), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n280), .A2(new_n281), .A3(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT71), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n280), .A2(new_n290), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT13), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n280), .A2(KEYINPUT71), .A3(new_n281), .A4(new_n290), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n293), .A2(new_n295), .A3(G179), .A4(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT14), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n281), .B1(new_n280), .B2(new_n290), .ZN(new_n299));
  AOI211_X1 g0099(.A(KEYINPUT13), .B(new_n289), .C1(new_n276), .C2(new_n279), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n298), .B(G169), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G169), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n303), .B1(new_n295), .B2(new_n291), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT73), .B1(new_n304), .B2(new_n298), .ZN(new_n305));
  OAI21_X1  g0105(.A(G169), .B1(new_n299), .B2(new_n300), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT73), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n306), .A2(new_n307), .A3(KEYINPUT14), .ZN(new_n308));
  AOI211_X1 g0108(.A(new_n265), .B(new_n302), .C1(new_n305), .C2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n305), .A2(new_n308), .ZN(new_n310));
  INV_X1    g0110(.A(new_n302), .ZN(new_n311));
  AOI21_X1  g0111(.A(KEYINPUT74), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n264), .B1(new_n309), .B2(new_n312), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n293), .A2(new_n295), .A3(G190), .A4(new_n296), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n314), .A2(new_n263), .ZN(new_n315));
  OAI21_X1  g0115(.A(G200), .B1(new_n299), .B2(new_n300), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT70), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI211_X1 g0118(.A(KEYINPUT70), .B(G200), .C1(new_n299), .C2(new_n300), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT72), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n315), .A2(KEYINPUT72), .A3(new_n320), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n313), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT9), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n255), .A2(new_n216), .ZN(new_n328));
  XOR2_X1   g0128(.A(KEYINPUT8), .B(G58), .Z(new_n329));
  INV_X1    g0129(.A(new_n253), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n329), .A2(new_n330), .B1(G150), .B2(new_n250), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n203), .A2(G20), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n328), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n245), .A2(new_n216), .A3(new_n255), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n259), .A2(G50), .ZN(new_n335));
  OAI22_X1  g0135(.A1(new_n334), .A2(new_n335), .B1(G50), .B2(new_n245), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT67), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n337), .A2(new_n338), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n327), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n272), .A2(G222), .A3(new_n266), .ZN(new_n343));
  INV_X1    g0143(.A(new_n219), .ZN(new_n344));
  INV_X1    g0144(.A(G223), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n272), .A2(G1698), .ZN(new_n346));
  OAI221_X1 g0146(.A(new_n343), .B1(new_n344), .B2(new_n272), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n279), .ZN(new_n348));
  INV_X1    g0148(.A(new_n285), .ZN(new_n349));
  INV_X1    g0149(.A(new_n288), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n349), .B1(G226), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT66), .B(G200), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  OR2_X1    g0155(.A1(new_n333), .A2(new_n336), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT67), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n357), .A2(KEYINPUT9), .A3(new_n339), .ZN(new_n358));
  INV_X1    g0158(.A(new_n352), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G190), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n342), .A2(new_n355), .A3(new_n358), .A4(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT68), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n342), .A2(new_n362), .A3(new_n358), .A4(new_n360), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT10), .ZN(new_n364));
  AND3_X1   g0164(.A1(new_n361), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n361), .B1(new_n364), .B2(new_n363), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n356), .B1(new_n359), .B2(G169), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n352), .A2(G179), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  XNOR2_X1  g0171(.A(KEYINPUT8), .B(G58), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n372), .B1(new_n206), .B2(G20), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n373), .A2(new_n258), .B1(new_n246), .B2(new_n372), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT75), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n374), .B(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT16), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT7), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(new_n272), .B2(G20), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n267), .A2(new_n268), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n380), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n247), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G58), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(new_n247), .ZN(new_n384));
  OAI21_X1  g0184(.A(G20), .B1(new_n384), .B2(new_n201), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n250), .A2(G159), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n377), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(KEYINPUT7), .B1(new_n380), .B2(new_n207), .ZN(new_n389));
  NOR4_X1   g0189(.A1(new_n267), .A2(new_n268), .A3(new_n378), .A4(G20), .ZN(new_n390));
  OAI21_X1  g0190(.A(G68), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n387), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n391), .A2(KEYINPUT16), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n388), .A2(new_n393), .A3(new_n256), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n376), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n345), .A2(new_n266), .ZN(new_n396));
  OAI221_X1 g0196(.A(new_n396), .B1(G226), .B2(new_n266), .C1(new_n267), .C2(new_n268), .ZN(new_n397));
  NAND2_X1  g0197(.A1(G33), .A2(G87), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n279), .ZN(new_n400));
  INV_X1    g0200(.A(G232), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n285), .B1(new_n401), .B2(new_n288), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n400), .A2(G179), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n278), .B1(new_n397), .B2(new_n398), .ZN(new_n405));
  OAI21_X1  g0205(.A(G169), .B1(new_n405), .B2(new_n402), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n395), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT18), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n376), .A2(new_n394), .B1(new_n406), .B2(new_n404), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT18), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(G200), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n414), .B1(new_n400), .B2(new_n403), .ZN(new_n415));
  INV_X1    g0215(.A(G190), .ZN(new_n416));
  NOR3_X1   g0216(.A1(new_n405), .A2(new_n402), .A3(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n418), .A2(new_n376), .A3(new_n394), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT17), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n418), .A2(new_n376), .A3(KEYINPUT17), .A4(new_n394), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n413), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g0224(.A(KEYINPUT15), .B(G87), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n426), .A2(new_n330), .B1(new_n219), .B2(G20), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n329), .A2(new_n250), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n256), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n259), .A2(G77), .ZN(new_n431));
  OAI221_X1 g0231(.A(new_n430), .B1(new_n219), .B2(new_n245), .C1(new_n334), .C2(new_n431), .ZN(new_n432));
  AND2_X1   g0232(.A1(new_n350), .A2(G244), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n272), .A2(G232), .A3(new_n266), .ZN(new_n434));
  INV_X1    g0234(.A(G107), .ZN(new_n435));
  OAI221_X1 g0235(.A(new_n434), .B1(new_n435), .B2(new_n272), .C1(new_n346), .C2(new_n286), .ZN(new_n436));
  AOI211_X1 g0236(.A(new_n349), .B(new_n433), .C1(new_n436), .C2(new_n279), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n432), .B1(new_n437), .B2(G190), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n438), .B1(new_n353), .B2(new_n437), .ZN(new_n439));
  INV_X1    g0239(.A(G179), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n441), .B(new_n432), .C1(G169), .C2(new_n437), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n367), .A2(new_n371), .A3(new_n424), .A4(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n326), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n206), .A2(G33), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n328), .A2(new_n245), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT25), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(new_n245), .B2(G107), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n246), .A2(KEYINPUT25), .A3(new_n435), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n448), .A2(G107), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n207), .B(G87), .C1(new_n267), .C2(new_n268), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT22), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT22), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n272), .A2(new_n456), .A3(new_n207), .A4(G87), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT23), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n459), .A2(new_n435), .A3(G20), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT81), .ZN(new_n461));
  NAND2_X1  g0261(.A1(KEYINPUT23), .A2(G107), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n464));
  OAI22_X1  g0264(.A1(new_n460), .A2(KEYINPUT81), .B1(new_n464), .B2(G20), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n458), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT24), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT24), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n458), .A2(new_n466), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n453), .B1(new_n471), .B2(new_n256), .ZN(new_n472));
  OAI211_X1 g0272(.A(G257), .B(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT82), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n272), .A2(KEYINPUT82), .A3(G257), .A4(G1698), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n272), .A2(G250), .A3(new_n266), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G294), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n475), .A2(new_n476), .A3(new_n477), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n279), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT83), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n479), .A2(KEYINPUT83), .A3(new_n279), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n206), .A2(G45), .ZN(new_n484));
  OR2_X1    g0284(.A1(KEYINPUT5), .A2(G41), .ZN(new_n485));
  NAND2_X1  g0285(.A1(KEYINPUT5), .A2(G41), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n487), .A2(new_n279), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G264), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n485), .A2(new_n486), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n283), .A2(G1), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n490), .A2(G274), .A3(new_n278), .A4(new_n491), .ZN(new_n492));
  AND2_X1   g0292(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n482), .A2(new_n483), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G169), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n479), .A2(new_n279), .B1(G264), .B2(new_n488), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n496), .A2(G179), .A3(new_n492), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n472), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n458), .A2(new_n466), .A3(new_n469), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n469), .B1(new_n458), .B2(new_n466), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n256), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n452), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n482), .A2(new_n416), .A3(new_n483), .A4(new_n493), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n480), .A2(new_n492), .A3(new_n489), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n414), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n502), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n498), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n278), .A2(G274), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n488), .A2(G270), .B1(new_n508), .B2(new_n487), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n272), .A2(G257), .A3(new_n266), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n380), .A2(G303), .ZN(new_n511));
  OAI211_X1 g0311(.A(G264), .B(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n279), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n509), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n448), .A2(G116), .ZN(new_n516));
  INV_X1    g0316(.A(G116), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n246), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G283), .ZN(new_n519));
  INV_X1    g0319(.A(G97), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n519), .B(new_n207), .C1(G33), .C2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n517), .A2(G20), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(new_n256), .A3(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT20), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n523), .A2(new_n524), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n516), .B(new_n518), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT79), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n515), .A2(new_n528), .A3(new_n529), .A4(G179), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n509), .A2(new_n514), .A3(G179), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n518), .B1(new_n447), .B2(new_n517), .ZN(new_n532));
  INV_X1    g0332(.A(new_n527), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n532), .B1(new_n533), .B2(new_n525), .ZN(new_n534));
  OAI21_X1  g0334(.A(KEYINPUT79), .B1(new_n531), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n509), .A2(new_n514), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n528), .A2(new_n537), .A3(G169), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT21), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n538), .A2(KEYINPUT80), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(KEYINPUT80), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n528), .A2(new_n537), .A3(G169), .A4(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n537), .A2(G200), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n543), .B(new_n534), .C1(new_n416), .C2(new_n537), .ZN(new_n544));
  AND4_X1   g0344(.A1(new_n536), .A2(new_n540), .A3(new_n542), .A4(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT19), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n207), .B1(new_n274), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(G97), .A2(G107), .ZN(new_n548));
  INV_X1    g0348(.A(G87), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n207), .B(G68), .C1(new_n267), .C2(new_n268), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n546), .B1(new_n253), .B2(new_n520), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT78), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n551), .A2(new_n552), .A3(KEYINPUT78), .A4(new_n553), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n556), .A2(new_n256), .A3(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n426), .A2(new_n245), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n448), .A2(G87), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n558), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n278), .A2(G274), .A3(new_n491), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n278), .A2(G250), .A3(new_n484), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(G244), .B(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n566));
  OAI211_X1 g0366(.A(G238), .B(new_n266), .C1(new_n267), .C2(new_n268), .ZN(new_n567));
  NAND2_X1  g0367(.A1(G33), .A2(G116), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n565), .B1(new_n279), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n570), .A2(new_n353), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n279), .ZN(new_n572));
  INV_X1    g0372(.A(new_n565), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n572), .A2(G190), .A3(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n572), .A2(new_n440), .A3(new_n573), .ZN(new_n576));
  AOI21_X1  g0376(.A(G169), .B1(new_n572), .B2(new_n573), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n448), .A2(new_n426), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n558), .A2(new_n579), .A3(new_n560), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n562), .A2(new_n575), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(G244), .B(new_n266), .C1(new_n267), .C2(new_n268), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT4), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n272), .A2(KEYINPUT4), .A3(G244), .A4(new_n266), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n272), .A2(G250), .A3(G1698), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n584), .A2(new_n585), .A3(new_n519), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n279), .ZN(new_n588));
  INV_X1    g0388(.A(new_n486), .ZN(new_n589));
  NOR2_X1   g0389(.A1(KEYINPUT5), .A2(G41), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n491), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n591), .A2(G257), .A3(new_n278), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n492), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n588), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n595), .A2(KEYINPUT77), .A3(G200), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n245), .A2(G97), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n597), .B1(new_n448), .B2(G97), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT76), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT6), .ZN(new_n601));
  AND2_X1   g0401(.A1(G97), .A2(G107), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n601), .B1(new_n602), .B2(new_n548), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n435), .A2(KEYINPUT6), .A3(G97), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n207), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n250), .A2(G77), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n600), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n435), .A2(KEYINPUT6), .A3(G97), .ZN(new_n609));
  XNOR2_X1  g0409(.A(G97), .B(G107), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n609), .B1(new_n610), .B2(new_n601), .ZN(new_n611));
  OAI211_X1 g0411(.A(KEYINPUT76), .B(new_n606), .C1(new_n611), .C2(new_n207), .ZN(new_n612));
  OAI21_X1  g0412(.A(G107), .B1(new_n389), .B2(new_n390), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n608), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n599), .B1(new_n614), .B2(new_n256), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT77), .ZN(new_n616));
  AOI21_X1  g0416(.A(G190), .B1(new_n616), .B2(G200), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n596), .B(new_n615), .C1(new_n595), .C2(new_n617), .ZN(new_n618));
  AOI211_X1 g0418(.A(G179), .B(new_n593), .C1(new_n587), .C2(new_n279), .ZN(new_n619));
  AOI21_X1  g0419(.A(G169), .B1(new_n588), .B2(new_n594), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n614), .A2(new_n256), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n598), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n581), .A2(new_n618), .A3(new_n624), .ZN(new_n625));
  AND4_X1   g0425(.A1(new_n445), .A2(new_n507), .A3(new_n545), .A4(new_n625), .ZN(G372));
  AND2_X1   g0426(.A1(new_n421), .A2(new_n422), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n306), .A2(new_n307), .A3(KEYINPUT14), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n307), .B1(new_n306), .B2(KEYINPUT14), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n265), .B1(new_n630), .B2(new_n302), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n310), .A2(KEYINPUT74), .A3(new_n311), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n263), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n442), .B1(new_n323), .B2(new_n324), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n627), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  XNOR2_X1  g0435(.A(new_n410), .B(KEYINPUT18), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n370), .B1(new_n637), .B2(new_n367), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n565), .A2(KEYINPUT84), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT84), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n563), .A2(new_n564), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n572), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n303), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n570), .A2(new_n440), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT85), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n643), .A2(KEYINPUT85), .A3(new_n644), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n328), .B1(new_n554), .B2(new_n555), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n559), .B1(new_n649), .B2(new_n557), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n647), .A2(new_n648), .B1(new_n579), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n577), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n580), .A2(new_n652), .A3(new_n644), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n572), .A2(new_n573), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n354), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n570), .A2(G190), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n650), .A2(new_n655), .A3(new_n561), .A4(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n621), .A2(new_n653), .A3(new_n657), .A4(new_n623), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n651), .B1(KEYINPUT26), .B2(new_n658), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n643), .A2(KEYINPUT85), .A3(new_n644), .ZN(new_n660));
  AOI21_X1  g0460(.A(KEYINPUT85), .B1(new_n643), .B2(new_n644), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n580), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n593), .B1(new_n587), .B2(new_n279), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n440), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(G169), .B2(new_n663), .ZN(new_n665));
  OAI21_X1  g0465(.A(KEYINPUT86), .B1(new_n665), .B2(new_n615), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n650), .A2(new_n561), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n642), .A2(new_n354), .ZN(new_n668));
  OR3_X1    g0468(.A1(new_n667), .A2(new_n668), .A3(new_n574), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT86), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n621), .A2(new_n670), .A3(new_n623), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n662), .A2(new_n666), .A3(new_n669), .A4(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n659), .B1(KEYINPUT26), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n536), .A2(new_n540), .A3(new_n542), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n498), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n503), .A2(new_n505), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n472), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n677), .A2(new_n624), .A3(new_n618), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n662), .A2(new_n669), .ZN(new_n679));
  NOR3_X1   g0479(.A1(new_n675), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n673), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n445), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n638), .A2(new_n682), .ZN(G369));
  NAND3_X1  g0483(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(G213), .A3(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(G343), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n502), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT87), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n495), .A2(new_n497), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n502), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n677), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT88), .ZN(new_n695));
  OR3_X1    g0495(.A1(new_n691), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n695), .B1(new_n691), .B2(new_n694), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n498), .A2(new_n689), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n528), .A2(new_n689), .ZN(new_n701));
  MUX2_X1   g0501(.A(new_n674), .B(new_n545), .S(new_n701), .Z(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G330), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n689), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n498), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n674), .A2(new_n706), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n696), .A2(new_n697), .A3(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n705), .A2(new_n707), .A3(new_n710), .ZN(G399));
  NOR2_X1   g0511(.A1(new_n210), .A2(G41), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n550), .A2(G116), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n713), .A2(G1), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n715), .B1(new_n214), .B2(new_n713), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT28), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT29), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT26), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n666), .A2(new_n671), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n667), .A2(new_n668), .A3(new_n574), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n647), .A2(new_n648), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n721), .B1(new_n722), .B2(new_n580), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n719), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n662), .B1(new_n658), .B2(KEYINPUT26), .ZN(new_n725));
  OAI21_X1  g0525(.A(KEYINPUT91), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n538), .B(new_n541), .ZN(new_n727));
  INV_X1    g0527(.A(new_n497), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n728), .B1(G169), .B2(new_n494), .ZN(new_n729));
  OAI211_X1 g0529(.A(new_n727), .B(new_n536), .C1(new_n729), .C2(new_n472), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n618), .A2(new_n624), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n730), .A2(new_n677), .A3(new_n731), .A4(new_n723), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n725), .B1(new_n672), .B2(KEYINPUT26), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT91), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n726), .A2(new_n732), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n718), .B1(new_n736), .B2(new_n706), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n681), .A2(new_n718), .A3(new_n706), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AND3_X1   g0539(.A1(new_n537), .A2(new_n440), .A3(new_n642), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT89), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n740), .A2(new_n741), .A3(new_n504), .A4(new_n595), .ZN(new_n742));
  AOI21_X1  g0542(.A(G179), .B1(new_n509), .B2(new_n514), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n504), .A2(new_n743), .A3(new_n595), .A4(new_n642), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(KEYINPUT89), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT30), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n496), .A2(new_n663), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n570), .A2(new_n509), .A3(new_n514), .A4(G179), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n748), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n750), .A2(KEYINPUT30), .A3(new_n496), .A4(new_n663), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n742), .A2(new_n745), .A3(new_n749), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(new_n689), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT31), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(KEYINPUT90), .ZN(new_n756));
  AOI21_X1  g0556(.A(KEYINPUT31), .B1(new_n752), .B2(new_n689), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT90), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n507), .A2(new_n625), .A3(new_n545), .A4(new_n706), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n751), .A2(new_n744), .A3(new_n749), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n761), .A2(KEYINPUT31), .A3(new_n689), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n756), .A2(new_n759), .A3(new_n760), .A4(new_n762), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n763), .A2(G330), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n739), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n717), .B1(new_n767), .B2(G1), .ZN(G364));
  OR3_X1    g0568(.A1(KEYINPUT95), .A2(G13), .A3(G33), .ZN(new_n769));
  OAI21_X1  g0569(.A(KEYINPUT95), .B1(G13), .B2(G33), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n216), .B1(G20), .B2(new_n303), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n210), .A2(new_n380), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT94), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G355), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(G116), .B2(new_n211), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n210), .A2(new_n272), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(G45), .B2(new_n214), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(G45), .B2(new_n243), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n775), .B1(new_n779), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n207), .A2(G13), .ZN(new_n784));
  OAI21_X1  g0584(.A(G1), .B1(new_n784), .B2(new_n283), .ZN(new_n785));
  OR3_X1    g0585(.A1(new_n712), .A2(KEYINPUT93), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(KEYINPUT93), .B1(new_n712), .B2(new_n785), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n783), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT96), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n207), .A2(G190), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G179), .A2(G200), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G159), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT32), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n207), .A2(new_n440), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR3_X1   g0599(.A1(new_n799), .A2(new_n416), .A3(new_n414), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n793), .A2(G190), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G20), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n801), .A2(new_n202), .B1(new_n520), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n797), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(G200), .B1(new_n799), .B2(KEYINPUT97), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(KEYINPUT97), .B2(new_n799), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n416), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n808), .A2(G190), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n806), .B1(new_n383), .B2(new_n810), .C1(new_n344), .C2(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n354), .A2(new_n440), .A3(new_n792), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(G107), .ZN(new_n816));
  NOR4_X1   g0616(.A1(new_n353), .A2(new_n207), .A3(G179), .A4(new_n416), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(G87), .ZN(new_n818));
  NOR3_X1   g0618(.A1(new_n799), .A2(G190), .A3(new_n414), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n380), .B1(new_n819), .B2(G68), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n816), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n813), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n794), .B(KEYINPUT98), .ZN(new_n823));
  AOI22_X1  g0623(.A1(G283), .A2(new_n815), .B1(new_n823), .B2(G329), .ZN(new_n824));
  INV_X1    g0624(.A(G303), .ZN(new_n825));
  INV_X1    g0625(.A(new_n817), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n809), .A2(G322), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n272), .B1(new_n800), .B2(G326), .ZN(new_n829));
  XNOR2_X1  g0629(.A(KEYINPUT33), .B(G317), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n819), .A2(new_n830), .B1(new_n803), .B2(G294), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n828), .A2(new_n829), .A3(new_n831), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n827), .B(new_n832), .C1(G311), .C2(new_n811), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n822), .B1(new_n834), .B2(KEYINPUT99), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(KEYINPUT99), .B2(new_n834), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n791), .B1(new_n836), .B2(new_n774), .ZN(new_n837));
  INV_X1    g0637(.A(new_n773), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n837), .B1(new_n702), .B2(new_n838), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n839), .B(KEYINPUT100), .Z(new_n840));
  XNOR2_X1  g0640(.A(new_n703), .B(KEYINPUT92), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n841), .B(new_n788), .C1(G330), .C2(new_n702), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n840), .A2(new_n842), .ZN(G396));
  NOR2_X1   g0643(.A1(new_n442), .A2(new_n689), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n432), .A2(new_n689), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n439), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n844), .B1(new_n846), .B2(new_n442), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n681), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n848), .B1(new_n849), .B2(new_n689), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n706), .B(new_n847), .C1(new_n673), .C2(new_n680), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n789), .B1(new_n852), .B2(new_n765), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n765), .B2(new_n852), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n771), .A2(new_n774), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n788), .B1(new_n252), .B2(new_n855), .ZN(new_n856));
  AOI22_X1  g0656(.A1(G137), .A2(new_n800), .B1(new_n819), .B2(G150), .ZN(new_n857));
  INV_X1    g0657(.A(G159), .ZN(new_n858));
  XOR2_X1   g0658(.A(KEYINPUT101), .B(G143), .Z(new_n859));
  OAI221_X1 g0659(.A(new_n857), .B1(new_n812), .B2(new_n858), .C1(new_n810), .C2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT34), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n815), .A2(G68), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n823), .A2(G132), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n380), .B1(new_n803), .B2(G58), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n817), .A2(G50), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n863), .A2(new_n864), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n860), .A2(new_n861), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n815), .A2(G87), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n435), .B2(new_n826), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(G311), .B2(new_n823), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n272), .B1(new_n803), .B2(G97), .ZN(new_n873));
  AOI22_X1  g0673(.A1(G303), .A2(new_n800), .B1(new_n819), .B2(G283), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n873), .B(new_n874), .C1(new_n812), .C2(new_n517), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(G294), .B2(new_n809), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n868), .A2(new_n869), .B1(new_n872), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n774), .ZN(new_n878));
  OAI221_X1 g0678(.A(new_n856), .B1(new_n877), .B2(new_n878), .C1(new_n772), .C2(new_n847), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n854), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(G384));
  INV_X1    g0681(.A(new_n611), .ZN(new_n882));
  OR2_X1    g0682(.A1(new_n882), .A2(KEYINPUT35), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(KEYINPUT35), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n883), .A2(new_n884), .A3(G116), .A4(new_n217), .ZN(new_n885));
  XOR2_X1   g0685(.A(new_n885), .B(KEYINPUT36), .Z(new_n886));
  OAI211_X1 g0686(.A(new_n219), .B(new_n215), .C1(new_n383), .C2(new_n247), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n202), .A2(G68), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n206), .B(G13), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n752), .A2(KEYINPUT31), .A3(new_n689), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n760), .A2(new_n755), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n445), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n893), .B(KEYINPUT102), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n263), .A2(new_n706), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n313), .A2(new_n325), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n631), .A2(new_n632), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n315), .A2(KEYINPUT72), .A3(new_n320), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT72), .B1(new_n315), .B2(new_n320), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n264), .B(new_n689), .C1(new_n898), .C2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n897), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT38), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT37), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n418), .A2(new_n376), .A3(new_n394), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n906), .A2(new_n410), .ZN(new_n907));
  INV_X1    g0707(.A(new_n687), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n395), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n905), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n408), .A2(new_n909), .A3(new_n905), .A4(new_n419), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n909), .B1(new_n636), .B2(new_n627), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n904), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n394), .A2(new_n374), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n908), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n413), .B2(new_n423), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n916), .A2(new_n407), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n917), .A2(new_n920), .A3(new_n419), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n911), .B1(new_n921), .B2(new_n905), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n919), .A2(KEYINPUT38), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n915), .A2(new_n923), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n892), .A2(new_n847), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n903), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(KEYINPUT40), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT38), .B1(new_n919), .B2(new_n922), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT40), .B1(new_n929), .B2(new_n923), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n903), .A2(new_n925), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n894), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n894), .A2(new_n932), .ZN(new_n934));
  INV_X1    g0734(.A(G330), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n844), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n851), .A2(new_n937), .ZN(new_n938));
  NOR3_X1   g0738(.A1(new_n633), .A2(new_n901), .A3(new_n895), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n896), .B1(new_n313), .B2(new_n325), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n923), .B2(new_n929), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT39), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n924), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n929), .A2(KEYINPUT39), .A3(new_n923), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n633), .A2(new_n706), .ZN(new_n947));
  OAI22_X1  g0747(.A1(new_n946), .A2(new_n947), .B1(new_n636), .B2(new_n908), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n942), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n445), .B1(new_n737), .B2(new_n738), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n638), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n949), .B(new_n951), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n936), .A2(new_n952), .B1(G1), .B2(new_n784), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT103), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n953), .A2(new_n954), .B1(new_n952), .B2(new_n936), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n953), .A2(new_n954), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n890), .B1(new_n955), .B2(new_n956), .ZN(G367));
  OAI21_X1  g0757(.A(new_n710), .B1(new_n700), .B2(new_n709), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n958), .A2(new_n703), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n841), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n961), .A2(new_n766), .ZN(new_n962));
  INV_X1    g0762(.A(new_n731), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n615), .A2(new_n706), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n963), .A2(new_n964), .B1(new_n624), .B2(new_n706), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT104), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n966), .A2(new_n707), .A3(new_n710), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT45), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n967), .A2(new_n968), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n710), .A2(new_n707), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT104), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n965), .B(new_n972), .ZN(new_n973));
  AND3_X1   g0773(.A1(new_n971), .A2(KEYINPUT44), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(KEYINPUT44), .B1(new_n971), .B2(new_n973), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n969), .A2(new_n970), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n976), .A2(new_n704), .A3(new_n700), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n705), .B1(new_n974), .B2(new_n975), .C1(new_n969), .C2(new_n970), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n962), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n767), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n712), .B(KEYINPUT41), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n785), .B(KEYINPUT106), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n973), .A2(new_n710), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n624), .B1(new_n973), .B2(new_n693), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n985), .A2(KEYINPUT42), .B1(new_n986), .B2(new_n706), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n985), .A2(KEYINPUT42), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n562), .A2(new_n706), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n651), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n679), .B2(new_n990), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT43), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n992), .A2(KEYINPUT43), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n989), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n705), .A2(new_n973), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n987), .A2(new_n988), .A3(new_n994), .A4(new_n993), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(KEYINPUT105), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n997), .A2(new_n999), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n998), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT105), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n997), .A2(new_n1005), .A3(new_n998), .A4(new_n999), .ZN(new_n1006));
  AND3_X1   g0806(.A1(new_n1001), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n984), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(G317), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n819), .ZN(new_n1010));
  INV_X1    g0810(.A(G294), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n380), .B1(new_n794), .B2(new_n1009), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n814), .A2(new_n520), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n800), .A2(G311), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n435), .B2(new_n804), .ZN(new_n1015));
  NOR3_X1   g0815(.A1(new_n1012), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G283), .A2(new_n811), .B1(new_n809), .B2(G303), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT46), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n826), .B2(new_n517), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n817), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1016), .A2(new_n1017), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n804), .A2(new_n247), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n801), .A2(new_n859), .B1(new_n1010), .B2(new_n858), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1022), .B(new_n1023), .C1(G150), .C2(new_n809), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n272), .B1(new_n814), .B2(new_n344), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT107), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1024), .B(new_n1026), .C1(new_n202), .C2(new_n812), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n817), .A2(G58), .B1(G137), .B2(new_n795), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT108), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1021), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT109), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT47), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n774), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n993), .A2(new_n773), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n775), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n210), .B2(new_n426), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n231), .A2(new_n780), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n788), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1033), .A2(new_n1034), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1008), .A2(new_n1039), .ZN(G387));
  INV_X1    g0840(.A(new_n983), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n959), .A2(new_n960), .A3(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n780), .B1(new_n236), .B2(new_n283), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n777), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1043), .B1(new_n714), .B2(new_n1044), .ZN(new_n1045));
  OR3_X1    g0845(.A1(new_n372), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1046));
  OAI21_X1  g0846(.A(KEYINPUT50), .B1(new_n372), .B2(G50), .ZN(new_n1047));
  AOI21_X1  g0847(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1046), .A2(new_n714), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n1045), .A2(new_n1049), .B1(new_n435), .B2(new_n210), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n789), .B1(new_n1050), .B2(new_n1035), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n826), .A2(new_n344), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(G150), .B2(new_n795), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT110), .Z(new_n1054));
  OAI21_X1  g0854(.A(new_n272), .B1(new_n801), .B2(new_n858), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1010), .A2(new_n372), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n804), .A2(new_n425), .ZN(new_n1057));
  NOR4_X1   g0857(.A1(new_n1055), .A2(new_n1056), .A3(new_n1013), .A4(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(G50), .A2(new_n809), .B1(new_n811), .B2(G68), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1054), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n272), .B1(new_n795), .B2(G326), .ZN(new_n1061));
  INV_X1    g0861(.A(G283), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n826), .A2(new_n1011), .B1(new_n1062), .B2(new_n804), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(G322), .A2(new_n800), .B1(new_n819), .B2(G311), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1064), .B1(new_n812), .B2(new_n825), .C1(new_n1009), .C2(new_n810), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT48), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1063), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n1066), .B2(new_n1065), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT49), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1061), .B1(new_n517), .B2(new_n814), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1060), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1051), .B1(new_n1072), .B2(new_n774), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n700), .B2(new_n838), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n1042), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n767), .B1(new_n960), .B2(new_n959), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n712), .B1(new_n961), .B2(new_n766), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1075), .B1(new_n1076), .B2(new_n1077), .ZN(G393));
  NAND2_X1  g0878(.A1(new_n977), .A2(new_n978), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n766), .B2(new_n961), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1080), .A2(new_n712), .A3(new_n979), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n977), .A2(new_n978), .A3(new_n1041), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n775), .B1(new_n520), .B2(new_n211), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n240), .B2(new_n780), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n819), .A2(G50), .B1(new_n803), .B2(G77), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n812), .B2(new_n372), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT111), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n809), .A2(G159), .B1(G150), .B2(new_n800), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT51), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n859), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n380), .B1(new_n1090), .B2(new_n795), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n870), .B(new_n1091), .C1(new_n247), .C2(new_n826), .ZN(new_n1092));
  OR3_X1    g0892(.A1(new_n1087), .A2(new_n1089), .A3(new_n1092), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n809), .A2(G311), .B1(G317), .B2(new_n800), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT113), .ZN(new_n1095));
  XOR2_X1   g0895(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n1096));
  XNOR2_X1  g0896(.A(new_n1095), .B(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n272), .B1(new_n795), .B2(G322), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n517), .B2(new_n804), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n816), .B1(new_n1062), .B2(new_n826), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1099), .B(new_n1100), .C1(G303), .C2(new_n819), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n1011), .B2(new_n812), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1093), .B1(new_n1097), .B2(new_n1102), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n788), .B(new_n1084), .C1(new_n1103), .C2(new_n774), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n966), .B2(new_n838), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1082), .A2(KEYINPUT114), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(KEYINPUT114), .B1(new_n1082), .B2(new_n1105), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1081), .B1(new_n1107), .B2(new_n1108), .ZN(G390));
  AOI21_X1  g0909(.A(new_n272), .B1(new_n803), .B2(G77), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(G283), .A2(new_n800), .B1(new_n819), .B2(G107), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1110), .B(new_n1111), .C1(new_n810), .C2(new_n517), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G97), .B2(new_n811), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n823), .A2(G294), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1113), .A2(new_n818), .A3(new_n863), .A4(new_n1114), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n819), .A2(G137), .B1(new_n803), .B2(G159), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(KEYINPUT54), .B(G143), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1116), .B1(new_n812), .B2(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1118), .B(KEYINPUT117), .ZN(new_n1119));
  INV_X1    g0919(.A(G128), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n272), .B1(new_n814), .B2(new_n202), .C1(new_n801), .C2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(G125), .B2(new_n823), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n817), .A2(G150), .ZN(new_n1123));
  OR2_X1    g0923(.A1(new_n1123), .A2(KEYINPUT53), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n809), .A2(G132), .B1(KEYINPUT53), .B2(new_n1123), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1119), .A2(new_n1122), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1115), .B1(new_n1127), .B2(KEYINPUT118), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT118), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n774), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n855), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1131), .B(new_n789), .C1(new_n329), .C2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(new_n946), .B2(new_n771), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n892), .A2(G330), .A3(new_n847), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n897), .B2(new_n902), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n919), .A2(KEYINPUT38), .A3(new_n922), .ZN(new_n1138));
  NOR3_X1   g0938(.A1(new_n1138), .A2(new_n928), .A3(new_n943), .ZN(new_n1139));
  AOI21_X1  g0939(.A(KEYINPUT39), .B1(new_n915), .B2(new_n923), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(new_n941), .B2(new_n947), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n924), .A2(new_n947), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n846), .A2(new_n442), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n1145));
  AOI211_X1 g0945(.A(KEYINPUT91), .B(new_n725), .C1(KEYINPUT26), .C2(new_n672), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n706), .B(new_n1144), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n937), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1143), .B1(new_n1148), .B2(new_n903), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1137), .B1(new_n1142), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1148), .A2(new_n903), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1143), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n903), .A2(new_n764), .A3(new_n847), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n897), .A2(new_n902), .B1(new_n937), .B2(new_n851), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n947), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n946), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1153), .A2(new_n1154), .A3(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1150), .A2(new_n1041), .A3(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT116), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1159), .B(new_n1160), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n760), .B(new_n762), .C1(new_n758), .C2(new_n757), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n759), .ZN(new_n1163));
  OAI211_X1 g0963(.A(G330), .B(new_n847), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1164));
  AND3_X1   g0964(.A1(new_n1164), .A2(new_n897), .A3(new_n902), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n938), .B1(new_n1165), .B2(new_n1137), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1148), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n897), .A2(new_n902), .A3(new_n1136), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1154), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n445), .A2(G330), .A3(new_n892), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n950), .A2(new_n638), .A3(new_n1171), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1150), .A2(new_n1170), .A3(new_n1158), .A4(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1173), .A2(KEYINPUT115), .A3(new_n712), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1150), .A2(new_n1158), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1174), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(KEYINPUT115), .B1(new_n1173), .B2(new_n712), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1135), .B(new_n1161), .C1(new_n1178), .C2(new_n1179), .ZN(G378));
  INV_X1    g0980(.A(G132), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n826), .A2(new_n1117), .B1(new_n1010), .B2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(G137), .B2(new_n811), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n1120), .B2(new_n810), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n800), .A2(G125), .B1(new_n803), .B2(G150), .ZN(new_n1185));
  XOR2_X1   g0985(.A(new_n1185), .B(KEYINPUT119), .Z(new_n1186));
  NOR2_X1   g0986(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(G33), .A2(G41), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT120), .B(G124), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1191), .B1(new_n794), .B2(new_n1192), .C1(new_n814), .C2(new_n858), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1189), .A2(new_n1190), .A3(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n272), .A2(G41), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n804), .B2(new_n247), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n1010), .A2(new_n520), .B1(new_n801), .B2(new_n517), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1196), .B(new_n1197), .C1(G107), .C2(new_n809), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n425), .B2(new_n812), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n823), .A2(G283), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n814), .A2(new_n383), .ZN(new_n1201));
  NOR4_X1   g1001(.A1(new_n1199), .A2(new_n1052), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  AND2_X1   g1002(.A1(new_n1202), .A2(KEYINPUT58), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1202), .A2(KEYINPUT58), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(new_n1195), .A2(G50), .A3(new_n1191), .ZN(new_n1205));
  NOR4_X1   g1005(.A1(new_n1194), .A2(new_n1203), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n789), .B1(G50), .B2(new_n1132), .C1(new_n1206), .C2(new_n878), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n367), .A2(new_n371), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n687), .B1(new_n357), .B2(new_n339), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  OR3_X1    g1013(.A1(new_n1210), .A2(new_n1211), .A3(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1213), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1215));
  AND2_X1   g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1207), .B1(new_n1216), .B2(new_n771), .ZN(new_n1217));
  AND2_X1   g1017(.A1(new_n903), .A2(new_n925), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1218), .A2(new_n930), .B1(new_n926), .B2(KEYINPUT40), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1216), .B1(new_n1219), .B2(new_n935), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n932), .A2(G330), .A3(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n949), .B1(new_n1220), .B2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1220), .A2(new_n949), .A3(new_n1222), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1217), .B1(new_n1226), .B2(new_n1041), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n1173), .A2(KEYINPUT121), .A3(new_n1172), .ZN(new_n1228));
  AOI21_X1  g1028(.A(KEYINPUT121), .B1(new_n1173), .B2(new_n1172), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1225), .ZN(new_n1231));
  OAI21_X1  g1031(.A(KEYINPUT57), .B1(new_n1231), .B2(new_n1223), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n712), .B1(new_n1230), .B2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1170), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1172), .B1(new_n1175), .B2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT121), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1173), .A2(KEYINPUT121), .A3(new_n1172), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(KEYINPUT57), .B1(new_n1239), .B2(new_n1226), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1227), .B1(new_n1233), .B2(new_n1240), .ZN(G375));
  OR2_X1    g1041(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1242), .A2(new_n981), .A3(new_n1176), .ZN(new_n1243));
  XOR2_X1   g1043(.A(new_n1243), .B(KEYINPUT122), .Z(new_n1244));
  AOI21_X1  g1044(.A(new_n788), .B1(new_n247), .B2(new_n855), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(KEYINPUT124), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(G294), .A2(new_n800), .B1(new_n819), .B2(G116), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n812), .B2(new_n435), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(new_n1248), .B(KEYINPUT125), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n272), .B(new_n1057), .C1(G77), .C2(new_n815), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n823), .A2(G303), .B1(G97), .B2(new_n817), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1250), .B(new_n1251), .C1(new_n1062), .C2(new_n810), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n272), .B1(new_n801), .B2(new_n1181), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n1010), .A2(new_n1117), .B1(new_n202), .B2(new_n804), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n1253), .B(new_n1254), .C1(G150), .C2(new_n811), .ZN(new_n1255));
  INV_X1    g1055(.A(G137), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1255), .B1(new_n1256), .B2(new_n810), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1201), .B1(G128), .B2(new_n823), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1258), .B1(new_n858), .B2(new_n826), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n1249), .A2(new_n1252), .B1(new_n1257), .B2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1246), .B1(new_n1260), .B2(new_n774), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1261), .B1(new_n903), .B2(new_n772), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n983), .B(KEYINPUT123), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1262), .B1(new_n1234), .B2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1244), .A2(new_n1265), .ZN(G381));
  INV_X1    g1066(.A(G396), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1075), .B(new_n1267), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1268));
  OR4_X1    g1068(.A1(G384), .A2(G387), .A3(G390), .A4(new_n1268), .ZN(new_n1269));
  OR4_X1    g1069(.A1(G378), .A2(new_n1269), .A3(G375), .A4(G381), .ZN(G407));
  INV_X1    g1070(.A(G378), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n688), .A2(G213), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1274));
  OAI211_X1 g1074(.A(G407), .B(G213), .C1(G375), .C2(new_n1274), .ZN(G409));
  NAND2_X1  g1075(.A1(G393), .A2(G396), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1268), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(G390), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1108), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n1106), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1277), .B1(new_n1281), .B2(new_n1081), .ZN(new_n1282));
  OAI21_X1  g1082(.A(G387), .B1(new_n1279), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(G390), .A2(new_n1278), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1039), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1285), .B1(new_n984), .B2(new_n1007), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1281), .A2(new_n1081), .A3(new_n1277), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1284), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1283), .A2(new_n1288), .ZN(new_n1289));
  OAI211_X1 g1089(.A(G378), .B(new_n1227), .C1(new_n1233), .C2(new_n1240), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1231), .A2(new_n1223), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n981), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1291), .B1(new_n1292), .B2(new_n1263), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1271), .B1(new_n1293), .B2(new_n1217), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1290), .A2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1272), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1176), .A2(KEYINPUT60), .ZN(new_n1297));
  AND2_X1   g1097(.A1(new_n1297), .A2(new_n1242), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n712), .B1(new_n1297), .B2(new_n1242), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n880), .B1(new_n1300), .B2(new_n1264), .ZN(new_n1301));
  OAI211_X1 g1101(.A(G384), .B(new_n1265), .C1(new_n1298), .C2(new_n1299), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1273), .A2(G2897), .ZN(new_n1303));
  AND3_X1   g1103(.A1(new_n1301), .A2(new_n1302), .A3(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1303), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(KEYINPUT61), .B1(new_n1296), .B2(new_n1306), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1295), .A2(new_n1308), .A3(new_n1272), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(KEYINPUT62), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1307), .A2(new_n1310), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1309), .A2(KEYINPUT62), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1289), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  AND3_X1   g1113(.A1(new_n1301), .A2(new_n1302), .A3(KEYINPUT63), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1295), .A2(new_n1272), .A3(new_n1314), .ZN(new_n1315));
  AND2_X1   g1115(.A1(new_n1283), .A2(new_n1288), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  XNOR2_X1  g1117(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1273), .B1(new_n1290), .B2(new_n1294), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1319), .B1(new_n1320), .B2(new_n1308), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1317), .A2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(KEYINPUT127), .B1(new_n1322), .B2(new_n1307), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1309), .A2(new_n1318), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1289), .B1(new_n1320), .B2(new_n1314), .ZN(new_n1325));
  AND4_X1   g1125(.A1(KEYINPUT127), .A2(new_n1307), .A3(new_n1324), .A4(new_n1325), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1313), .B1(new_n1323), .B2(new_n1326), .ZN(G405));
  XNOR2_X1  g1127(.A(G375), .B(G378), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1308), .ZN(new_n1329));
  AND2_X1   g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1331));
  OR3_X1    g1131(.A1(new_n1330), .A2(new_n1331), .A3(new_n1289), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1289), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1332), .A2(new_n1333), .ZN(G402));
endmodule


