

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U553 ( .A1(n530), .A2(n529), .ZN(G160) );
  XNOR2_X1 U554 ( .A(n690), .B(n689), .ZN(n693) );
  NAND2_X1 U555 ( .A1(n718), .A2(G2072), .ZN(n690) );
  INV_X1 U556 ( .A(n807), .ZN(n759) );
  XOR2_X1 U557 ( .A(G543), .B(KEYINPUT0), .Z(n518) );
  INV_X1 U558 ( .A(KEYINPUT27), .ZN(n689) );
  INV_X1 U559 ( .A(KEYINPUT92), .ZN(n694) );
  XNOR2_X1 U560 ( .A(KEYINPUT91), .B(n742), .ZN(n718) );
  INV_X1 U561 ( .A(KEYINPUT29), .ZN(n716) );
  XNOR2_X1 U562 ( .A(n717), .B(n716), .ZN(n722) );
  AND2_X1 U563 ( .A1(n741), .A2(n735), .ZN(n736) );
  AND2_X1 U564 ( .A1(n749), .A2(n748), .ZN(n751) );
  NAND2_X1 U565 ( .A1(n688), .A2(n765), .ZN(n742) );
  OR2_X1 U566 ( .A1(n534), .A2(n638), .ZN(n535) );
  NOR2_X1 U567 ( .A1(n764), .A2(n763), .ZN(n799) );
  XOR2_X1 U568 ( .A(KEYINPUT15), .B(n585), .Z(n959) );
  AND2_X2 U569 ( .A1(n524), .A2(n523), .ZN(n883) );
  XOR2_X1 U570 ( .A(KEYINPUT1), .B(n531), .Z(n658) );
  NOR2_X1 U571 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U572 ( .A1(G2104), .A2(G2105), .ZN(n519) );
  XOR2_X1 U573 ( .A(KEYINPUT17), .B(n519), .Z(n520) );
  XNOR2_X1 U574 ( .A(KEYINPUT66), .B(n520), .ZN(n768) );
  NAND2_X1 U575 ( .A1(G137), .A2(n768), .ZN(n530) );
  XNOR2_X1 U576 ( .A(KEYINPUT64), .B(G2104), .ZN(n524) );
  INV_X1 U577 ( .A(G2105), .ZN(n523) );
  NAND2_X1 U578 ( .A1(G101), .A2(n883), .ZN(n521) );
  XNOR2_X1 U579 ( .A(n521), .B(KEYINPUT23), .ZN(n528) );
  NAND2_X1 U580 ( .A1(G2105), .A2(G2104), .ZN(n522) );
  XNOR2_X1 U581 ( .A(n522), .B(KEYINPUT65), .ZN(n887) );
  NAND2_X1 U582 ( .A1(G113), .A2(n887), .ZN(n526) );
  NOR2_X2 U583 ( .A1(n524), .A2(n523), .ZN(n888) );
  NAND2_X1 U584 ( .A1(G125), .A2(n888), .ZN(n525) );
  NAND2_X1 U585 ( .A1(n526), .A2(n525), .ZN(n527) );
  INV_X1 U586 ( .A(G651), .ZN(n534) );
  NOR2_X1 U587 ( .A1(G543), .A2(n534), .ZN(n531) );
  NAND2_X1 U588 ( .A1(G64), .A2(n658), .ZN(n533) );
  XOR2_X1 U589 ( .A(KEYINPUT67), .B(n518), .Z(n638) );
  NOR2_X1 U590 ( .A1(G651), .A2(n638), .ZN(n653) );
  NAND2_X1 U591 ( .A1(G52), .A2(n653), .ZN(n532) );
  NAND2_X1 U592 ( .A1(n533), .A2(n532), .ZN(n540) );
  NOR2_X1 U593 ( .A1(G651), .A2(G543), .ZN(n652) );
  NAND2_X1 U594 ( .A1(G90), .A2(n652), .ZN(n537) );
  XOR2_X1 U595 ( .A(KEYINPUT68), .B(n535), .Z(n651) );
  NAND2_X1 U596 ( .A1(G77), .A2(n651), .ZN(n536) );
  NAND2_X1 U597 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U598 ( .A(KEYINPUT9), .B(n538), .Z(n539) );
  NOR2_X1 U599 ( .A1(n540), .A2(n539), .ZN(G171) );
  XOR2_X1 U600 ( .A(G2443), .B(G2446), .Z(n542) );
  XNOR2_X1 U601 ( .A(G2427), .B(G2451), .ZN(n541) );
  XNOR2_X1 U602 ( .A(n542), .B(n541), .ZN(n548) );
  XOR2_X1 U603 ( .A(G2430), .B(G2454), .Z(n544) );
  XNOR2_X1 U604 ( .A(G1341), .B(G1348), .ZN(n543) );
  XNOR2_X1 U605 ( .A(n544), .B(n543), .ZN(n546) );
  XOR2_X1 U606 ( .A(G2435), .B(G2438), .Z(n545) );
  XNOR2_X1 U607 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U608 ( .A(n548), .B(n547), .Z(n549) );
  AND2_X1 U609 ( .A1(G14), .A2(n549), .ZN(G401) );
  AND2_X1 U610 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U611 ( .A(G57), .ZN(G237) );
  INV_X1 U612 ( .A(G132), .ZN(G219) );
  INV_X1 U613 ( .A(G82), .ZN(G220) );
  NAND2_X1 U614 ( .A1(G138), .A2(n768), .ZN(n551) );
  NAND2_X1 U615 ( .A1(n887), .A2(G114), .ZN(n550) );
  NAND2_X1 U616 ( .A1(n551), .A2(n550), .ZN(n555) );
  NAND2_X1 U617 ( .A1(G126), .A2(n888), .ZN(n553) );
  NAND2_X1 U618 ( .A1(G102), .A2(n883), .ZN(n552) );
  NAND2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U620 ( .A1(n555), .A2(n554), .ZN(G164) );
  NAND2_X1 U621 ( .A1(n652), .A2(G89), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(KEYINPUT4), .ZN(n558) );
  NAND2_X1 U623 ( .A1(G76), .A2(n651), .ZN(n557) );
  NAND2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U625 ( .A(KEYINPUT5), .B(n559), .ZN(n565) );
  NAND2_X1 U626 ( .A1(G63), .A2(n658), .ZN(n561) );
  NAND2_X1 U627 ( .A1(G51), .A2(n653), .ZN(n560) );
  NAND2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n563) );
  XOR2_X1 U629 ( .A(KEYINPUT6), .B(KEYINPUT72), .Z(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n564) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(KEYINPUT7), .B(n566), .ZN(G168) );
  XOR2_X1 U633 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U634 ( .A1(G7), .A2(G661), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n567), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U636 ( .A(G223), .ZN(n832) );
  NAND2_X1 U637 ( .A1(n832), .A2(G567), .ZN(n568) );
  XOR2_X1 U638 ( .A(KEYINPUT11), .B(n568), .Z(G234) );
  NAND2_X1 U639 ( .A1(n652), .A2(G81), .ZN(n569) );
  XNOR2_X1 U640 ( .A(n569), .B(KEYINPUT12), .ZN(n571) );
  NAND2_X1 U641 ( .A1(G68), .A2(n651), .ZN(n570) );
  NAND2_X1 U642 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U643 ( .A(KEYINPUT13), .B(n572), .ZN(n578) );
  NAND2_X1 U644 ( .A1(G56), .A2(n658), .ZN(n573) );
  XOR2_X1 U645 ( .A(KEYINPUT14), .B(n573), .Z(n576) );
  NAND2_X1 U646 ( .A1(G43), .A2(n653), .ZN(n574) );
  XNOR2_X1 U647 ( .A(KEYINPUT69), .B(n574), .ZN(n575) );
  NOR2_X1 U648 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U649 ( .A1(n578), .A2(n577), .ZN(n954) );
  INV_X1 U650 ( .A(G860), .ZN(n598) );
  OR2_X1 U651 ( .A1(n954), .A2(n598), .ZN(G153) );
  XOR2_X1 U652 ( .A(G171), .B(KEYINPUT70), .Z(G301) );
  INV_X1 U653 ( .A(G868), .ZN(n671) );
  NOR2_X1 U654 ( .A1(G301), .A2(n671), .ZN(n587) );
  NAND2_X1 U655 ( .A1(n651), .A2(G79), .ZN(n580) );
  NAND2_X1 U656 ( .A1(G92), .A2(n652), .ZN(n579) );
  NAND2_X1 U657 ( .A1(n580), .A2(n579), .ZN(n584) );
  NAND2_X1 U658 ( .A1(G66), .A2(n658), .ZN(n582) );
  NAND2_X1 U659 ( .A1(G54), .A2(n653), .ZN(n581) );
  NAND2_X1 U660 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U661 ( .A1(n584), .A2(n583), .ZN(n585) );
  AND2_X1 U662 ( .A1(n671), .A2(n959), .ZN(n586) );
  NOR2_X1 U663 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U664 ( .A(KEYINPUT71), .B(n588), .Z(G284) );
  NAND2_X1 U665 ( .A1(G65), .A2(n658), .ZN(n590) );
  NAND2_X1 U666 ( .A1(G53), .A2(n653), .ZN(n589) );
  NAND2_X1 U667 ( .A1(n590), .A2(n589), .ZN(n594) );
  NAND2_X1 U668 ( .A1(G91), .A2(n652), .ZN(n592) );
  NAND2_X1 U669 ( .A1(G78), .A2(n651), .ZN(n591) );
  NAND2_X1 U670 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U671 ( .A1(n594), .A2(n593), .ZN(n699) );
  INV_X1 U672 ( .A(n699), .ZN(G299) );
  NOR2_X1 U673 ( .A1(G286), .A2(n671), .ZN(n596) );
  NOR2_X1 U674 ( .A1(G868), .A2(G299), .ZN(n595) );
  NOR2_X1 U675 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U676 ( .A(KEYINPUT73), .B(n597), .Z(G297) );
  NAND2_X1 U677 ( .A1(n598), .A2(G559), .ZN(n599) );
  NAND2_X1 U678 ( .A1(n599), .A2(n959), .ZN(n600) );
  XNOR2_X1 U679 ( .A(n600), .B(KEYINPUT16), .ZN(n601) );
  XNOR2_X1 U680 ( .A(KEYINPUT74), .B(n601), .ZN(G148) );
  NOR2_X1 U681 ( .A1(G868), .A2(n954), .ZN(n602) );
  XOR2_X1 U682 ( .A(KEYINPUT75), .B(n602), .Z(n605) );
  NAND2_X1 U683 ( .A1(G868), .A2(n959), .ZN(n603) );
  NOR2_X1 U684 ( .A1(G559), .A2(n603), .ZN(n604) );
  NOR2_X1 U685 ( .A1(n605), .A2(n604), .ZN(G282) );
  XOR2_X1 U686 ( .A(KEYINPUT18), .B(KEYINPUT76), .Z(n607) );
  NAND2_X1 U687 ( .A1(G123), .A2(n888), .ZN(n606) );
  XNOR2_X1 U688 ( .A(n607), .B(n606), .ZN(n610) );
  NAND2_X1 U689 ( .A1(G135), .A2(n768), .ZN(n608) );
  XNOR2_X1 U690 ( .A(KEYINPUT77), .B(n608), .ZN(n609) );
  NOR2_X1 U691 ( .A1(n610), .A2(n609), .ZN(n615) );
  NAND2_X1 U692 ( .A1(G111), .A2(n887), .ZN(n612) );
  NAND2_X1 U693 ( .A1(G99), .A2(n883), .ZN(n611) );
  NAND2_X1 U694 ( .A1(n612), .A2(n611), .ZN(n613) );
  XOR2_X1 U695 ( .A(KEYINPUT78), .B(n613), .Z(n614) );
  NAND2_X1 U696 ( .A1(n615), .A2(n614), .ZN(n616) );
  XOR2_X1 U697 ( .A(KEYINPUT79), .B(n616), .Z(n920) );
  XOR2_X1 U698 ( .A(G2096), .B(KEYINPUT80), .Z(n617) );
  XNOR2_X1 U699 ( .A(n920), .B(n617), .ZN(n619) );
  INV_X1 U700 ( .A(G2100), .ZN(n618) );
  NAND2_X1 U701 ( .A1(n619), .A2(n618), .ZN(G156) );
  NAND2_X1 U702 ( .A1(G67), .A2(n658), .ZN(n620) );
  XNOR2_X1 U703 ( .A(n620), .B(KEYINPUT82), .ZN(n627) );
  NAND2_X1 U704 ( .A1(n653), .A2(G55), .ZN(n622) );
  NAND2_X1 U705 ( .A1(G80), .A2(n651), .ZN(n621) );
  NAND2_X1 U706 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U707 ( .A1(G93), .A2(n652), .ZN(n623) );
  XNOR2_X1 U708 ( .A(KEYINPUT81), .B(n623), .ZN(n624) );
  NOR2_X1 U709 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U710 ( .A1(n627), .A2(n626), .ZN(n670) );
  NAND2_X1 U711 ( .A1(G559), .A2(n959), .ZN(n628) );
  XNOR2_X1 U712 ( .A(n628), .B(n954), .ZN(n668) );
  NOR2_X1 U713 ( .A1(n668), .A2(G860), .ZN(n629) );
  XNOR2_X1 U714 ( .A(n629), .B(KEYINPUT83), .ZN(n630) );
  XNOR2_X1 U715 ( .A(n670), .B(n630), .ZN(G145) );
  NAND2_X1 U716 ( .A1(G86), .A2(n652), .ZN(n632) );
  NAND2_X1 U717 ( .A1(G48), .A2(n653), .ZN(n631) );
  NAND2_X1 U718 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U719 ( .A1(n651), .A2(G73), .ZN(n633) );
  XOR2_X1 U720 ( .A(KEYINPUT2), .B(n633), .Z(n634) );
  NOR2_X1 U721 ( .A1(n635), .A2(n634), .ZN(n637) );
  NAND2_X1 U722 ( .A1(n658), .A2(G61), .ZN(n636) );
  NAND2_X1 U723 ( .A1(n637), .A2(n636), .ZN(G305) );
  NAND2_X1 U724 ( .A1(G87), .A2(n638), .ZN(n639) );
  XNOR2_X1 U725 ( .A(n639), .B(KEYINPUT84), .ZN(n644) );
  NAND2_X1 U726 ( .A1(G49), .A2(n653), .ZN(n641) );
  NAND2_X1 U727 ( .A1(G74), .A2(G651), .ZN(n640) );
  NAND2_X1 U728 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U729 ( .A1(n658), .A2(n642), .ZN(n643) );
  NAND2_X1 U730 ( .A1(n644), .A2(n643), .ZN(G288) );
  NAND2_X1 U731 ( .A1(G88), .A2(n652), .ZN(n646) );
  NAND2_X1 U732 ( .A1(G75), .A2(n651), .ZN(n645) );
  NAND2_X1 U733 ( .A1(n646), .A2(n645), .ZN(n650) );
  NAND2_X1 U734 ( .A1(G62), .A2(n658), .ZN(n648) );
  NAND2_X1 U735 ( .A1(G50), .A2(n653), .ZN(n647) );
  NAND2_X1 U736 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U737 ( .A1(n650), .A2(n649), .ZN(G166) );
  AND2_X1 U738 ( .A1(G72), .A2(n651), .ZN(n657) );
  NAND2_X1 U739 ( .A1(G85), .A2(n652), .ZN(n655) );
  NAND2_X1 U740 ( .A1(G47), .A2(n653), .ZN(n654) );
  NAND2_X1 U741 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U742 ( .A1(n657), .A2(n656), .ZN(n660) );
  NAND2_X1 U743 ( .A1(n658), .A2(G60), .ZN(n659) );
  NAND2_X1 U744 ( .A1(n660), .A2(n659), .ZN(G290) );
  XNOR2_X1 U745 ( .A(KEYINPUT19), .B(KEYINPUT86), .ZN(n662) );
  XNOR2_X1 U746 ( .A(G288), .B(KEYINPUT85), .ZN(n661) );
  XNOR2_X1 U747 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U748 ( .A(G305), .B(n663), .ZN(n665) );
  XNOR2_X1 U749 ( .A(n699), .B(G166), .ZN(n664) );
  XNOR2_X1 U750 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U751 ( .A(n666), .B(G290), .ZN(n667) );
  XNOR2_X1 U752 ( .A(n667), .B(n670), .ZN(n903) );
  XNOR2_X1 U753 ( .A(n668), .B(n903), .ZN(n669) );
  NAND2_X1 U754 ( .A1(n669), .A2(G868), .ZN(n673) );
  NAND2_X1 U755 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U756 ( .A1(n673), .A2(n672), .ZN(G295) );
  NAND2_X1 U757 ( .A1(G2084), .A2(G2078), .ZN(n674) );
  XNOR2_X1 U758 ( .A(n674), .B(KEYINPUT87), .ZN(n675) );
  XNOR2_X1 U759 ( .A(n675), .B(KEYINPUT20), .ZN(n676) );
  NAND2_X1 U760 ( .A1(n676), .A2(G2090), .ZN(n677) );
  XNOR2_X1 U761 ( .A(KEYINPUT21), .B(n677), .ZN(n678) );
  NAND2_X1 U762 ( .A1(n678), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U763 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U764 ( .A1(G220), .A2(G219), .ZN(n679) );
  XOR2_X1 U765 ( .A(KEYINPUT22), .B(n679), .Z(n680) );
  NOR2_X1 U766 ( .A1(G218), .A2(n680), .ZN(n681) );
  NAND2_X1 U767 ( .A1(G96), .A2(n681), .ZN(n837) );
  NAND2_X1 U768 ( .A1(n837), .A2(G2106), .ZN(n685) );
  NAND2_X1 U769 ( .A1(G69), .A2(G120), .ZN(n682) );
  NOR2_X1 U770 ( .A1(G237), .A2(n682), .ZN(n683) );
  NAND2_X1 U771 ( .A1(G108), .A2(n683), .ZN(n838) );
  NAND2_X1 U772 ( .A1(n838), .A2(G567), .ZN(n684) );
  NAND2_X1 U773 ( .A1(n685), .A2(n684), .ZN(n839) );
  NAND2_X1 U774 ( .A1(G483), .A2(G661), .ZN(n686) );
  NOR2_X1 U775 ( .A1(n839), .A2(n686), .ZN(n834) );
  NAND2_X1 U776 ( .A1(n834), .A2(G36), .ZN(G176) );
  INV_X1 U777 ( .A(G166), .ZN(G303) );
  NAND2_X1 U778 ( .A1(G160), .A2(G40), .ZN(n766) );
  INV_X1 U779 ( .A(KEYINPUT90), .ZN(n687) );
  XNOR2_X1 U780 ( .A(n766), .B(n687), .ZN(n688) );
  NOR2_X1 U781 ( .A1(G164), .A2(G1384), .ZN(n765) );
  INV_X1 U782 ( .A(n718), .ZN(n691) );
  NAND2_X1 U783 ( .A1(G1956), .A2(n691), .ZN(n692) );
  NAND2_X1 U784 ( .A1(n693), .A2(n692), .ZN(n695) );
  XNOR2_X1 U785 ( .A(n695), .B(n694), .ZN(n698) );
  NOR2_X1 U786 ( .A1(n698), .A2(n699), .ZN(n697) );
  INV_X1 U787 ( .A(KEYINPUT28), .ZN(n696) );
  XNOR2_X1 U788 ( .A(n697), .B(n696), .ZN(n715) );
  NAND2_X1 U789 ( .A1(n699), .A2(n698), .ZN(n713) );
  INV_X1 U790 ( .A(G1996), .ZN(n1002) );
  NOR2_X1 U791 ( .A1(n742), .A2(n1002), .ZN(n700) );
  XOR2_X1 U792 ( .A(n700), .B(KEYINPUT26), .Z(n702) );
  NAND2_X1 U793 ( .A1(n742), .A2(G1341), .ZN(n701) );
  NAND2_X1 U794 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U795 ( .A1(n954), .A2(n703), .ZN(n704) );
  OR2_X1 U796 ( .A1(n959), .A2(n704), .ZN(n710) );
  NAND2_X1 U797 ( .A1(n959), .A2(n704), .ZN(n708) );
  NAND2_X1 U798 ( .A1(G2067), .A2(n718), .ZN(n706) );
  NAND2_X1 U799 ( .A1(G1348), .A2(n742), .ZN(n705) );
  NAND2_X1 U800 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U801 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U802 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U803 ( .A(KEYINPUT93), .B(n711), .Z(n712) );
  NAND2_X1 U804 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U805 ( .A1(n715), .A2(n714), .ZN(n717) );
  INV_X1 U806 ( .A(G1961), .ZN(n983) );
  NAND2_X1 U807 ( .A1(n983), .A2(n742), .ZN(n720) );
  XNOR2_X1 U808 ( .A(G2078), .B(KEYINPUT25), .ZN(n1009) );
  NAND2_X1 U809 ( .A1(n718), .A2(n1009), .ZN(n719) );
  NAND2_X1 U810 ( .A1(n720), .A2(n719), .ZN(n727) );
  NAND2_X1 U811 ( .A1(n727), .A2(G171), .ZN(n721) );
  NAND2_X1 U812 ( .A1(n722), .A2(n721), .ZN(n733) );
  XNOR2_X1 U813 ( .A(KEYINPUT31), .B(KEYINPUT95), .ZN(n731) );
  NOR2_X1 U814 ( .A1(G2084), .A2(n742), .ZN(n737) );
  NAND2_X1 U815 ( .A1(G8), .A2(n742), .ZN(n807) );
  NOR2_X1 U816 ( .A1(G1966), .A2(n807), .ZN(n734) );
  NOR2_X1 U817 ( .A1(n737), .A2(n734), .ZN(n723) );
  XNOR2_X1 U818 ( .A(KEYINPUT94), .B(n723), .ZN(n724) );
  NAND2_X1 U819 ( .A1(n724), .A2(G8), .ZN(n725) );
  XNOR2_X1 U820 ( .A(KEYINPUT30), .B(n725), .ZN(n726) );
  NOR2_X1 U821 ( .A1(G168), .A2(n726), .ZN(n729) );
  NOR2_X1 U822 ( .A1(G171), .A2(n727), .ZN(n728) );
  NOR2_X1 U823 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U824 ( .A(n731), .B(n730), .ZN(n732) );
  NAND2_X1 U825 ( .A1(n733), .A2(n732), .ZN(n741) );
  INV_X1 U826 ( .A(n734), .ZN(n735) );
  XNOR2_X1 U827 ( .A(n736), .B(KEYINPUT96), .ZN(n739) );
  NAND2_X1 U828 ( .A1(n737), .A2(G8), .ZN(n738) );
  NAND2_X1 U829 ( .A1(n739), .A2(n738), .ZN(n753) );
  AND2_X1 U830 ( .A1(G286), .A2(G8), .ZN(n740) );
  NAND2_X1 U831 ( .A1(n741), .A2(n740), .ZN(n749) );
  INV_X1 U832 ( .A(G8), .ZN(n747) );
  NOR2_X1 U833 ( .A1(G2090), .A2(n742), .ZN(n744) );
  NOR2_X1 U834 ( .A1(G1971), .A2(n807), .ZN(n743) );
  NOR2_X1 U835 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U836 ( .A1(n745), .A2(G303), .ZN(n746) );
  OR2_X1 U837 ( .A1(n747), .A2(n746), .ZN(n748) );
  XOR2_X1 U838 ( .A(KEYINPUT32), .B(KEYINPUT97), .Z(n750) );
  XNOR2_X1 U839 ( .A(n751), .B(n750), .ZN(n752) );
  NAND2_X1 U840 ( .A1(n753), .A2(n752), .ZN(n803) );
  NOR2_X1 U841 ( .A1(G1976), .A2(G288), .ZN(n945) );
  NOR2_X1 U842 ( .A1(G1971), .A2(G303), .ZN(n754) );
  XNOR2_X1 U843 ( .A(KEYINPUT98), .B(n754), .ZN(n755) );
  NOR2_X1 U844 ( .A1(n945), .A2(n755), .ZN(n756) );
  NAND2_X1 U845 ( .A1(n803), .A2(n756), .ZN(n757) );
  NAND2_X1 U846 ( .A1(G1976), .A2(G288), .ZN(n946) );
  NAND2_X1 U847 ( .A1(n757), .A2(n946), .ZN(n758) );
  XNOR2_X1 U848 ( .A(n758), .B(KEYINPUT99), .ZN(n760) );
  AND2_X1 U849 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U850 ( .A1(KEYINPUT33), .A2(n761), .ZN(n764) );
  NAND2_X1 U851 ( .A1(n945), .A2(KEYINPUT33), .ZN(n762) );
  NOR2_X1 U852 ( .A1(n762), .A2(n807), .ZN(n763) );
  XOR2_X1 U853 ( .A(G1981), .B(G305), .Z(n964) );
  NOR2_X1 U854 ( .A1(n766), .A2(n765), .ZN(n767) );
  XOR2_X1 U855 ( .A(n767), .B(KEYINPUT88), .Z(n794) );
  NAND2_X1 U856 ( .A1(n883), .A2(G95), .ZN(n770) );
  BUF_X1 U857 ( .A(n768), .Z(n884) );
  NAND2_X1 U858 ( .A1(G131), .A2(n884), .ZN(n769) );
  NAND2_X1 U859 ( .A1(n770), .A2(n769), .ZN(n774) );
  NAND2_X1 U860 ( .A1(G107), .A2(n887), .ZN(n772) );
  NAND2_X1 U861 ( .A1(G119), .A2(n888), .ZN(n771) );
  NAND2_X1 U862 ( .A1(n772), .A2(n771), .ZN(n773) );
  NOR2_X1 U863 ( .A1(n774), .A2(n773), .ZN(n875) );
  INV_X1 U864 ( .A(G1991), .ZN(n813) );
  NOR2_X1 U865 ( .A1(n875), .A2(n813), .ZN(n783) );
  NAND2_X1 U866 ( .A1(G105), .A2(n883), .ZN(n775) );
  XNOR2_X1 U867 ( .A(n775), .B(KEYINPUT38), .ZN(n777) );
  NAND2_X1 U868 ( .A1(n888), .A2(G129), .ZN(n776) );
  NAND2_X1 U869 ( .A1(n777), .A2(n776), .ZN(n781) );
  NAND2_X1 U870 ( .A1(n887), .A2(G117), .ZN(n779) );
  NAND2_X1 U871 ( .A1(G141), .A2(n884), .ZN(n778) );
  NAND2_X1 U872 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U873 ( .A1(n781), .A2(n780), .ZN(n876) );
  NOR2_X1 U874 ( .A1(n1002), .A2(n876), .ZN(n782) );
  NOR2_X1 U875 ( .A1(n783), .A2(n782), .ZN(n923) );
  NOR2_X1 U876 ( .A1(n794), .A2(n923), .ZN(n816) );
  INV_X1 U877 ( .A(n816), .ZN(n795) );
  NAND2_X1 U878 ( .A1(n883), .A2(G104), .ZN(n785) );
  NAND2_X1 U879 ( .A1(G140), .A2(n884), .ZN(n784) );
  NAND2_X1 U880 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U881 ( .A(KEYINPUT34), .B(n786), .ZN(n792) );
  NAND2_X1 U882 ( .A1(n888), .A2(G128), .ZN(n787) );
  XOR2_X1 U883 ( .A(KEYINPUT89), .B(n787), .Z(n789) );
  NAND2_X1 U884 ( .A1(n887), .A2(G116), .ZN(n788) );
  NAND2_X1 U885 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U886 ( .A(KEYINPUT35), .B(n790), .Z(n791) );
  NOR2_X1 U887 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U888 ( .A(KEYINPUT36), .B(n793), .ZN(n900) );
  XNOR2_X1 U889 ( .A(KEYINPUT37), .B(G2067), .ZN(n812) );
  NOR2_X1 U890 ( .A1(n900), .A2(n812), .ZN(n926) );
  INV_X1 U891 ( .A(n794), .ZN(n824) );
  NAND2_X1 U892 ( .A1(n926), .A2(n824), .ZN(n822) );
  NAND2_X1 U893 ( .A1(n795), .A2(n822), .ZN(n797) );
  XNOR2_X1 U894 ( .A(G1986), .B(G290), .ZN(n950) );
  AND2_X1 U895 ( .A1(n950), .A2(n824), .ZN(n796) );
  NOR2_X1 U896 ( .A1(n797), .A2(n796), .ZN(n800) );
  AND2_X1 U897 ( .A1(n964), .A2(n800), .ZN(n798) );
  NAND2_X1 U898 ( .A1(n799), .A2(n798), .ZN(n829) );
  INV_X1 U899 ( .A(n800), .ZN(n811) );
  NOR2_X1 U900 ( .A1(G2090), .A2(G303), .ZN(n801) );
  NAND2_X1 U901 ( .A1(G8), .A2(n801), .ZN(n802) );
  NAND2_X1 U902 ( .A1(n803), .A2(n802), .ZN(n804) );
  NAND2_X1 U903 ( .A1(n804), .A2(n807), .ZN(n809) );
  NOR2_X1 U904 ( .A1(G1981), .A2(G305), .ZN(n805) );
  XOR2_X1 U905 ( .A(n805), .B(KEYINPUT24), .Z(n806) );
  OR2_X1 U906 ( .A1(n807), .A2(n806), .ZN(n808) );
  AND2_X1 U907 ( .A1(n809), .A2(n808), .ZN(n810) );
  OR2_X1 U908 ( .A1(n811), .A2(n810), .ZN(n827) );
  NAND2_X1 U909 ( .A1(n900), .A2(n812), .ZN(n937) );
  AND2_X1 U910 ( .A1(n813), .A2(n875), .ZN(n919) );
  NOR2_X1 U911 ( .A1(G1986), .A2(G290), .ZN(n814) );
  NOR2_X1 U912 ( .A1(n919), .A2(n814), .ZN(n815) );
  NOR2_X1 U913 ( .A1(n816), .A2(n815), .ZN(n818) );
  AND2_X1 U914 ( .A1(n876), .A2(n1002), .ZN(n817) );
  XNOR2_X1 U915 ( .A(n817), .B(KEYINPUT100), .ZN(n916) );
  NOR2_X1 U916 ( .A1(n818), .A2(n916), .ZN(n820) );
  XOR2_X1 U917 ( .A(KEYINPUT39), .B(KEYINPUT101), .Z(n819) );
  XNOR2_X1 U918 ( .A(n820), .B(n819), .ZN(n821) );
  NAND2_X1 U919 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U920 ( .A1(n937), .A2(n823), .ZN(n825) );
  NAND2_X1 U921 ( .A1(n825), .A2(n824), .ZN(n826) );
  AND2_X1 U922 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U923 ( .A1(n829), .A2(n828), .ZN(n831) );
  XNOR2_X1 U924 ( .A(KEYINPUT40), .B(KEYINPUT102), .ZN(n830) );
  XNOR2_X1 U925 ( .A(n831), .B(n830), .ZN(G329) );
  NAND2_X1 U926 ( .A1(G2106), .A2(n832), .ZN(G217) );
  AND2_X1 U927 ( .A1(G15), .A2(G2), .ZN(n833) );
  NAND2_X1 U928 ( .A1(G661), .A2(n833), .ZN(G259) );
  NAND2_X1 U929 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U930 ( .A1(n835), .A2(n834), .ZN(n836) );
  XOR2_X1 U931 ( .A(KEYINPUT103), .B(n836), .Z(G188) );
  INV_X1 U933 ( .A(G120), .ZN(G236) );
  INV_X1 U934 ( .A(G96), .ZN(G221) );
  INV_X1 U935 ( .A(G69), .ZN(G235) );
  NOR2_X1 U936 ( .A1(n838), .A2(n837), .ZN(G325) );
  INV_X1 U937 ( .A(G325), .ZN(G261) );
  INV_X1 U938 ( .A(n839), .ZN(G319) );
  XOR2_X1 U939 ( .A(G2096), .B(KEYINPUT43), .Z(n841) );
  XNOR2_X1 U940 ( .A(G2072), .B(G2678), .ZN(n840) );
  XNOR2_X1 U941 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U942 ( .A(n842), .B(KEYINPUT42), .Z(n844) );
  XNOR2_X1 U943 ( .A(G2067), .B(G2090), .ZN(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U945 ( .A(KEYINPUT104), .B(G2100), .Z(n846) );
  XNOR2_X1 U946 ( .A(G2084), .B(G2078), .ZN(n845) );
  XNOR2_X1 U947 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(G227) );
  XOR2_X1 U949 ( .A(G1956), .B(G1961), .Z(n850) );
  XNOR2_X1 U950 ( .A(G1986), .B(G1966), .ZN(n849) );
  XNOR2_X1 U951 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U952 ( .A(G1976), .B(G1971), .Z(n852) );
  XNOR2_X1 U953 ( .A(G1996), .B(G1991), .ZN(n851) );
  XNOR2_X1 U954 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U955 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U956 ( .A(G2474), .B(KEYINPUT41), .ZN(n855) );
  XNOR2_X1 U957 ( .A(n856), .B(n855), .ZN(n858) );
  XOR2_X1 U958 ( .A(G1981), .B(KEYINPUT105), .Z(n857) );
  XNOR2_X1 U959 ( .A(n858), .B(n857), .ZN(G229) );
  NAND2_X1 U960 ( .A1(n883), .A2(G100), .ZN(n860) );
  NAND2_X1 U961 ( .A1(G136), .A2(n884), .ZN(n859) );
  NAND2_X1 U962 ( .A1(n860), .A2(n859), .ZN(n865) );
  NAND2_X1 U963 ( .A1(G124), .A2(n888), .ZN(n861) );
  XNOR2_X1 U964 ( .A(n861), .B(KEYINPUT44), .ZN(n863) );
  NAND2_X1 U965 ( .A1(n887), .A2(G112), .ZN(n862) );
  NAND2_X1 U966 ( .A1(n863), .A2(n862), .ZN(n864) );
  NOR2_X1 U967 ( .A1(n865), .A2(n864), .ZN(G162) );
  NAND2_X1 U968 ( .A1(n883), .A2(G106), .ZN(n866) );
  XOR2_X1 U969 ( .A(KEYINPUT107), .B(n866), .Z(n868) );
  NAND2_X1 U970 ( .A1(G142), .A2(n884), .ZN(n867) );
  NAND2_X1 U971 ( .A1(n868), .A2(n867), .ZN(n869) );
  XNOR2_X1 U972 ( .A(n869), .B(KEYINPUT45), .ZN(n871) );
  NAND2_X1 U973 ( .A1(G130), .A2(n888), .ZN(n870) );
  NAND2_X1 U974 ( .A1(n871), .A2(n870), .ZN(n874) );
  NAND2_X1 U975 ( .A1(n887), .A2(G118), .ZN(n872) );
  XOR2_X1 U976 ( .A(KEYINPUT106), .B(n872), .Z(n873) );
  NOR2_X1 U977 ( .A1(n874), .A2(n873), .ZN(n898) );
  XOR2_X1 U978 ( .A(G162), .B(n875), .Z(n878) );
  XNOR2_X1 U979 ( .A(G160), .B(n876), .ZN(n877) );
  XNOR2_X1 U980 ( .A(n878), .B(n877), .ZN(n882) );
  XOR2_X1 U981 ( .A(KEYINPUT110), .B(KEYINPUT108), .Z(n880) );
  XNOR2_X1 U982 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n879) );
  XNOR2_X1 U983 ( .A(n880), .B(n879), .ZN(n881) );
  XOR2_X1 U984 ( .A(n882), .B(n881), .Z(n896) );
  NAND2_X1 U985 ( .A1(n883), .A2(G103), .ZN(n886) );
  NAND2_X1 U986 ( .A1(G139), .A2(n884), .ZN(n885) );
  NAND2_X1 U987 ( .A1(n886), .A2(n885), .ZN(n894) );
  NAND2_X1 U988 ( .A1(G115), .A2(n887), .ZN(n890) );
  NAND2_X1 U989 ( .A1(G127), .A2(n888), .ZN(n889) );
  NAND2_X1 U990 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U991 ( .A(KEYINPUT109), .B(n891), .ZN(n892) );
  XNOR2_X1 U992 ( .A(KEYINPUT47), .B(n892), .ZN(n893) );
  NOR2_X1 U993 ( .A1(n894), .A2(n893), .ZN(n930) );
  XNOR2_X1 U994 ( .A(G164), .B(n930), .ZN(n895) );
  XNOR2_X1 U995 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U996 ( .A(n898), .B(n897), .Z(n899) );
  XNOR2_X1 U997 ( .A(n920), .B(n899), .ZN(n901) );
  XOR2_X1 U998 ( .A(n901), .B(n900), .Z(n902) );
  NOR2_X1 U999 ( .A1(G37), .A2(n902), .ZN(G395) );
  XNOR2_X1 U1000 ( .A(n954), .B(n903), .ZN(n905) );
  XNOR2_X1 U1001 ( .A(G171), .B(n959), .ZN(n904) );
  XNOR2_X1 U1002 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1003 ( .A(G286), .B(n906), .Z(n907) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n907), .ZN(n908) );
  XOR2_X1 U1005 ( .A(KEYINPUT111), .B(n908), .Z(G397) );
  NOR2_X1 U1006 ( .A1(G227), .A2(G229), .ZN(n909) );
  XOR2_X1 U1007 ( .A(KEYINPUT49), .B(n909), .Z(n910) );
  NAND2_X1 U1008 ( .A1(G319), .A2(n910), .ZN(n911) );
  NOR2_X1 U1009 ( .A1(G401), .A2(n911), .ZN(n912) );
  XNOR2_X1 U1010 ( .A(KEYINPUT112), .B(n912), .ZN(n914) );
  NOR2_X1 U1011 ( .A1(G395), .A2(G397), .ZN(n913) );
  NAND2_X1 U1012 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1015 ( .A(G2090), .B(G162), .Z(n915) );
  NOR2_X1 U1016 ( .A1(n916), .A2(n915), .ZN(n917) );
  XOR2_X1 U1017 ( .A(KEYINPUT51), .B(n917), .Z(n929) );
  XOR2_X1 U1018 ( .A(G160), .B(G2084), .Z(n918) );
  NOR2_X1 U1019 ( .A1(n919), .A2(n918), .ZN(n921) );
  NAND2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(KEYINPUT113), .B(n922), .ZN(n924) );
  NAND2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n925) );
  NOR2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1024 ( .A(n927), .B(KEYINPUT114), .ZN(n928) );
  NAND2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n935) );
  XOR2_X1 U1026 ( .A(G2072), .B(n930), .Z(n932) );
  XOR2_X1 U1027 ( .A(G164), .B(G2078), .Z(n931) );
  NOR2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1029 ( .A(KEYINPUT50), .B(n933), .Z(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1032 ( .A(n938), .B(KEYINPUT52), .ZN(n939) );
  XNOR2_X1 U1033 ( .A(KEYINPUT115), .B(n939), .ZN(n941) );
  INV_X1 U1034 ( .A(KEYINPUT55), .ZN(n940) );
  NAND2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1036 ( .A1(n942), .A2(G29), .ZN(n1027) );
  XNOR2_X1 U1037 ( .A(G16), .B(KEYINPUT56), .ZN(n970) );
  XNOR2_X1 U1038 ( .A(G299), .B(G1956), .ZN(n944) );
  XNOR2_X1 U1039 ( .A(G303), .B(G1971), .ZN(n943) );
  NOR2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n952) );
  XNOR2_X1 U1041 ( .A(n945), .B(KEYINPUT119), .ZN(n947) );
  NAND2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1043 ( .A(n948), .B(KEYINPUT120), .ZN(n949) );
  NOR2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1045 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1046 ( .A(KEYINPUT121), .B(n953), .ZN(n958) );
  XOR2_X1 U1047 ( .A(G171), .B(G1961), .Z(n956) );
  XNOR2_X1 U1048 ( .A(n954), .B(G1341), .ZN(n955) );
  NOR2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1050 ( .A1(n958), .A2(n957), .ZN(n962) );
  XOR2_X1 U1051 ( .A(G1348), .B(n959), .Z(n960) );
  XNOR2_X1 U1052 ( .A(KEYINPUT118), .B(n960), .ZN(n961) );
  NOR2_X1 U1053 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1054 ( .A(KEYINPUT122), .B(n963), .ZN(n968) );
  XNOR2_X1 U1055 ( .A(G1966), .B(G168), .ZN(n965) );
  NAND2_X1 U1056 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1057 ( .A(KEYINPUT57), .B(n966), .ZN(n967) );
  NAND2_X1 U1058 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1059 ( .A1(n970), .A2(n969), .ZN(n999) );
  INV_X1 U1060 ( .A(G16), .ZN(n997) );
  XNOR2_X1 U1061 ( .A(G1348), .B(KEYINPUT59), .ZN(n971) );
  XNOR2_X1 U1062 ( .A(n971), .B(G4), .ZN(n975) );
  XNOR2_X1 U1063 ( .A(G1956), .B(G20), .ZN(n973) );
  XNOR2_X1 U1064 ( .A(G19), .B(G1341), .ZN(n972) );
  NOR2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n978) );
  XOR2_X1 U1067 ( .A(KEYINPUT123), .B(G1981), .Z(n976) );
  XNOR2_X1 U1068 ( .A(G6), .B(n976), .ZN(n977) );
  NOR2_X1 U1069 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1070 ( .A(KEYINPUT60), .B(n979), .Z(n981) );
  XNOR2_X1 U1071 ( .A(G1966), .B(G21), .ZN(n980) );
  NOR2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(KEYINPUT124), .B(n982), .ZN(n985) );
  XNOR2_X1 U1074 ( .A(n983), .B(G5), .ZN(n984) );
  NAND2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n993) );
  XNOR2_X1 U1076 ( .A(G1986), .B(G24), .ZN(n987) );
  XNOR2_X1 U1077 ( .A(G23), .B(G1976), .ZN(n986) );
  NOR2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n990) );
  XNOR2_X1 U1079 ( .A(G1971), .B(KEYINPUT125), .ZN(n988) );
  XNOR2_X1 U1080 ( .A(n988), .B(G22), .ZN(n989) );
  NAND2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1082 ( .A(KEYINPUT58), .B(n991), .ZN(n992) );
  NOR2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(n994), .B(KEYINPUT61), .ZN(n995) );
  XNOR2_X1 U1085 ( .A(n995), .B(KEYINPUT126), .ZN(n996) );
  NAND2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1024) );
  XNOR2_X1 U1088 ( .A(G1991), .B(G25), .ZN(n1001) );
  XNOR2_X1 U1089 ( .A(G33), .B(G2072), .ZN(n1000) );
  NOR2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1008) );
  XNOR2_X1 U1091 ( .A(G32), .B(n1002), .ZN(n1003) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(G28), .ZN(n1006) );
  XNOR2_X1 U1093 ( .A(KEYINPUT116), .B(G2067), .ZN(n1004) );
  XNOR2_X1 U1094 ( .A(G26), .B(n1004), .ZN(n1005) );
  NOR2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1011) );
  XOR2_X1 U1097 ( .A(G27), .B(n1009), .Z(n1010) );
  NOR2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1099 ( .A(KEYINPUT53), .B(n1012), .Z(n1015) );
  XOR2_X1 U1100 ( .A(KEYINPUT54), .B(G34), .Z(n1013) );
  XNOR2_X1 U1101 ( .A(G2084), .B(n1013), .ZN(n1014) );
  NAND2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1017) );
  XNOR2_X1 U1103 ( .A(G35), .B(G2090), .ZN(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1105 ( .A(KEYINPUT55), .B(n1018), .ZN(n1020) );
  INV_X1 U1106 ( .A(G29), .ZN(n1019) );
  NAND2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1108 ( .A1(n1021), .A2(G11), .ZN(n1022) );
  XOR2_X1 U1109 ( .A(KEYINPUT117), .B(n1022), .Z(n1023) );
  NOR2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1111 ( .A(KEYINPUT127), .B(n1025), .Z(n1026) );
  NAND2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XOR2_X1 U1113 ( .A(KEYINPUT62), .B(n1028), .Z(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

