//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 0 1 0 1 1 0 0 0 1 0 1 1 1 1 1 1 1 0 1 1 1 0 0 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NOR3_X1   g0007(.A1(new_n207), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0009(.A(G97), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  INV_X1    g0011(.A(G107), .ZN(new_n212));
  INV_X1    g0012(.A(G264), .ZN(new_n213));
  OAI22_X1  g0013(.A1(new_n210), .A2(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G77), .A2(G244), .ZN(new_n215));
  INV_X1    g0015(.A(G50), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  INV_X1    g0017(.A(G232), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n202), .C2(new_n218), .ZN(new_n219));
  AOI211_X1 g0019(.A(new_n214), .B(new_n219), .C1(G87), .C2(G250), .ZN(new_n220));
  XOR2_X1   g0020(.A(KEYINPUT65), .B(G238), .Z(new_n221));
  INV_X1    g0021(.A(G116), .ZN(new_n222));
  INV_X1    g0022(.A(G270), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n220), .B1(new_n203), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G20), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT1), .Z(new_n227));
  NOR2_X1   g0027(.A1(new_n225), .A2(G13), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G250), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(new_n211), .B2(new_n213), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n206), .A2(new_n216), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  INV_X1    g0032(.A(G20), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  AOI22_X1  g0034(.A1(new_n230), .A2(KEYINPUT0), .B1(new_n231), .B2(new_n234), .ZN(new_n235));
  OAI211_X1 g0035(.A(new_n227), .B(new_n235), .C1(KEYINPUT0), .C2(new_n230), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G226), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G264), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n223), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(G107), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G77), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n212), .A2(KEYINPUT6), .A3(G97), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n210), .A2(new_n212), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G97), .A2(G107), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n256), .B1(new_n259), .B2(KEYINPUT6), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G20), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  OAI21_X1  g0062(.A(KEYINPUT78), .B1(new_n262), .B2(KEYINPUT3), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT78), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT3), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n264), .A2(new_n265), .A3(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n263), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(KEYINPUT7), .A3(new_n233), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT7), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT3), .B(G33), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n270), .B1(new_n271), .B2(G20), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n255), .B(new_n261), .C1(new_n273), .C2(new_n212), .ZN(new_n274));
  NAND3_X1  g0074(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n232), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G13), .ZN(new_n278));
  NOR3_X1   g0078(.A1(new_n278), .A2(new_n233), .A3(G1), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(G97), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n276), .ZN(new_n283));
  INV_X1    g0083(.A(G1), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G33), .ZN(new_n285));
  AND3_X1   g0085(.A1(new_n280), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G97), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n277), .A2(new_n282), .A3(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT81), .ZN(new_n289));
  INV_X1    g0089(.A(G41), .ZN(new_n290));
  OAI211_X1 g0090(.A(G1), .B(G13), .C1(new_n262), .C2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n265), .A2(G33), .ZN(new_n292));
  INV_X1    g0092(.A(G1698), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n267), .A2(new_n292), .A3(G244), .A4(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT80), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT4), .ZN(new_n296));
  AND3_X1   g0096(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n296), .B1(new_n294), .B2(new_n295), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n267), .A2(new_n292), .A3(G250), .A4(G1698), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G33), .A2(G283), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n291), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n291), .A2(G274), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n290), .A2(KEYINPUT5), .ZN(new_n305));
  INV_X1    g0105(.A(G45), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n306), .A2(G1), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n290), .A2(KEYINPUT67), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT67), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G41), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT5), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n308), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n304), .A2(new_n305), .A3(new_n307), .A4(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n312), .A2(new_n305), .A3(new_n307), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n314), .A2(G257), .A3(new_n291), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n289), .B1(new_n303), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n294), .A2(new_n295), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT4), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(new_n302), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n232), .B1(G33), .B2(G41), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n316), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n323), .A2(new_n324), .A3(KEYINPUT81), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n317), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n288), .B1(new_n326), .B2(G190), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n323), .A2(new_n324), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G200), .ZN(new_n329));
  INV_X1    g0129(.A(G179), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n323), .A2(new_n324), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT82), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT82), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n323), .A2(new_n324), .A3(new_n333), .A4(new_n330), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n281), .B1(new_n274), .B2(new_n276), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n332), .A2(new_n334), .B1(new_n335), .B2(new_n287), .ZN(new_n336));
  INV_X1    g0136(.A(G169), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n317), .A2(new_n337), .A3(new_n325), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n327), .A2(new_n329), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT71), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT8), .B(G58), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n233), .A2(G33), .ZN(new_n342));
  INV_X1    g0142(.A(G150), .ZN(new_n343));
  INV_X1    g0143(.A(new_n254), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n341), .A2(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT69), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n233), .B1(new_n206), .B2(new_n216), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n276), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n279), .A2(new_n216), .ZN(new_n349));
  AND2_X1   g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n283), .B1(G1), .B2(new_n233), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(G50), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n350), .A2(KEYINPUT9), .A3(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(KEYINPUT9), .B1(new_n350), .B2(new_n353), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n340), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n350), .A2(new_n353), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT9), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n360), .A2(KEYINPUT71), .A3(new_n354), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n271), .A2(G223), .A3(G1698), .ZN(new_n362));
  INV_X1    g0162(.A(G77), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n271), .A2(new_n293), .ZN(new_n364));
  INV_X1    g0164(.A(G222), .ZN(new_n365));
  OAI221_X1 g0165(.A(new_n362), .B1(new_n363), .B2(new_n271), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n322), .ZN(new_n367));
  AOI21_X1  g0167(.A(G45), .B1(new_n308), .B2(new_n310), .ZN(new_n368));
  OAI21_X1  g0168(.A(KEYINPUT68), .B1(new_n368), .B2(G1), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT68), .ZN(new_n370));
  XNOR2_X1  g0170(.A(KEYINPUT67), .B(G41), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n370), .B(new_n284), .C1(new_n371), .C2(G45), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n369), .A2(new_n304), .A3(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n284), .B1(G41), .B2(G45), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n291), .A2(new_n374), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n367), .B(new_n373), .C1(new_n217), .C2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G190), .ZN(new_n377));
  OR2_X1    g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT73), .ZN(new_n379));
  XNOR2_X1  g0179(.A(new_n378), .B(new_n379), .ZN(new_n380));
  AND3_X1   g0180(.A1(new_n376), .A2(KEYINPUT72), .A3(G200), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT72), .B1(new_n376), .B2(G200), .ZN(new_n382));
  NOR3_X1   g0182(.A1(new_n381), .A2(new_n382), .A3(KEYINPUT10), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n357), .A2(new_n361), .A3(new_n380), .A4(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n376), .A2(G200), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n360), .A2(new_n385), .A3(new_n354), .ZN(new_n386));
  XNOR2_X1  g0186(.A(new_n378), .B(KEYINPUT73), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT10), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n384), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n376), .A2(new_n337), .ZN(new_n390));
  OR2_X1    g0190(.A1(new_n376), .A2(G179), .ZN(new_n391));
  AND3_X1   g0191(.A1(new_n358), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT74), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n373), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n369), .A2(KEYINPUT74), .A3(new_n304), .A4(new_n372), .ZN(new_n397));
  XOR2_X1   g0197(.A(new_n375), .B(KEYINPUT75), .Z(new_n398));
  AOI22_X1  g0198(.A1(new_n396), .A2(new_n397), .B1(new_n398), .B2(G238), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT13), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n271), .A2(G232), .A3(G1698), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G33), .A2(G97), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n401), .B(new_n402), .C1(new_n364), .C2(new_n217), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n322), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n399), .A2(new_n400), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n400), .B1(new_n399), .B2(new_n404), .ZN(new_n407));
  OAI21_X1  g0207(.A(G169), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT14), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n399), .A2(new_n404), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT13), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n405), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT14), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(new_n413), .A3(G169), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n411), .A2(G179), .A3(new_n405), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n409), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n203), .A2(G20), .ZN(new_n417));
  OAI221_X1 g0217(.A(new_n417), .B1(new_n342), .B2(new_n363), .C1(new_n344), .C2(new_n216), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n418), .A2(KEYINPUT11), .A3(new_n276), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n203), .B2(new_n351), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n279), .A2(new_n203), .ZN(new_n421));
  XOR2_X1   g0221(.A(new_n421), .B(KEYINPUT12), .Z(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT11), .B1(new_n418), .B2(new_n276), .ZN(new_n423));
  NOR3_X1   g0223(.A1(new_n420), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n416), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n412), .A2(G200), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n411), .A2(G190), .A3(new_n405), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n427), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G20), .A2(G77), .ZN(new_n430));
  XOR2_X1   g0230(.A(KEYINPUT15), .B(G87), .Z(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  OAI221_X1 g0232(.A(new_n430), .B1(new_n344), .B2(new_n341), .C1(new_n432), .C2(new_n342), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n433), .A2(new_n276), .B1(new_n363), .B2(new_n279), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n363), .B2(new_n351), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n271), .A2(G232), .A3(new_n293), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n271), .A2(G1698), .ZN(new_n437));
  OAI221_X1 g0237(.A(new_n436), .B1(new_n212), .B2(new_n271), .C1(new_n437), .C2(new_n221), .ZN(new_n438));
  XOR2_X1   g0238(.A(new_n438), .B(KEYINPUT70), .Z(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n322), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n291), .A2(G244), .A3(new_n374), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n373), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n435), .B1(new_n443), .B2(G200), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(new_n377), .B2(new_n443), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n426), .A2(new_n429), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n443), .A2(new_n337), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n440), .A2(new_n330), .A3(new_n442), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n447), .A2(new_n435), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n271), .A2(G223), .A3(new_n293), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G33), .A2(G87), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n451), .B(new_n452), .C1(new_n437), .C2(new_n217), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n322), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT79), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n455), .B1(new_n375), .B2(new_n218), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n291), .A2(KEYINPUT79), .A3(G232), .A4(new_n374), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n454), .A2(new_n458), .A3(new_n373), .ZN(new_n459));
  OR2_X1    g0259(.A1(new_n459), .A2(new_n377), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(G200), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT16), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n203), .B1(new_n269), .B2(new_n272), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n204), .B(new_n205), .C1(new_n202), .C2(new_n203), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G20), .ZN(new_n465));
  INV_X1    g0265(.A(G159), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT77), .B1(new_n344), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT77), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n254), .A2(new_n468), .A3(G159), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n462), .B1(new_n463), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(KEYINPUT7), .A2(G20), .ZN(new_n473));
  AND3_X1   g0273(.A1(new_n267), .A2(new_n292), .A3(KEYINPUT76), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT76), .B1(new_n267), .B2(new_n292), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(KEYINPUT7), .B1(new_n271), .B2(G20), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n476), .A2(G68), .A3(new_n477), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n464), .A2(G20), .B1(new_n467), .B2(new_n469), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n478), .A2(KEYINPUT16), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n472), .A2(new_n480), .A3(new_n276), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n280), .A2(new_n341), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(new_n352), .B2(new_n341), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n460), .A2(new_n461), .A3(new_n481), .A4(new_n483), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n484), .A2(KEYINPUT17), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n484), .A2(KEYINPUT17), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n481), .A2(new_n483), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n459), .A2(G169), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n454), .A2(new_n458), .A3(new_n373), .A4(G179), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT18), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(KEYINPUT18), .B1(new_n487), .B2(new_n490), .ZN(new_n494));
  OAI22_X1  g0294(.A1(new_n485), .A2(new_n486), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OR2_X1    g0295(.A1(new_n450), .A2(new_n495), .ZN(new_n496));
  NOR3_X1   g0296(.A1(new_n394), .A2(new_n446), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n271), .A2(new_n233), .A3(G68), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT19), .ZN(new_n499));
  INV_X1    g0299(.A(G87), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n258), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n402), .A2(new_n233), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NOR3_X1   g0303(.A1(new_n402), .A2(KEYINPUT19), .A3(G20), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n498), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT83), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT83), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n498), .B(new_n507), .C1(new_n503), .C2(new_n504), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n506), .A2(new_n276), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n286), .A2(new_n431), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n432), .A2(new_n279), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n271), .A2(G238), .A3(new_n293), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n271), .A2(G244), .A3(G1698), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G116), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n322), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n307), .A2(G274), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n291), .B(G250), .C1(G1), .C2(new_n306), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n337), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n517), .A2(new_n330), .A3(new_n518), .A4(new_n519), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n512), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n517), .A2(G190), .A3(new_n518), .A4(new_n519), .ZN(new_n524));
  INV_X1    g0324(.A(new_n520), .ZN(new_n525));
  INV_X1    g0325(.A(G200), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n286), .A2(G87), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n509), .A2(new_n511), .A3(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n523), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n515), .A2(G20), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n267), .A2(new_n292), .A3(new_n233), .A4(G87), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(KEYINPUT22), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT22), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n271), .A2(new_n534), .A3(new_n233), .A4(G87), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n531), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT24), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n233), .A2(G107), .ZN(new_n538));
  XNOR2_X1  g0338(.A(new_n538), .B(KEYINPUT23), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n537), .B1(new_n536), .B2(new_n539), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n276), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n286), .A2(G107), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n279), .A2(new_n212), .ZN(new_n544));
  XOR2_X1   g0344(.A(new_n544), .B(KEYINPUT25), .Z(new_n545));
  NAND3_X1  g0345(.A1(new_n542), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n267), .A2(new_n292), .A3(G257), .A4(G1698), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n267), .A2(new_n292), .A3(G250), .A4(new_n293), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G33), .A2(G294), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(KEYINPUT84), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT84), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n547), .A2(new_n548), .A3(new_n552), .A4(new_n549), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n551), .A2(new_n322), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n314), .A2(G264), .A3(new_n291), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n554), .A2(new_n555), .A3(new_n313), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n557), .A2(new_n526), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n546), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n557), .A2(G190), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n530), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n556), .A2(new_n337), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n557), .A2(new_n330), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n546), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT21), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n267), .A2(new_n292), .A3(G257), .A4(new_n293), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n267), .A2(new_n292), .A3(G264), .A4(G1698), .ZN(new_n567));
  INV_X1    g0367(.A(G303), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n566), .B(new_n567), .C1(new_n568), .C2(new_n271), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n322), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n314), .A2(G270), .A3(new_n291), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n570), .A2(new_n313), .A3(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n280), .A2(G116), .A3(new_n283), .A4(new_n285), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n279), .A2(new_n222), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n275), .A2(new_n232), .B1(G20), .B2(new_n222), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n301), .B(new_n233), .C1(G33), .C2(new_n210), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n576), .A2(KEYINPUT20), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT20), .B1(new_n576), .B2(new_n577), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n574), .B(new_n575), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(G169), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n565), .B1(new_n573), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n573), .A2(G179), .A3(new_n580), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n572), .A2(KEYINPUT21), .A3(G169), .A4(new_n580), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n580), .B1(new_n572), .B2(G200), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(new_n377), .B2(new_n572), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n564), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  AND4_X1   g0389(.A1(new_n339), .A2(new_n497), .A3(new_n561), .A4(new_n589), .ZN(G372));
  NAND2_X1  g0390(.A1(new_n426), .A2(new_n449), .ZN(new_n591));
  OR2_X1    g0391(.A1(new_n485), .A2(new_n486), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(new_n429), .A3(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT86), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n487), .A2(new_n490), .A3(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n594), .B1(new_n487), .B2(new_n490), .ZN(new_n597));
  NOR3_X1   g0397(.A1(new_n596), .A2(new_n597), .A3(KEYINPUT87), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT87), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n491), .A2(KEYINPUT86), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n599), .B1(new_n600), .B2(new_n595), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n492), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(KEYINPUT87), .B1(new_n596), .B2(new_n597), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n600), .A2(new_n599), .A3(new_n595), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n603), .A2(new_n604), .A3(KEYINPUT18), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n593), .A2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n389), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n393), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n339), .A2(new_n561), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(KEYINPUT85), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n564), .A2(new_n586), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT85), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n339), .A2(new_n613), .A3(new_n561), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n611), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n523), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n336), .A2(new_n338), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n530), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n618), .A2(KEYINPUT26), .A3(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT26), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n617), .B2(new_n530), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n616), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n615), .A2(new_n623), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n497), .A2(new_n624), .ZN(new_n625));
  OR2_X1    g0425(.A1(new_n609), .A2(new_n625), .ZN(G369));
  NOR2_X1   g0426(.A1(new_n278), .A2(G20), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n284), .ZN(new_n628));
  OR2_X1    g0428(.A1(new_n628), .A2(KEYINPUT27), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(KEYINPUT27), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n629), .A2(G213), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(G343), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n633), .A2(new_n580), .ZN(new_n634));
  XNOR2_X1  g0434(.A(new_n585), .B(new_n634), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n635), .A2(new_n588), .ZN(new_n636));
  XNOR2_X1  g0436(.A(new_n636), .B(KEYINPUT88), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(G330), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT89), .ZN(new_n639));
  XNOR2_X1  g0439(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n564), .A2(new_n633), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n559), .A2(new_n560), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n546), .A2(new_n633), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n641), .B1(new_n644), .B2(new_n564), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n640), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n586), .A2(new_n633), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(new_n564), .B2(new_n633), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n651), .B(KEYINPUT90), .ZN(G399));
  NOR2_X1   g0452(.A1(new_n501), .A2(G116), .ZN(new_n653));
  XOR2_X1   g0453(.A(new_n653), .B(KEYINPUT91), .Z(new_n654));
  INV_X1    g0454(.A(new_n228), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(new_n371), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n654), .A2(new_n284), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n657), .B1(new_n231), .B2(new_n656), .ZN(new_n658));
  XOR2_X1   g0458(.A(new_n658), .B(KEYINPUT28), .Z(new_n659));
  AOI21_X1  g0459(.A(new_n633), .B1(new_n615), .B2(new_n623), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT29), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n612), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n623), .B1(new_n610), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n632), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(KEYINPUT29), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(G330), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n554), .A2(new_n555), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n570), .A2(G179), .A3(new_n313), .A4(new_n571), .ZN(new_n670));
  NOR3_X1   g0470(.A1(new_n669), .A2(new_n520), .A3(new_n670), .ZN(new_n671));
  NOR3_X1   g0471(.A1(new_n303), .A2(new_n289), .A3(new_n316), .ZN(new_n672));
  AOI21_X1  g0472(.A(KEYINPUT81), .B1(new_n323), .B2(new_n324), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT30), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n525), .A2(new_n573), .A3(G179), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n677), .A2(new_n328), .A3(new_n556), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n326), .A2(KEYINPUT30), .A3(new_n671), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n676), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n633), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(KEYINPUT31), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT31), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n680), .A2(new_n683), .A3(new_n633), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n339), .A2(new_n589), .A3(new_n561), .A4(new_n632), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n668), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n667), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n659), .B1(new_n688), .B2(G1), .ZN(G364));
  XNOR2_X1  g0489(.A(new_n638), .B(KEYINPUT89), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n284), .B1(new_n627), .B2(G45), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n656), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g0493(.A(new_n693), .B(KEYINPUT92), .Z(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n690), .B(new_n695), .C1(G330), .C2(new_n637), .ZN(new_n696));
  NOR2_X1   g0496(.A1(G179), .A2(G200), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G190), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G20), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(G294), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(new_n377), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n271), .B1(new_n704), .B2(G326), .ZN(new_n705));
  INV_X1    g0505(.A(G311), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n330), .A2(G200), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n233), .A2(G190), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n705), .B1(new_n706), .B2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n703), .A2(G190), .ZN(new_n711));
  XNOR2_X1  g0511(.A(KEYINPUT33), .B(G317), .ZN(new_n712));
  AOI211_X1 g0512(.A(new_n702), .B(new_n710), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n233), .A2(new_n377), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n526), .A2(G179), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G303), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n708), .A2(new_n715), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT96), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G283), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n714), .A2(new_n707), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n708), .A2(new_n697), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  AOI22_X1  g0525(.A1(G322), .A2(new_n723), .B1(new_n725), .B2(G329), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n713), .A2(new_n718), .A3(new_n721), .A4(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n271), .B1(new_n716), .B2(new_n500), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n725), .A2(G159), .ZN(new_n729));
  INV_X1    g0529(.A(new_n704), .ZN(new_n730));
  OAI22_X1  g0530(.A1(new_n729), .A2(KEYINPUT32), .B1(new_n216), .B2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n709), .ZN(new_n732));
  AOI211_X1 g0532(.A(new_n728), .B(new_n731), .C1(G77), .C2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n699), .A2(G97), .ZN(new_n734));
  AOI22_X1  g0534(.A1(new_n729), .A2(KEYINPUT32), .B1(G68), .B2(new_n711), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n720), .A2(G107), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n733), .A2(new_n734), .A3(new_n735), .A4(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n722), .A2(new_n202), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n727), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n232), .B1(G20), .B2(new_n337), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n474), .ZN(new_n742));
  INV_X1    g0542(.A(new_n475), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(new_n228), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n745), .B(KEYINPUT95), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n249), .A2(G45), .ZN(new_n747));
  INV_X1    g0547(.A(new_n231), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n746), .B(new_n747), .C1(G45), .C2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n271), .A2(new_n228), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT93), .ZN(new_n751));
  XOR2_X1   g0551(.A(G355), .B(KEYINPUT94), .Z(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n749), .B(new_n753), .C1(G116), .C2(new_n228), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G13), .A2(G33), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(G20), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n740), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n695), .B1(new_n754), .B2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n757), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n741), .B(new_n759), .C1(new_n636), .C2(new_n760), .ZN(new_n761));
  AND2_X1   g0561(.A1(new_n696), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(G396));
  AND2_X1   g0563(.A1(new_n720), .A2(G68), .ZN(new_n764));
  INV_X1    g0564(.A(new_n744), .ZN(new_n765));
  OAI221_X1 g0565(.A(new_n765), .B1(new_n216), .B2(new_n716), .C1(new_n202), .C2(new_n700), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n732), .A2(G159), .B1(G137), .B2(new_n704), .ZN(new_n767));
  INV_X1    g0567(.A(G143), .ZN(new_n768));
  INV_X1    g0568(.A(new_n711), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n767), .B1(new_n768), .B2(new_n722), .C1(new_n343), .C2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT34), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n764), .B(new_n766), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G132), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n772), .B1(new_n771), .B2(new_n770), .C1(new_n773), .C2(new_n724), .ZN(new_n774));
  INV_X1    g0574(.A(G283), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n775), .A2(new_n769), .B1(new_n730), .B2(new_n568), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n267), .A2(new_n292), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n734), .A2(new_n777), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n776), .B(new_n778), .C1(G294), .C2(new_n723), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n716), .A2(new_n212), .B1(new_n724), .B2(new_n706), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n780), .B1(new_n720), .B2(G87), .ZN(new_n781));
  OAI211_X1 g0581(.A(new_n779), .B(new_n781), .C1(new_n222), .C2(new_n709), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n774), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n695), .B1(new_n783), .B2(new_n740), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n740), .A2(new_n755), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n435), .A2(new_n633), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n445), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(new_n449), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n450), .A2(new_n632), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n784), .B1(G77), .B2(new_n786), .C1(new_n792), .C2(new_n756), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n660), .B(new_n791), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n687), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n694), .B1(new_n795), .B2(KEYINPUT97), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(KEYINPUT97), .B2(new_n795), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n794), .A2(new_n687), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n793), .B1(new_n797), .B2(new_n798), .ZN(G384));
  XNOR2_X1  g0599(.A(new_n790), .B(KEYINPUT99), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n800), .B1(new_n660), .B2(new_n792), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n425), .A2(new_n633), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n426), .A2(new_n429), .A3(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n429), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n425), .B(new_n633), .C1(new_n804), .C2(new_n416), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n801), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n480), .A2(new_n276), .ZN(new_n809));
  AOI21_X1  g0609(.A(KEYINPUT16), .B1(new_n478), .B2(new_n479), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n483), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n495), .A2(new_n631), .A3(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n631), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n488), .A2(new_n489), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(new_n487), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT37), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n815), .A2(new_n484), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n814), .A2(new_n811), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n818), .A2(new_n484), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n817), .B1(new_n819), .B2(new_n816), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n812), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT38), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n812), .A2(KEYINPUT38), .A3(new_n820), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n808), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n487), .A2(new_n631), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(new_n606), .B2(new_n592), .ZN(new_n828));
  INV_X1    g0628(.A(new_n817), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n600), .A2(new_n484), .A3(new_n595), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(KEYINPUT100), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT100), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n600), .A2(new_n832), .A3(new_n484), .A4(new_n595), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n831), .A2(new_n833), .A3(new_n827), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n829), .B1(new_n834), .B2(KEYINPUT37), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n822), .B1(new_n828), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n824), .A2(KEYINPUT101), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT101), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n812), .A2(new_n838), .A3(KEYINPUT38), .A4(new_n820), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n841), .A2(KEYINPUT39), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(KEYINPUT39), .B2(new_n825), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n416), .A2(new_n425), .A3(new_n632), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n826), .B1(new_n606), .B2(new_n631), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n609), .B1(new_n497), .B2(new_n667), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n845), .B(new_n846), .ZN(new_n847));
  AND3_X1   g0647(.A1(new_n680), .A2(new_n683), .A3(new_n633), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n683), .B1(new_n680), .B2(new_n633), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n686), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT102), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n686), .B(KEYINPUT102), .C1(new_n848), .C2(new_n849), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n791), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT40), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n823), .A2(new_n855), .A3(new_n824), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT103), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(KEYINPUT40), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n854), .A2(new_n806), .A3(new_n856), .A4(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT102), .B1(new_n685), .B2(new_n686), .ZN(new_n860));
  INV_X1    g0660(.A(new_n853), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n792), .B(new_n806), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n862), .A2(new_n857), .B1(new_n836), .B2(new_n840), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n859), .B1(new_n863), .B2(new_n855), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n852), .A2(new_n853), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n497), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n864), .B(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(G330), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n847), .B(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n284), .B2(new_n627), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n222), .B1(new_n260), .B2(KEYINPUT35), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n871), .B(new_n234), .C1(KEYINPUT35), .C2(new_n260), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n872), .B(KEYINPUT36), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n363), .B(new_n748), .C1(G58), .C2(G68), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n203), .A2(G50), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n875), .B(KEYINPUT98), .ZN(new_n876));
  OAI211_X1 g0676(.A(G1), .B(new_n278), .C1(new_n874), .C2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n870), .A2(new_n873), .A3(new_n877), .ZN(G367));
  OR2_X1    g0678(.A1(new_n339), .A2(new_n633), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n327), .A2(new_n329), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n617), .B(new_n633), .C1(new_n880), .C2(new_n288), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n650), .A2(new_n882), .ZN(new_n883));
  XOR2_X1   g0683(.A(new_n883), .B(KEYINPUT104), .Z(new_n884));
  OR2_X1    g0684(.A1(new_n884), .A2(KEYINPUT44), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(KEYINPUT44), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n650), .A2(new_n882), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n887), .B(KEYINPUT45), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n885), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n889), .B(new_n647), .ZN(new_n890));
  INV_X1    g0690(.A(new_n645), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n690), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n646), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n893), .B(new_n648), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n688), .ZN(new_n895));
  OR2_X1    g0695(.A1(new_n890), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n688), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n656), .B(KEYINPUT41), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n691), .ZN(new_n900));
  INV_X1    g0700(.A(new_n882), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n647), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n882), .A2(new_n649), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n903), .B(KEYINPUT42), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n617), .B1(new_n880), .B2(new_n564), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n632), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n529), .A2(new_n633), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n619), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n523), .B2(new_n907), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n904), .A2(new_n906), .B1(KEYINPUT43), .B2(new_n909), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n902), .B(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n909), .A2(KEYINPUT43), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n911), .B(new_n912), .ZN(new_n913));
  OR2_X1    g0713(.A1(new_n909), .A2(new_n760), .ZN(new_n914));
  INV_X1    g0714(.A(new_n746), .ZN(new_n915));
  OAI221_X1 g0715(.A(new_n758), .B1(new_n228), .B2(new_n432), .C1(new_n915), .C2(new_n245), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n694), .ZN(new_n917));
  XOR2_X1   g0717(.A(new_n917), .B(KEYINPUT105), .Z(new_n918));
  INV_X1    g0718(.A(new_n740), .ZN(new_n919));
  AOI22_X1  g0719(.A1(G150), .A2(new_n723), .B1(new_n732), .B2(G50), .ZN(new_n920));
  INV_X1    g0720(.A(G137), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n920), .B1(new_n921), .B2(new_n724), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n769), .A2(new_n466), .B1(new_n730), .B2(new_n768), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n271), .B1(new_n716), .B2(new_n202), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n700), .A2(new_n203), .ZN(new_n925));
  NOR4_X1   g0725(.A1(new_n922), .A2(new_n923), .A3(new_n924), .A4(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n719), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(G77), .ZN(new_n928));
  AOI22_X1  g0728(.A1(G97), .A2(new_n927), .B1(new_n725), .B2(G317), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n568), .B2(new_n722), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n744), .B1(new_n769), .B2(new_n701), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n717), .A2(KEYINPUT46), .A3(G116), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n704), .A2(G311), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n699), .A2(G107), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT46), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n716), .B2(new_n222), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n932), .A2(new_n933), .A3(new_n934), .A4(new_n936), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n930), .A2(new_n931), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n732), .A2(G283), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n926), .A2(new_n928), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT47), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n918), .B1(new_n919), .B2(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT106), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n900), .A2(new_n913), .B1(new_n914), .B2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(G387));
  OR2_X1    g0745(.A1(new_n894), .A2(new_n688), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n946), .A2(new_n656), .A3(new_n895), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n654), .A2(new_n751), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n746), .B1(new_n242), .B2(new_n306), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n341), .A2(G50), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT50), .ZN(new_n951));
  AOI21_X1  g0751(.A(G45), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n951), .B2(new_n950), .ZN(new_n953));
  AOI211_X1 g0753(.A(new_n654), .B(new_n953), .C1(G68), .C2(G77), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n948), .B1(G107), .B2(new_n228), .C1(new_n949), .C2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT107), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n758), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(new_n956), .B2(new_n955), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n725), .A2(G326), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n723), .A2(G317), .B1(G311), .B2(new_n711), .ZN(new_n960));
  XNOR2_X1  g0760(.A(KEYINPUT108), .B(G322), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n704), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n960), .B(new_n962), .C1(new_n568), .C2(new_n709), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT48), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n964), .B1(new_n775), .B2(new_n700), .C1(new_n701), .C2(new_n716), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT49), .ZN(new_n966));
  AOI211_X1 g0766(.A(new_n765), .B(new_n959), .C1(new_n965), .C2(new_n966), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n967), .B1(new_n966), .B2(new_n965), .C1(new_n222), .C2(new_n719), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n716), .A2(new_n363), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n765), .B1(new_n341), .B2(new_n769), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(G159), .B2(new_n704), .ZN(new_n971));
  AOI22_X1  g0771(.A1(G50), .A2(new_n723), .B1(new_n732), .B2(G68), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n343), .B2(new_n724), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(G97), .B2(new_n720), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n971), .B(new_n974), .C1(new_n432), .C2(new_n700), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n968), .B1(new_n969), .B2(new_n975), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT109), .Z(new_n977));
  OAI21_X1  g0777(.A(new_n694), .B1(new_n977), .B2(new_n919), .ZN(new_n978));
  AOI211_X1 g0778(.A(new_n958), .B(new_n978), .C1(new_n891), .C2(new_n757), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(new_n894), .B2(new_n692), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n947), .A2(new_n980), .ZN(G393));
  NAND2_X1  g0781(.A1(new_n890), .A2(new_n895), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n896), .A2(new_n982), .A3(new_n656), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n890), .A2(new_n691), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n271), .B1(new_n725), .B2(new_n961), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n736), .B(new_n985), .C1(new_n775), .C2(new_n716), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT110), .Z(new_n987));
  AOI22_X1  g0787(.A1(new_n723), .A2(G311), .B1(G317), .B2(new_n704), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT52), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(G294), .B2(new_n732), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n699), .A2(G116), .B1(G303), .B2(new_n711), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT111), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n987), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n769), .A2(new_n216), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n994), .B(new_n744), .C1(G77), .C2(new_n699), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n717), .A2(G68), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n730), .A2(new_n343), .B1(new_n722), .B2(new_n466), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT51), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n709), .A2(new_n341), .B1(new_n724), .B2(new_n768), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(new_n720), .B2(G87), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n995), .A2(new_n996), .A3(new_n998), .A4(new_n1000), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n993), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n694), .B1(new_n1002), .B2(new_n919), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n746), .A2(new_n252), .B1(G97), .B2(new_n655), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1003), .B1(new_n758), .B2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT112), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n760), .B2(new_n901), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n983), .A2(new_n984), .A3(new_n1007), .ZN(G390));
  NAND3_X1  g0808(.A1(new_n497), .A2(G330), .A3(new_n865), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n1009), .A2(KEYINPUT113), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1009), .A2(KEYINPUT113), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n846), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT114), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1015));
  AOI21_X1  g0815(.A(KEYINPUT114), .B1(new_n1015), .B2(new_n846), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n844), .B1(new_n801), .B2(new_n807), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n825), .A2(KEYINPUT39), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1018), .B(new_n1019), .C1(KEYINPUT39), .C2(new_n841), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n800), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n665), .B2(new_n791), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(new_n806), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1023), .A2(new_n844), .A3(new_n841), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n792), .A2(new_n687), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1025), .A2(new_n807), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1020), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1027));
  AND2_X1   g0827(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n862), .A2(new_n668), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1025), .A2(new_n807), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1031), .A2(KEYINPUT115), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1032), .A2(new_n801), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1031), .B(KEYINPUT115), .C1(new_n862), .C2(new_n668), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n806), .B1(new_n854), .B2(G330), .ZN(new_n1036));
  OR3_X1    g0836(.A1(new_n1036), .A2(new_n1022), .A3(new_n1026), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1017), .A2(new_n1030), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1029), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n1028), .B2(new_n1026), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1015), .A2(KEYINPUT114), .A3(new_n846), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1042), .A2(new_n1043), .A3(new_n1038), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1041), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1039), .A2(new_n656), .A3(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(KEYINPUT116), .B1(new_n1041), .B2(new_n691), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT116), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1030), .A2(new_n1048), .A3(new_n692), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n843), .A2(new_n755), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n700), .A2(new_n363), .B1(new_n775), .B2(new_n730), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n777), .B1(new_n722), .B2(new_n222), .C1(new_n500), .C2(new_n716), .ZN(new_n1053));
  NOR3_X1   g0853(.A1(new_n764), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n732), .A2(G97), .B1(G107), .B2(new_n711), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT117), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1054), .B(new_n1056), .C1(new_n701), .C2(new_n724), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT118), .Z(new_n1058));
  NOR3_X1   g0858(.A1(new_n716), .A2(KEYINPUT53), .A3(new_n343), .ZN(new_n1059));
  OAI21_X1  g0859(.A(KEYINPUT53), .B1(new_n716), .B2(new_n343), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n769), .B2(new_n921), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n1059), .B(new_n1061), .C1(G128), .C2(new_n704), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n725), .A2(G125), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n722), .A2(new_n773), .B1(new_n719), .B2(new_n216), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n271), .B1(new_n700), .B2(new_n466), .ZN(new_n1065));
  XOR2_X1   g0865(.A(KEYINPUT54), .B(G143), .Z(new_n1066));
  AOI211_X1 g0866(.A(new_n1064), .B(new_n1065), .C1(new_n732), .C2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1062), .A2(new_n1063), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n919), .B1(new_n1058), .B2(new_n1068), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n695), .B(new_n1069), .C1(new_n341), .C2(new_n785), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT119), .Z(new_n1071));
  NAND2_X1  g0871(.A1(new_n1051), .A2(new_n1071), .ZN(new_n1072));
  AND3_X1   g0872(.A1(new_n1046), .A2(new_n1050), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(G378));
  INV_X1    g0874(.A(new_n845), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT122), .ZN(new_n1076));
  AND3_X1   g0876(.A1(new_n864), .A2(new_n1076), .A3(G330), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1076), .B1(new_n864), .B2(G330), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n392), .B1(new_n384), .B2(new_n388), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n358), .A2(new_n631), .ZN(new_n1080));
  AND2_X1   g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1082));
  NOR3_X1   g0882(.A1(new_n1081), .A2(new_n1082), .A3(KEYINPUT55), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(KEYINPUT55), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1085));
  AND3_X1   g0885(.A1(new_n1084), .A2(KEYINPUT56), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(KEYINPUT56), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n1077), .A2(new_n1078), .A3(new_n1088), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1088), .A2(new_n1076), .A3(G330), .A4(new_n864), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1075), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n864), .A2(G330), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(KEYINPUT122), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n864), .A2(new_n1076), .A3(G330), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1088), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1097), .A2(new_n845), .A3(new_n1090), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1092), .A2(KEYINPUT123), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n845), .B1(new_n1097), .B2(new_n1090), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT123), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1038), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1017), .B1(new_n1041), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1099), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT57), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  AND3_X1   g0907(.A1(new_n1097), .A2(new_n845), .A3(new_n1090), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1104), .B(KEYINPUT57), .C1(new_n1108), .C2(new_n1100), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n1109), .A2(new_n656), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1099), .A2(new_n692), .A3(new_n1102), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT124), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n694), .B1(G50), .B2(new_n786), .ZN(new_n1114));
  XOR2_X1   g0914(.A(new_n1114), .B(KEYINPUT121), .Z(new_n1115));
  INV_X1    g0915(.A(new_n371), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n744), .B(new_n1116), .C1(new_n212), .C2(new_n722), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n711), .A2(G97), .B1(new_n704), .B2(G116), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n1118), .B1(new_n363), .B2(new_n716), .C1(new_n432), .C2(new_n709), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n719), .A2(new_n202), .B1(new_n724), .B2(new_n775), .ZN(new_n1120));
  NOR4_X1   g0920(.A1(new_n1117), .A2(new_n1119), .A3(new_n925), .A4(new_n1120), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n1121), .B(KEYINPUT58), .Z(new_n1122));
  AOI22_X1  g0922(.A1(G128), .A2(new_n723), .B1(new_n732), .B2(G137), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n699), .A2(G150), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n717), .A2(new_n1066), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n711), .A2(G132), .B1(new_n704), .B2(G125), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  OR2_X1    g0927(.A1(new_n1127), .A2(KEYINPUT59), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n725), .A2(G124), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1127), .A2(KEYINPUT59), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(G33), .A2(G41), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT120), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(G159), .B2(new_n927), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .A4(new_n1133), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n216), .B(new_n1132), .C1(new_n765), .C2(new_n371), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n1122), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n1115), .B1(new_n919), .B2(new_n1136), .C1(new_n1096), .C2(new_n756), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n1112), .A2(new_n1113), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1113), .B1(new_n1112), .B2(new_n1137), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1111), .B1(new_n1138), .B2(new_n1139), .ZN(G375));
  AOI21_X1  g0940(.A(new_n1038), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1142), .A2(new_n898), .A3(new_n1044), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n222), .A2(new_n769), .B1(new_n730), .B2(new_n701), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n777), .B1(new_n700), .B2(new_n432), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1144), .B(new_n1145), .C1(G283), .C2(new_n723), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n716), .A2(new_n210), .B1(new_n724), .B2(new_n568), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(new_n720), .B2(G77), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1146), .B(new_n1148), .C1(new_n212), .C2(new_n709), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n730), .A2(new_n773), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n744), .B1(G159), .B2(new_n717), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n927), .A2(G58), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(G50), .A2(new_n699), .B1(new_n1066), .B2(new_n711), .ZN(new_n1153));
  INV_X1    g0953(.A(G128), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n709), .A2(new_n343), .B1(new_n724), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(G137), .B2(new_n723), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .A4(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1149), .B1(new_n1150), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n695), .B1(new_n1158), .B2(new_n740), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n806), .B2(new_n756), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n203), .B2(new_n785), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n1038), .B2(new_n692), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1143), .A2(new_n1162), .ZN(G381));
  NAND2_X1  g0963(.A1(new_n1112), .A2(new_n1137), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(KEYINPUT124), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1112), .A2(new_n1113), .A3(new_n1137), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n1165), .A2(new_n1166), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n1073), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n947), .A2(new_n762), .A3(new_n980), .ZN(new_n1169));
  OR3_X1    g0969(.A1(G390), .A2(G384), .A3(new_n1169), .ZN(new_n1170));
  OR4_X1    g0970(.A1(G387), .A2(new_n1168), .A3(G381), .A4(new_n1170), .ZN(G407));
  OAI211_X1 g0971(.A(G407), .B(G213), .C1(G343), .C2(new_n1168), .ZN(G409));
  NAND4_X1  g0972(.A1(new_n1099), .A2(new_n898), .A3(new_n1102), .A4(new_n1104), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n692), .B1(new_n1108), .B2(new_n1100), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1073), .A2(new_n1173), .A3(new_n1137), .A4(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(G343), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(G213), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1141), .A2(KEYINPUT60), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n656), .B(new_n1044), .C1(new_n1141), .C2(KEYINPUT60), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1162), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(G384), .B(KEYINPUT125), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT125), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(G384), .A2(new_n1186), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1162), .B(new_n1187), .C1(new_n1181), .C2(new_n1182), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1185), .A2(new_n1188), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1179), .B(new_n1189), .C1(new_n1167), .C2(new_n1073), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(KEYINPUT62), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1178), .B1(G375), .B2(G378), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT62), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1192), .A2(new_n1193), .A3(new_n1189), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT61), .ZN(new_n1195));
  INV_X1    g0995(.A(G2897), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1177), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT126), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1185), .A2(new_n1200), .A3(new_n1188), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1201), .A2(new_n1203), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1185), .A2(KEYINPUT126), .A3(new_n1197), .A4(new_n1188), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1073), .B1(new_n1208), .B2(new_n1111), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1207), .B1(new_n1209), .B2(new_n1178), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1191), .A2(new_n1194), .A3(new_n1195), .A4(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(G393), .A2(G396), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(G390), .A2(new_n1169), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1169), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1214), .A2(new_n984), .A3(new_n983), .A4(new_n1007), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n944), .A2(new_n1213), .A3(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n944), .B1(new_n1213), .B2(new_n1215), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1211), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(G375), .A2(G378), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1206), .B1(new_n1221), .B2(new_n1179), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT63), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1190), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  NOR3_X1   g1024(.A1(new_n1216), .A2(new_n1217), .A3(KEYINPUT61), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT127), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n1190), .B2(new_n1223), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1192), .A2(KEYINPUT127), .A3(KEYINPUT63), .A4(new_n1189), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1224), .A2(new_n1225), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1220), .A2(new_n1229), .ZN(G405));
  NAND2_X1  g1030(.A1(new_n1168), .A2(new_n1221), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1231), .A2(new_n1185), .A3(new_n1188), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1168), .A2(new_n1221), .A3(new_n1189), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n1219), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1232), .A2(new_n1218), .A3(new_n1233), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(G402));
endmodule


