//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 1 0 0 1 0 0 1 1 0 0 1 1 0 0 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0 1 1 1 1 0 1 1 1 1 1 0 1 1 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n815, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1035, new_n1036;
  XNOR2_X1  g000(.A(KEYINPUT70), .B(G113gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G120gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G127gat), .B(G134gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT71), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OR2_X1    g005(.A1(G113gat), .A2(G120gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT1), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT72), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT72), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT1), .ZN(new_n211));
  AND3_X1   g010(.A1(new_n207), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G127gat), .ZN(new_n213));
  INV_X1    g012(.A(G134gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G127gat), .A2(G134gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n215), .A2(KEYINPUT71), .A3(new_n216), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n203), .A2(new_n206), .A3(new_n212), .A4(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT73), .ZN(new_n219));
  AOI22_X1  g018(.A1(new_n205), .A2(new_n204), .B1(new_n202), .B2(G120gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT73), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n220), .A2(new_n221), .A3(new_n217), .A4(new_n212), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n204), .A2(KEYINPUT69), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT69), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n215), .A2(new_n225), .A3(new_n216), .ZN(new_n226));
  NAND2_X1  g025(.A1(G113gat), .A2(G120gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n207), .A2(new_n208), .A3(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n224), .A2(new_n226), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n223), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT74), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n233), .B1(KEYINPUT23), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT24), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n236), .A2(G183gat), .A3(G190gat), .ZN(new_n237));
  INV_X1    g036(.A(G183gat), .ZN(new_n238));
  INV_X1    g037(.A(G190gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n237), .B1(new_n240), .B2(new_n236), .ZN(new_n241));
  NOR2_X1   g040(.A1(G183gat), .A2(G190gat), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n235), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n233), .A2(KEYINPUT23), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT64), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT25), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  OR2_X1    g049(.A1(new_n242), .A2(KEYINPUT65), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n242), .A2(KEYINPUT65), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n241), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n245), .A2(KEYINPUT25), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n254), .A2(new_n235), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT28), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT27), .B(G183gat), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n238), .A2(KEYINPUT27), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(new_n259), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(new_n239), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n257), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n257), .A2(G190gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n258), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT67), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT67), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n258), .A2(new_n268), .A3(new_n265), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n264), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G169gat), .ZN(new_n271));
  INV_X1    g070(.A(G176gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT68), .B1(new_n273), .B2(KEYINPUT26), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT68), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT26), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n233), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n234), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n279), .B1(KEYINPUT26), .B2(new_n273), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n240), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  AOI22_X1  g080(.A1(new_n250), .A2(new_n256), .B1(new_n270), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n229), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n283), .B1(new_n219), .B2(new_n222), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT74), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n232), .A2(new_n282), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n267), .A2(new_n269), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT27), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(G183gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n261), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT66), .ZN(new_n291));
  AOI21_X1  g090(.A(G190gat), .B1(new_n261), .B2(new_n259), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT28), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n281), .B1(new_n287), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n256), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT25), .B1(new_n244), .B2(new_n247), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n284), .A2(KEYINPUT74), .ZN(new_n298));
  AOI211_X1 g097(.A(new_n231), .B(new_n283), .C1(new_n219), .C2(new_n222), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n286), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(G227gat), .A2(G233gat), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT33), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G15gat), .B(G43gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(G71gat), .B(G99gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n305), .B(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT34), .B1(new_n301), .B2(new_n303), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT34), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n286), .A2(new_n300), .A3(new_n310), .A4(new_n302), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n301), .A2(new_n303), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT32), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n309), .B(new_n311), .C1(new_n304), .C2(new_n307), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n313), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n316), .B1(new_n313), .B2(new_n317), .ZN(new_n320));
  XNOR2_X1  g119(.A(G197gat), .B(G204gat), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT22), .ZN(new_n322));
  INV_X1    g121(.A(G211gat), .ZN(new_n323));
  INV_X1    g122(.A(G218gat), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G211gat), .B(G218gat), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n326), .B(new_n328), .ZN(new_n329));
  XOR2_X1   g128(.A(G141gat), .B(G148gat), .Z(new_n330));
  INV_X1    g129(.A(G155gat), .ZN(new_n331));
  INV_X1    g130(.A(G162gat), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT2), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G155gat), .B(G162gat), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT3), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n330), .A2(new_n335), .A3(new_n333), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT29), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n329), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  AND2_X1   g141(.A1(G228gat), .A2(G233gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n341), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT3), .B1(new_n345), .B2(KEYINPUT77), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n326), .B(new_n327), .ZN(new_n347));
  OR3_X1    g146(.A1(new_n347), .A2(KEYINPUT77), .A3(KEYINPUT29), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n337), .A2(new_n339), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n344), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n351), .B1(new_n345), .B2(new_n338), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n343), .B1(new_n353), .B2(new_n342), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(KEYINPUT31), .B(G50gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n356), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n352), .A2(new_n354), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(G78gat), .B(G106gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(G22gat), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n357), .A2(new_n362), .A3(new_n359), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NOR3_X1   g165(.A1(new_n319), .A2(new_n320), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(G225gat), .A2(G233gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n350), .A2(KEYINPUT3), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(new_n340), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n368), .B1(new_n370), .B2(new_n284), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT4), .B1(new_n284), .B2(new_n351), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n232), .A2(KEYINPUT4), .A3(new_n285), .A4(new_n351), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT5), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n230), .A2(new_n350), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n284), .A2(new_n351), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n368), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n376), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n375), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n284), .A2(KEYINPUT4), .A3(new_n351), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n376), .B(new_n368), .C1(new_n370), .C2(new_n284), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n298), .A2(new_n299), .A3(new_n350), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n383), .B(new_n385), .C1(new_n386), .C2(KEYINPUT4), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n382), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G1gat), .B(G29gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n389), .B(KEYINPUT0), .ZN(new_n390));
  XNOR2_X1  g189(.A(G57gat), .B(G85gat), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n390), .B(new_n391), .Z(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n388), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT6), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n382), .A2(new_n387), .A3(new_n392), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n388), .A2(KEYINPUT6), .A3(new_n393), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  XOR2_X1   g198(.A(G8gat), .B(G36gat), .Z(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(KEYINPUT76), .ZN(new_n401));
  XNOR2_X1  g200(.A(G64gat), .B(G92gat), .ZN(new_n402));
  XOR2_X1   g201(.A(new_n401), .B(new_n402), .Z(new_n403));
  INV_X1    g202(.A(G226gat), .ZN(new_n404));
  INV_X1    g203(.A(G233gat), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n406), .B1(new_n297), .B2(new_n341), .ZN(new_n407));
  INV_X1    g206(.A(new_n406), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n282), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n347), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT75), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n297), .A2(new_n406), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n250), .A2(new_n256), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT29), .B1(new_n413), .B2(new_n294), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n329), .B(new_n412), .C1(new_n414), .C2(new_n406), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n410), .A2(new_n411), .A3(new_n415), .ZN(new_n416));
  OAI211_X1 g215(.A(KEYINPUT75), .B(new_n347), .C1(new_n407), .C2(new_n409), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n403), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n410), .A2(new_n411), .A3(new_n415), .ZN(new_n420));
  INV_X1    g219(.A(new_n403), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n420), .A2(new_n417), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n419), .A2(KEYINPUT30), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT30), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n424), .B(new_n403), .C1(new_n416), .C2(new_n418), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  AND2_X1   g225(.A1(new_n399), .A2(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(KEYINPUT83), .A2(KEYINPUT35), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(KEYINPUT83), .A2(KEYINPUT35), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n367), .A2(new_n427), .A3(new_n429), .A4(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n313), .A2(new_n317), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n315), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n364), .A2(new_n365), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n433), .A2(new_n434), .A3(new_n318), .A4(new_n430), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n399), .A2(new_n426), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n428), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n431), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT38), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n421), .A2(KEYINPUT37), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n422), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n420), .A2(KEYINPUT37), .A3(new_n417), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n439), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT81), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n410), .A2(new_n444), .ZN(new_n445));
  OAI211_X1 g244(.A(KEYINPUT81), .B(new_n347), .C1(new_n407), .C2(new_n409), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n445), .A2(new_n415), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT38), .B1(new_n447), .B2(KEYINPUT37), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n441), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n449), .A2(new_n397), .A3(new_n419), .A4(new_n398), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT82), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n443), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n397), .A2(new_n398), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n453), .A2(KEYINPUT82), .A3(new_n449), .A4(new_n419), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n230), .A2(new_n340), .A3(new_n369), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n456), .B(new_n383), .C1(new_n386), .C2(KEYINPUT4), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n380), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT39), .B1(new_n379), .B2(new_n380), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT39), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n457), .A2(new_n462), .A3(new_n380), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n461), .A2(KEYINPUT40), .A3(new_n392), .A4(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n423), .A2(new_n464), .A3(new_n394), .A4(new_n425), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT80), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT40), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n463), .A2(new_n392), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n459), .B1(new_n457), .B2(new_n380), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT79), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT79), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n473), .B(new_n468), .C1(new_n469), .C2(new_n470), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n466), .A2(new_n467), .A3(new_n472), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n472), .A2(new_n474), .ZN(new_n476));
  OAI21_X1  g275(.A(KEYINPUT80), .B1(new_n476), .B2(new_n465), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n455), .A2(new_n475), .A3(new_n434), .A4(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n433), .A2(KEYINPUT36), .A3(new_n318), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT36), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n480), .B1(new_n319), .B2(new_n320), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n364), .A2(KEYINPUT78), .A3(new_n365), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT78), .B1(new_n364), .B2(new_n365), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n479), .A2(new_n481), .B1(new_n484), .B2(new_n436), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n438), .B1(new_n478), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(G22gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(G15gat), .ZN(new_n488));
  INV_X1    g287(.A(G15gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(G22gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(G1gat), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT87), .B1(new_n492), .B2(KEYINPUT16), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n492), .A2(KEYINPUT87), .A3(KEYINPUT16), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n491), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(G8gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(G15gat), .B(G22gat), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n497), .B1(new_n498), .B2(G1gat), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT88), .B1(new_n498), .B2(G1gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT88), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n492), .A2(KEYINPUT87), .A3(KEYINPUT16), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n498), .B(new_n503), .C1(new_n504), .C2(new_n493), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(G8gat), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT89), .B1(new_n502), .B2(new_n506), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n505), .A2(G8gat), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT89), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n498), .B1(new_n504), .B2(new_n493), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n510), .B(KEYINPUT88), .C1(G1gat), .C2(new_n498), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n508), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n500), .B1(new_n507), .B2(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(G43gat), .B(G50gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT15), .ZN(new_n515));
  INV_X1    g314(.A(G50gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n516), .A2(KEYINPUT86), .A3(G43gat), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT15), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT86), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n519), .B1(new_n520), .B2(new_n514), .ZN(new_n521));
  NAND2_X1  g320(.A1(KEYINPUT85), .A2(G36gat), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(KEYINPUT85), .A2(G36gat), .ZN(new_n524));
  OAI21_X1  g323(.A(G29gat), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT14), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n526), .B1(G29gat), .B2(G36gat), .ZN(new_n527));
  INV_X1    g326(.A(G29gat), .ZN(new_n528));
  INV_X1    g327(.A(G36gat), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(new_n529), .A3(KEYINPUT14), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n525), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n515), .B1(new_n521), .B2(new_n531), .ZN(new_n532));
  OR2_X1    g331(.A1(KEYINPUT85), .A2(G36gat), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n528), .B1(new_n533), .B2(new_n522), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n530), .A2(new_n527), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n515), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n532), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT90), .B1(new_n513), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n500), .ZN(new_n541));
  NOR3_X1   g340(.A1(new_n502), .A2(new_n506), .A3(KEYINPUT89), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n509), .B1(new_n508), .B2(new_n511), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n516), .A2(G43gat), .ZN(new_n545));
  INV_X1    g344(.A(G43gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(G50gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n518), .B(new_n517), .C1(new_n548), .C2(KEYINPUT86), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n537), .B1(new_n536), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n531), .A2(new_n515), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n544), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n540), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G229gat), .A2(G233gat), .ZN(new_n555));
  XOR2_X1   g354(.A(new_n555), .B(KEYINPUT13), .Z(new_n556));
  NAND3_X1  g355(.A1(new_n544), .A2(KEYINPUT90), .A3(new_n552), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n554), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT17), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n559), .B1(new_n550), .B2(new_n551), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n532), .A2(new_n538), .A3(KEYINPUT17), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n513), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n553), .A2(new_n555), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT18), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n553), .A2(KEYINPUT18), .A3(new_n563), .A4(new_n555), .ZN(new_n567));
  XNOR2_X1  g366(.A(G113gat), .B(G141gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G169gat), .B(G197gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT12), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n558), .A2(new_n566), .A3(new_n567), .A4(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT91), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n573), .B1(new_n564), .B2(new_n565), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n578), .A2(KEYINPUT91), .A3(new_n558), .A4(new_n567), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n558), .A2(new_n566), .A3(new_n567), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(new_n573), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G99gat), .A2(G106gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT8), .ZN(new_n586));
  NAND2_X1  g385(.A1(G85gat), .A2(G92gat), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT7), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(G85gat), .ZN(new_n590));
  INV_X1    g389(.A(G92gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n586), .A2(new_n589), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n585), .ZN(new_n595));
  NOR2_X1   g394(.A1(G99gat), .A2(G106gat), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n595), .A2(new_n596), .ZN(new_n599));
  INV_X1    g398(.A(new_n593), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI22_X1  g401(.A1(KEYINPUT8), .A2(new_n585), .B1(new_n590), .B2(new_n591), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n599), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n598), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n562), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(G232gat), .A2(G233gat), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n607), .B(KEYINPUT93), .Z(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT41), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n609), .B1(new_n539), .B2(new_n605), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n239), .B1(new_n606), .B2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n605), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n613), .B1(new_n560), .B2(new_n561), .ZN(new_n614));
  NOR3_X1   g413(.A1(new_n614), .A2(new_n610), .A3(G190gat), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n324), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT95), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n606), .A2(new_n611), .A3(new_n239), .ZN(new_n618));
  OAI21_X1  g417(.A(G190gat), .B1(new_n614), .B2(new_n610), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n618), .A2(G218gat), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n616), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  OR2_X1    g420(.A1(new_n608), .A2(KEYINPUT41), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n622), .B(KEYINPUT94), .Z(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G134gat), .B(G162gat), .ZN(new_n625));
  INV_X1    g424(.A(new_n623), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n616), .A2(new_n617), .A3(new_n626), .A4(new_n620), .ZN(new_n627));
  AND3_X1   g426(.A1(new_n624), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n625), .B1(new_n624), .B2(new_n627), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT92), .ZN(new_n631));
  AND2_X1   g430(.A1(G71gat), .A2(G78gat), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n631), .B1(new_n632), .B2(KEYINPUT9), .ZN(new_n633));
  INV_X1    g432(.A(G57gat), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(G64gat), .ZN(new_n635));
  INV_X1    g434(.A(G64gat), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(G57gat), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(KEYINPUT92), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n633), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G71gat), .B(G78gat), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  AOI22_X1  g443(.A1(new_n635), .A2(new_n637), .B1(new_n639), .B2(KEYINPUT92), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n645), .A2(new_n642), .A3(new_n633), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT21), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(G231gat), .A2(G233gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(G127gat), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n513), .B1(new_n648), .B2(new_n647), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(G155gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(G183gat), .B(G211gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n654), .B(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT96), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n594), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n599), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n594), .A2(new_n597), .A3(new_n661), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n663), .A2(new_n644), .A3(new_n646), .A4(new_n664), .ZN(new_n665));
  AND4_X1   g464(.A1(new_n642), .A2(new_n633), .A3(new_n638), .A4(new_n640), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n642), .B1(new_n645), .B2(new_n633), .ZN(new_n667));
  OAI22_X1  g466(.A1(new_n666), .A2(new_n667), .B1(new_n598), .B2(new_n604), .ZN(new_n668));
  INV_X1    g467(.A(G230gat), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n669), .A2(new_n405), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n665), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n671), .A2(KEYINPUT97), .ZN(new_n672));
  INV_X1    g471(.A(new_n670), .ZN(new_n673));
  AOI21_X1  g472(.A(KEYINPUT10), .B1(new_n665), .B2(new_n668), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT10), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n647), .A2(new_n605), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n673), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n671), .A2(KEYINPUT97), .ZN(new_n678));
  XNOR2_X1  g477(.A(G120gat), .B(G148gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(G176gat), .B(G204gat), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n679), .B(new_n680), .Z(new_n681));
  NAND4_X1  g480(.A1(new_n672), .A2(new_n677), .A3(new_n678), .A4(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n677), .A2(new_n671), .ZN(new_n683));
  INV_X1    g482(.A(new_n681), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT98), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT98), .ZN(new_n686));
  AOI211_X1 g485(.A(new_n686), .B(new_n681), .C1(new_n677), .C2(new_n671), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n682), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT99), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI211_X1 g489(.A(KEYINPUT99), .B(new_n682), .C1(new_n685), .C2(new_n687), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n630), .A2(new_n660), .A3(new_n693), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n486), .A2(new_n584), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n453), .A2(KEYINPUT100), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT100), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n399), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(G1gat), .ZN(G1324gat));
  INV_X1    g500(.A(new_n426), .ZN(new_n702));
  XOR2_X1   g501(.A(KEYINPUT16), .B(G8gat), .Z(new_n703));
  NAND3_X1  g502(.A1(new_n695), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT42), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n486), .A2(new_n584), .ZN(new_n707));
  INV_X1    g506(.A(new_n694), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(G8gat), .B1(new_n709), .B2(new_n426), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n710), .A2(new_n704), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n706), .B1(new_n711), .B2(new_n705), .ZN(G1325gat));
  NAND2_X1  g511(.A1(new_n481), .A2(new_n479), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT101), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(G15gat), .B1(new_n709), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n319), .A2(new_n320), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n695), .A2(new_n489), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(G1326gat));
  INV_X1    g519(.A(new_n484), .ZN(new_n721));
  OAI21_X1  g520(.A(KEYINPUT102), .B1(new_n709), .B2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT102), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n695), .A2(new_n723), .A3(new_n484), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g524(.A(KEYINPUT43), .B(G22gat), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n722), .A2(new_n724), .A3(new_n726), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(G1327gat));
  NOR3_X1   g529(.A1(new_n630), .A2(new_n660), .A3(new_n692), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n486), .A2(new_n584), .A3(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n733), .A2(new_n528), .A3(new_n699), .ZN(new_n734));
  XNOR2_X1  g533(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n734), .B(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n475), .A2(new_n477), .A3(new_n434), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n452), .A2(new_n454), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n485), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n438), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n630), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(KEYINPUT44), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(new_n486), .B2(new_n630), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n692), .B(KEYINPUT104), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n747), .A2(new_n584), .A3(new_n660), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n743), .A2(new_n745), .A3(new_n699), .A4(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT105), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G29gat), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n749), .A2(new_n750), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n737), .B1(new_n752), .B2(new_n753), .ZN(G1328gat));
  INV_X1    g553(.A(KEYINPUT46), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n523), .A2(new_n524), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n426), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n733), .A2(new_n755), .A3(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT106), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n743), .A2(new_n745), .A3(new_n748), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n757), .B1(new_n762), .B2(new_n426), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n733), .A2(new_n758), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(KEYINPUT46), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n761), .A2(new_n763), .A3(new_n765), .ZN(G1329gat));
  INV_X1    g565(.A(new_n713), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n743), .A2(new_n745), .A3(new_n767), .A4(new_n748), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(G43gat), .ZN(new_n769));
  INV_X1    g568(.A(new_n718), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n770), .A2(G43gat), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n733), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n769), .A2(KEYINPUT47), .A3(new_n772), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n743), .A2(new_n745), .A3(new_n715), .A4(new_n748), .ZN(new_n774));
  AOI22_X1  g573(.A1(new_n774), .A2(G43gat), .B1(new_n733), .B2(new_n771), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(KEYINPUT47), .B2(new_n775), .ZN(G1330gat));
  NAND4_X1  g575(.A1(new_n743), .A2(new_n745), .A3(new_n366), .A4(new_n748), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(G50gat), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n740), .A2(new_n741), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n779), .A2(new_n583), .A3(new_n731), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT107), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT107), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n707), .A2(new_n782), .A3(new_n731), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n721), .A2(G50gat), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n781), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n778), .A2(KEYINPUT48), .A3(new_n785), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n743), .A2(new_n745), .A3(new_n484), .A4(new_n748), .ZN(new_n787));
  INV_X1    g586(.A(new_n784), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n788), .B1(new_n733), .B2(new_n782), .ZN(new_n789));
  AOI22_X1  g588(.A1(G50gat), .A2(new_n787), .B1(new_n789), .B2(new_n781), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n786), .B1(new_n790), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g590(.A(new_n629), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n624), .A2(new_n625), .A3(new_n627), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n654), .B(new_n658), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n779), .A2(new_n584), .A3(new_n796), .A4(new_n747), .ZN(new_n797));
  INV_X1    g596(.A(new_n699), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(new_n634), .ZN(G1332gat));
  NOR2_X1   g599(.A1(new_n797), .A2(new_n426), .ZN(new_n801));
  NOR2_X1   g600(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n802));
  AND2_X1   g601(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n804), .B1(new_n801), .B2(new_n802), .ZN(G1333gat));
  INV_X1    g604(.A(KEYINPUT50), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n797), .A2(new_n716), .ZN(new_n807));
  INV_X1    g606(.A(G71gat), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n718), .A2(new_n808), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n797), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n806), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  OAI221_X1 g611(.A(KEYINPUT50), .B1(new_n797), .B2(new_n810), .C1(new_n807), .C2(new_n808), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(G1334gat));
  NOR2_X1   g613(.A1(new_n797), .A2(new_n721), .ZN(new_n815));
  XOR2_X1   g614(.A(new_n815), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g615(.A1(new_n660), .A2(new_n583), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n779), .A2(new_n794), .A3(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT51), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n742), .A2(KEYINPUT51), .A3(new_n817), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n822), .A2(new_n590), .A3(new_n692), .A4(new_n699), .ZN(new_n823));
  INV_X1    g622(.A(new_n817), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n824), .A2(new_n693), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n743), .A2(new_n745), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(G85gat), .B1(new_n826), .B2(new_n798), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n823), .A2(new_n827), .ZN(G1336gat));
  NAND4_X1  g627(.A1(new_n743), .A2(new_n745), .A3(new_n702), .A4(new_n825), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(G92gat), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT52), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n746), .A2(G92gat), .A3(new_n426), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(KEYINPUT108), .ZN(new_n833));
  AOI21_X1  g632(.A(KEYINPUT51), .B1(new_n742), .B2(new_n817), .ZN(new_n834));
  NOR4_X1   g633(.A1(new_n486), .A2(new_n819), .A3(new_n630), .A4(new_n824), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n830), .A2(new_n831), .A3(new_n836), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n833), .B(KEYINPUT109), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n822), .A2(new_n838), .B1(new_n829), .B2(G92gat), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n837), .B1(new_n839), .B2(new_n831), .ZN(G1337gat));
  NOR2_X1   g639(.A1(new_n770), .A2(G99gat), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n822), .A2(new_n692), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(G99gat), .B1(new_n826), .B2(new_n716), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(G1338gat));
  NAND4_X1  g643(.A1(new_n743), .A2(new_n745), .A3(new_n366), .A4(new_n825), .ZN(new_n845));
  XNOR2_X1  g644(.A(KEYINPUT110), .B(G106gat), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n746), .A2(G106gat), .A3(new_n434), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n848), .B1(new_n834), .B2(new_n835), .ZN(new_n849));
  XNOR2_X1  g648(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n847), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n743), .A2(new_n745), .A3(new_n484), .A4(new_n825), .ZN(new_n852));
  AOI22_X1  g651(.A1(new_n822), .A2(new_n848), .B1(new_n852), .B2(new_n846), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n851), .B1(new_n853), .B2(new_n854), .ZN(G1339gat));
  NAND2_X1  g654(.A1(new_n708), .A2(new_n584), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n556), .B1(new_n554), .B2(new_n557), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n555), .B1(new_n553), .B2(new_n563), .ZN(new_n858));
  OR2_X1    g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n572), .ZN(new_n860));
  AOI22_X1  g659(.A1(new_n577), .A2(new_n579), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n861), .B1(new_n628), .B2(new_n629), .ZN(new_n862));
  OR3_X1    g661(.A1(new_n674), .A2(new_n676), .A3(new_n673), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n863), .A2(KEYINPUT54), .A3(new_n677), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n865), .B(new_n673), .C1(new_n674), .C2(new_n676), .ZN(new_n866));
  AND3_X1   g665(.A1(new_n866), .A2(KEYINPUT112), .A3(new_n684), .ZN(new_n867));
  AOI21_X1  g666(.A(KEYINPUT112), .B1(new_n866), .B2(new_n684), .ZN(new_n868));
  OAI211_X1 g667(.A(KEYINPUT55), .B(new_n864), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT113), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n869), .A2(new_n870), .A3(new_n682), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n864), .B1(new_n867), .B2(new_n868), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT55), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n869), .A2(new_n682), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(KEYINPUT113), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n862), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n859), .A2(new_n860), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n692), .A2(new_n580), .A3(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT114), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n583), .A2(new_n877), .A3(new_n875), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n861), .A2(KEYINPUT114), .A3(new_n692), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n879), .B1(new_n886), .B2(new_n630), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n856), .B1(new_n887), .B2(new_n660), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n888), .A2(new_n699), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n367), .A2(new_n426), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OR3_X1    g690(.A1(new_n891), .A2(new_n584), .A3(new_n202), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n798), .A2(new_n702), .A3(new_n770), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n888), .A2(KEYINPUT115), .A3(new_n721), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(KEYINPUT115), .B1(new_n888), .B2(new_n721), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n583), .B(new_n893), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT116), .ZN(new_n898));
  AND3_X1   g697(.A1(new_n897), .A2(new_n898), .A3(G113gat), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(new_n897), .B2(G113gat), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n892), .B1(new_n899), .B2(new_n900), .ZN(G1340gat));
  NOR2_X1   g700(.A1(new_n891), .A2(new_n693), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n902), .A2(G120gat), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n721), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT115), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n894), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n893), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n747), .A2(G120gat), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n903), .B1(new_n909), .B2(new_n910), .ZN(G1341gat));
  NOR2_X1   g710(.A1(new_n795), .A2(new_n213), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n907), .A2(new_n893), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT117), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n213), .B1(new_n891), .B2(new_n795), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n913), .A2(KEYINPUT117), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n916), .A2(new_n917), .ZN(G1342gat));
  NAND4_X1  g717(.A1(new_n889), .A2(new_n214), .A3(new_n794), .A4(new_n890), .ZN(new_n919));
  XOR2_X1   g718(.A(new_n919), .B(KEYINPUT56), .Z(new_n920));
  OAI21_X1  g719(.A(G134gat), .B1(new_n908), .B2(new_n630), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1343gat));
  NOR3_X1   g721(.A1(new_n767), .A2(new_n798), .A3(new_n702), .ZN(new_n923));
  AOI21_X1  g722(.A(KEYINPUT57), .B1(new_n888), .B2(new_n366), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n484), .A2(KEYINPUT57), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT118), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n876), .B1(new_n873), .B2(new_n872), .ZN(new_n927));
  AOI22_X1  g726(.A1(new_n881), .A2(new_n926), .B1(new_n583), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n861), .A2(KEYINPUT118), .A3(new_n692), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n794), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n795), .B1(new_n930), .B2(new_n879), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n925), .B1(new_n931), .B2(new_n856), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n923), .B1(new_n924), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(G141gat), .B1(new_n933), .B2(new_n584), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n715), .A2(new_n702), .A3(new_n434), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n889), .A2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(G141gat), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n936), .A2(new_n937), .A3(new_n583), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n934), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(KEYINPUT58), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT58), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n934), .A2(new_n938), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n940), .A2(new_n942), .ZN(G1344gat));
  XOR2_X1   g742(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n944));
  INV_X1    g743(.A(KEYINPUT57), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n945), .B1(new_n888), .B2(new_n366), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n484), .A2(new_n945), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n796), .A2(KEYINPUT121), .A3(new_n584), .A4(new_n693), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT121), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n949), .B1(new_n694), .B2(new_n583), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n947), .B1(new_n951), .B2(new_n931), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n923), .A2(new_n692), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n946), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(G148gat), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n944), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI211_X1 g755(.A(new_n692), .B(new_n923), .C1(new_n924), .C2(new_n932), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT119), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n955), .A2(KEYINPUT59), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n958), .B1(new_n957), .B2(new_n959), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n956), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n936), .A2(new_n955), .A3(new_n692), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(G1345gat));
  NAND3_X1  g763(.A1(new_n889), .A2(new_n935), .A3(new_n660), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT122), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n331), .B1(new_n965), .B2(new_n966), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n660), .A2(G155gat), .ZN(new_n969));
  OAI22_X1  g768(.A1(new_n967), .A2(new_n968), .B1(new_n933), .B2(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(G1346gat));
  AND4_X1   g770(.A1(new_n332), .A2(new_n889), .A3(new_n935), .A4(new_n794), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT123), .ZN(new_n973));
  OAI21_X1  g772(.A(G162gat), .B1(new_n933), .B2(new_n630), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(G1347gat));
  AND2_X1   g774(.A1(new_n888), .A2(new_n798), .ZN(new_n976));
  AND2_X1   g775(.A1(new_n367), .A2(new_n702), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g777(.A(new_n978), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n979), .A2(new_n271), .A3(new_n583), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n699), .A2(new_n426), .ZN(new_n981));
  OR2_X1    g780(.A1(new_n981), .A2(KEYINPUT124), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(KEYINPUT124), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n982), .A2(new_n718), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n984), .B1(new_n906), .B2(new_n894), .ZN(new_n985));
  AOI211_X1 g784(.A(KEYINPUT125), .B(new_n271), .C1(new_n985), .C2(new_n583), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT125), .ZN(new_n987));
  INV_X1    g786(.A(new_n984), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n907), .A2(new_n583), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n987), .B1(new_n989), .B2(G169gat), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n980), .B1(new_n986), .B2(new_n990), .ZN(G1348gat));
  AOI21_X1  g790(.A(new_n272), .B1(new_n985), .B2(new_n747), .ZN(new_n992));
  NOR3_X1   g791(.A1(new_n978), .A2(G176gat), .A3(new_n693), .ZN(new_n993));
  OR2_X1    g792(.A1(new_n992), .A2(new_n993), .ZN(G1349gat));
  AOI21_X1  g793(.A(new_n238), .B1(new_n985), .B2(new_n660), .ZN(new_n995));
  NOR3_X1   g794(.A1(new_n978), .A2(new_n290), .A3(new_n795), .ZN(new_n996));
  OAI21_X1  g795(.A(KEYINPUT60), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g796(.A(new_n996), .ZN(new_n998));
  INV_X1    g797(.A(KEYINPUT60), .ZN(new_n999));
  OAI211_X1 g798(.A(new_n660), .B(new_n988), .C1(new_n895), .C2(new_n896), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n1000), .A2(G183gat), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n997), .A2(new_n1002), .ZN(G1350gat));
  NAND3_X1  g802(.A1(new_n907), .A2(new_n794), .A3(new_n988), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1004), .A2(G190gat), .ZN(new_n1005));
  INV_X1    g804(.A(KEYINPUT61), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n1004), .A2(KEYINPUT61), .A3(G190gat), .ZN(new_n1008));
  NAND4_X1  g807(.A1(new_n976), .A2(new_n239), .A3(new_n794), .A4(new_n977), .ZN(new_n1009));
  INV_X1    g808(.A(KEYINPUT126), .ZN(new_n1010));
  XNOR2_X1  g809(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  NAND3_X1  g810(.A1(new_n1007), .A2(new_n1008), .A3(new_n1011), .ZN(G1351gat));
  NOR3_X1   g811(.A1(new_n715), .A2(new_n426), .A3(new_n434), .ZN(new_n1013));
  AND2_X1   g812(.A1(new_n976), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g813(.A(G197gat), .B1(new_n1014), .B2(new_n583), .ZN(new_n1015));
  NOR2_X1   g814(.A1(new_n946), .A2(new_n952), .ZN(new_n1016));
  INV_X1    g815(.A(new_n1016), .ZN(new_n1017));
  AND2_X1   g816(.A1(new_n982), .A2(new_n983), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n1018), .A2(new_n716), .ZN(new_n1019));
  NOR2_X1   g818(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  AND2_X1   g819(.A1(new_n583), .A2(G197gat), .ZN(new_n1021));
  AOI21_X1  g820(.A(new_n1015), .B1(new_n1020), .B2(new_n1021), .ZN(G1352gat));
  XNOR2_X1  g821(.A(KEYINPUT127), .B(G204gat), .ZN(new_n1023));
  NAND3_X1  g822(.A1(new_n1014), .A2(new_n692), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g823(.A1(new_n1024), .A2(KEYINPUT62), .ZN(new_n1025));
  INV_X1    g824(.A(KEYINPUT62), .ZN(new_n1026));
  NAND4_X1  g825(.A1(new_n1014), .A2(new_n1026), .A3(new_n692), .A4(new_n1023), .ZN(new_n1027));
  NOR3_X1   g826(.A1(new_n1017), .A2(new_n746), .A3(new_n1019), .ZN(new_n1028));
  OAI211_X1 g827(.A(new_n1025), .B(new_n1027), .C1(new_n1028), .C2(new_n1023), .ZN(G1353gat));
  NAND3_X1  g828(.A1(new_n1014), .A2(new_n323), .A3(new_n660), .ZN(new_n1030));
  NAND4_X1  g829(.A1(new_n1016), .A2(new_n660), .A3(new_n716), .A4(new_n1018), .ZN(new_n1031));
  AND3_X1   g830(.A1(new_n1031), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1032));
  AOI21_X1  g831(.A(KEYINPUT63), .B1(new_n1031), .B2(G211gat), .ZN(new_n1033));
  OAI21_X1  g832(.A(new_n1030), .B1(new_n1032), .B2(new_n1033), .ZN(G1354gat));
  NAND3_X1  g833(.A1(new_n1014), .A2(new_n324), .A3(new_n794), .ZN(new_n1035));
  NOR3_X1   g834(.A1(new_n1017), .A2(new_n630), .A3(new_n1019), .ZN(new_n1036));
  OAI21_X1  g835(.A(new_n1035), .B1(new_n1036), .B2(new_n324), .ZN(G1355gat));
endmodule


