//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0 0 1 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 0 1 1 1 0 1 0 0 0 0 0 1 1 1 0 1 0 0 0 0 1 0 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n625, new_n626, new_n627, new_n630, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1187, new_n1188, new_n1189;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT66), .Z(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(new_n455), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(KEYINPUT69), .B1(new_n463), .B2(G2105), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT69), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(new_n466), .A3(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g043(.A(KEYINPUT70), .B1(new_n468), .B2(G101), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT70), .ZN(new_n470));
  INV_X1    g045(.A(G101), .ZN(new_n471));
  AOI211_X1 g046(.A(new_n470), .B(new_n471), .C1(new_n464), .C2(new_n467), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n473), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n474));
  OAI22_X1  g049(.A1(new_n469), .A2(new_n472), .B1(new_n466), .B2(new_n474), .ZN(new_n475));
  AND2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  OAI211_X1 g052(.A(G137), .B(new_n466), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n478), .B(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n475), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT71), .ZN(G160));
  OR2_X1    g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NAND2_X1  g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  AOI21_X1  g059(.A(G2105), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n466), .B1(new_n483), .B2(new_n484), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  OR2_X1    g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n486), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  OAI211_X1 g067(.A(G126), .B(G2105), .C1(new_n476), .C2(new_n477), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n495), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g072(.A(G138), .B(new_n466), .C1(new_n476), .C2(new_n477), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n473), .A2(new_n500), .A3(G138), .A4(new_n466), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n497), .B1(new_n499), .B2(new_n501), .ZN(G164));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT72), .A2(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT72), .A2(G651), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT6), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n503), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G50), .ZN(new_n510));
  XNOR2_X1  g085(.A(new_n510), .B(KEYINPUT73), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n514), .B1(new_n506), .B2(new_n508), .ZN(new_n515));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G62), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n504), .A2(new_n505), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n515), .A2(G88), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n511), .A2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  INV_X1    g098(.A(G63), .ZN(new_n524));
  INV_X1    g099(.A(G651), .ZN(new_n525));
  NOR3_X1   g100(.A1(new_n514), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n526), .B1(new_n509), .B2(G51), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(KEYINPUT74), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XOR2_X1   g104(.A(new_n529), .B(KEYINPUT7), .Z(new_n530));
  AOI21_X1  g105(.A(new_n530), .B1(new_n515), .B2(G89), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n527), .A2(KEYINPUT74), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(G168));
  INV_X1    g111(.A(new_n514), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n537), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n538), .A2(new_n519), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n515), .A2(G90), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n509), .A2(G52), .ZN(new_n541));
  AND3_X1   g116(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(G171));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n514), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(new_n520), .ZN(new_n546));
  XOR2_X1   g121(.A(new_n546), .B(KEYINPUT75), .Z(new_n547));
  AOI22_X1  g122(.A1(G43), .A2(new_n509), .B1(new_n515), .B2(G81), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT76), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  INV_X1    g131(.A(KEYINPUT6), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT72), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(new_n525), .ZN(new_n559));
  NAND2_X1  g134(.A1(KEYINPUT72), .A2(G651), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n557), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI211_X1 g136(.A(G53), .B(G543), .C1(new_n561), .C2(new_n507), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n562), .A2(KEYINPUT9), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n564), .B1(new_n509), .B2(G53), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g141(.A(KEYINPUT78), .B(G65), .ZN(new_n567));
  OR2_X1    g142(.A1(KEYINPUT5), .A2(G543), .ZN(new_n568));
  NAND2_X1  g143(.A1(KEYINPUT5), .A2(G543), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n568), .A2(KEYINPUT77), .A3(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT77), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n571), .B1(new_n512), .B2(new_n513), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n567), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  AND2_X1   g148(.A1(G78), .A2(G543), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n515), .A2(G91), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OR3_X1    g152(.A1(new_n566), .A2(new_n577), .A3(KEYINPUT79), .ZN(new_n578));
  OAI21_X1  g153(.A(KEYINPUT79), .B1(new_n566), .B2(new_n577), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G299));
  INV_X1    g156(.A(G171), .ZN(G301));
  INV_X1    g157(.A(KEYINPUT80), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n532), .A2(new_n583), .A3(new_n534), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n528), .A2(new_n531), .ZN(new_n585));
  OAI21_X1  g160(.A(KEYINPUT80), .B1(new_n585), .B2(new_n533), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G286));
  NAND2_X1  g163(.A1(new_n515), .A2(G87), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n509), .A2(G49), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n537), .B2(G74), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(G288));
  NAND2_X1  g167(.A1(new_n515), .A2(G86), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT82), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n515), .A2(KEYINPUT82), .A3(G86), .ZN(new_n596));
  AND2_X1   g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(G73), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G61), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n514), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(new_n520), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(KEYINPUT81), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT81), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n600), .A2(new_n603), .A3(new_n520), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n602), .A2(new_n604), .B1(G48), .B2(new_n509), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n597), .A2(new_n605), .ZN(G305));
  NAND2_X1  g181(.A1(new_n515), .A2(G85), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n509), .A2(G47), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n537), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n609));
  OAI211_X1 g184(.A(new_n607), .B(new_n608), .C1(new_n519), .C2(new_n609), .ZN(G290));
  NAND2_X1  g185(.A1(G301), .A2(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  AND2_X1   g187(.A1(new_n570), .A2(new_n572), .ZN(new_n613));
  INV_X1    g188(.A(G66), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G651), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n509), .A2(G54), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n515), .A2(G92), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT10), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n611), .B1(new_n621), .B2(G868), .ZN(G284));
  OAI21_X1  g197(.A(new_n611), .B1(new_n621), .B2(G868), .ZN(G321));
  AND3_X1   g198(.A1(G286), .A2(KEYINPUT83), .A3(G868), .ZN(new_n624));
  AOI21_X1  g199(.A(G868), .B1(new_n580), .B2(KEYINPUT84), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(KEYINPUT84), .B2(new_n580), .ZN(new_n626));
  AOI21_X1  g201(.A(KEYINPUT83), .B1(G286), .B2(G868), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n624), .B1(new_n626), .B2(new_n627), .ZN(G297));
  AOI21_X1  g203(.A(new_n624), .B1(new_n626), .B2(new_n627), .ZN(G280));
  INV_X1    g204(.A(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n621), .B1(new_n630), .B2(G860), .ZN(G148));
  NAND2_X1  g206(.A1(new_n621), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G868), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g210(.A1(new_n468), .A2(new_n473), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  INV_X1    g213(.A(G2100), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n485), .A2(G135), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n487), .A2(G123), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n466), .A2(G111), .ZN(new_n644));
  OAI21_X1  g219(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n642), .B(new_n643), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(G2096), .Z(new_n647));
  NAND3_X1  g222(.A1(new_n640), .A2(new_n641), .A3(new_n647), .ZN(G156));
  XOR2_X1   g223(.A(G2451), .B(G2454), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(KEYINPUT14), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2427), .B(G2438), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2430), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT15), .B(G2435), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n657), .B1(new_n656), .B2(new_n655), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n652), .B(new_n658), .Z(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2443), .B(G2446), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(G14), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n662), .B2(new_n660), .ZN(G401));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT85), .B(KEYINPUT18), .Z(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n665), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT86), .Z(new_n672));
  NAND2_X1  g247(.A1(new_n668), .A2(KEYINPUT17), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n666), .A2(new_n667), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n669), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n672), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2096), .B(G2100), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G227));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n681), .A2(KEYINPUT87), .ZN(new_n682));
  XOR2_X1   g257(.A(G1971), .B(G1976), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(KEYINPUT87), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n682), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT20), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n679), .A2(new_n680), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(new_n681), .ZN(new_n689));
  MUX2_X1   g264(.A(new_n689), .B(new_n688), .S(new_n684), .Z(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT88), .ZN(new_n692));
  XOR2_X1   g267(.A(G1991), .B(G1996), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(G1981), .B(G1986), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT89), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n694), .B(new_n698), .ZN(G229));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NOR2_X1   g275(.A1(G171), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(G5), .B2(new_n700), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G35), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G162), .B2(new_n704), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT29), .Z(new_n707));
  INV_X1    g282(.A(G2090), .ZN(new_n708));
  AOI22_X1  g283(.A1(G1961), .A2(new_n703), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT25), .Z(new_n711));
  INV_X1    g286(.A(G139), .ZN(new_n712));
  INV_X1    g287(.A(new_n485), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT94), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n473), .A2(G127), .ZN(new_n716));
  AND2_X1   g291(.A1(G115), .A2(G2104), .ZN(new_n717));
  OAI21_X1  g292(.A(G2105), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  MUX2_X1   g294(.A(G33), .B(new_n719), .S(G29), .Z(new_n720));
  OAI221_X1 g295(.A(new_n709), .B1(G1961), .B2(new_n703), .C1(G2072), .C2(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n550), .A2(new_n700), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n700), .B2(G19), .ZN(new_n723));
  INV_X1    g298(.A(G1341), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n723), .A2(new_n724), .ZN(new_n726));
  NOR2_X1   g301(.A1(G27), .A2(G29), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G164), .B2(G29), .ZN(new_n728));
  INV_X1    g303(.A(G2078), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n720), .A2(G2072), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n725), .A2(new_n726), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n621), .A2(G16), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G4), .B2(G16), .ZN(new_n734));
  INV_X1    g309(.A(G1348), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n734), .A2(new_n735), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n485), .A2(G140), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n487), .A2(G128), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n466), .A2(G116), .ZN(new_n740));
  OAI21_X1  g315(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n738), .B(new_n739), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(G29), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n704), .A2(G26), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT28), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G2067), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  XOR2_X1   g323(.A(KEYINPUT31), .B(G11), .Z(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT30), .B(G28), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n749), .B1(new_n704), .B2(new_n750), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n704), .A2(G32), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT96), .B(KEYINPUT26), .Z(new_n753));
  NAND3_X1  g328(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  AOI22_X1  g330(.A1(G129), .A2(new_n487), .B1(new_n485), .B2(G141), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n468), .A2(G105), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n755), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n752), .B1(new_n758), .B2(G29), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT27), .B(G1996), .Z(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT97), .ZN(new_n761));
  OAI221_X1 g336(.A(new_n751), .B1(new_n704), .B2(new_n646), .C1(new_n759), .C2(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n761), .B2(new_n759), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n737), .A2(new_n748), .A3(new_n763), .ZN(new_n764));
  NOR4_X1   g339(.A1(new_n721), .A2(new_n732), .A3(new_n736), .A4(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G34), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n766), .A2(KEYINPUT24), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n766), .A2(KEYINPUT24), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n704), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G160), .B2(new_n704), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT95), .B(G2084), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n700), .A2(G20), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT23), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n580), .B2(new_n700), .ZN(new_n775));
  INV_X1    g350(.A(G1956), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n707), .A2(new_n708), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT98), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n700), .A2(G21), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G168), .B2(new_n700), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n781), .A2(G1966), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n781), .A2(G1966), .ZN(new_n783));
  NOR3_X1   g358(.A1(new_n779), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n765), .A2(new_n772), .A3(new_n777), .A4(new_n784), .ZN(new_n785));
  MUX2_X1   g360(.A(G6), .B(G305), .S(G16), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT93), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT32), .B(G1981), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  MUX2_X1   g364(.A(G23), .B(G288), .S(G16), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT33), .ZN(new_n791));
  INV_X1    g366(.A(G1976), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(G16), .A2(G22), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G166), .B2(G16), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G1971), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n789), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(KEYINPUT34), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT34), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n789), .A2(new_n800), .A3(new_n797), .ZN(new_n801));
  MUX2_X1   g376(.A(G24), .B(G290), .S(G16), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1986), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n704), .A2(G25), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT90), .Z(new_n805));
  OAI21_X1  g380(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n806));
  INV_X1    g381(.A(G107), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(G2105), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT91), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n487), .A2(G119), .ZN(new_n810));
  INV_X1    g385(.A(G131), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(new_n713), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n805), .B1(new_n814), .B2(G29), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT35), .B(G1991), .Z(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT92), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n815), .B(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n803), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n799), .A2(new_n801), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(KEYINPUT36), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT36), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n799), .A2(new_n822), .A3(new_n801), .A4(new_n819), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n785), .B1(new_n821), .B2(new_n823), .ZN(G311));
  INV_X1    g399(.A(G311), .ZN(G150));
  NAND2_X1  g400(.A1(new_n621), .A2(G559), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT38), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n509), .A2(G55), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n537), .B1(new_n561), .B2(new_n507), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT99), .B(G93), .Z(new_n830));
  AOI22_X1  g405(.A1(new_n537), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n831));
  OAI221_X1 g406(.A(new_n828), .B1(new_n829), .B2(new_n830), .C1(new_n519), .C2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n549), .B(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n827), .B(new_n834), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n835), .A2(KEYINPUT39), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(KEYINPUT39), .ZN(new_n837));
  NOR3_X1   g412(.A1(new_n836), .A2(new_n837), .A3(G860), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n832), .A2(G860), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT37), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n838), .A2(new_n840), .ZN(G145));
  INV_X1    g416(.A(G37), .ZN(new_n842));
  AOI22_X1  g417(.A1(G130), .A2(new_n487), .B1(new_n485), .B2(G142), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT100), .ZN(new_n844));
  NOR3_X1   g419(.A1(new_n844), .A2(new_n466), .A3(G118), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n844), .B1(new_n466), .B2(G118), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n846), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n843), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT101), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n637), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n814), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n851), .A2(KEYINPUT102), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(KEYINPUT102), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n719), .B(new_n758), .ZN(new_n854));
  XNOR2_X1  g429(.A(G164), .B(new_n742), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n852), .A2(new_n853), .A3(new_n856), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n853), .A2(new_n856), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(G160), .B(new_n646), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n491), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n842), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n859), .A2(new_n861), .ZN(new_n864));
  AOI21_X1  g439(.A(KEYINPUT40), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n864), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT40), .ZN(new_n867));
  NOR3_X1   g442(.A1(new_n866), .A2(new_n862), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n865), .A2(new_n868), .ZN(G395));
  XNOR2_X1  g444(.A(new_n833), .B(new_n632), .ZN(new_n870));
  NAND2_X1  g445(.A1(G299), .A2(new_n621), .ZN(new_n871));
  INV_X1    g446(.A(new_n621), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n580), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n875), .A2(KEYINPUT103), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(KEYINPUT103), .ZN(new_n877));
  AND3_X1   g452(.A1(new_n871), .A2(KEYINPUT41), .A3(new_n873), .ZN(new_n878));
  AOI21_X1  g453(.A(KEYINPUT41), .B1(new_n871), .B2(new_n873), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n876), .B(new_n877), .C1(new_n870), .C2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(G166), .A2(G305), .ZN(new_n882));
  NAND3_X1  g457(.A1(G303), .A2(new_n605), .A3(new_n597), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(G290), .B(G288), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n884), .A2(new_n886), .ZN(new_n889));
  NOR3_X1   g464(.A1(new_n888), .A2(KEYINPUT42), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT104), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n891), .B1(new_n888), .B2(new_n889), .ZN(new_n892));
  INV_X1    g467(.A(new_n889), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n893), .A2(KEYINPUT104), .A3(new_n887), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n890), .B1(new_n895), .B2(KEYINPUT42), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n881), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n881), .A2(new_n896), .ZN(new_n898));
  OAI21_X1  g473(.A(G868), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(G868), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n832), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(G295));
  NAND2_X1  g477(.A1(new_n899), .A2(new_n901), .ZN(G331));
  NAND3_X1  g478(.A1(new_n584), .A2(G171), .A3(new_n586), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT105), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n905), .B1(new_n535), .B2(G171), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n584), .A2(new_n586), .A3(new_n905), .A4(G171), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(new_n833), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n833), .B1(new_n907), .B2(new_n908), .ZN(new_n911));
  OAI22_X1  g486(.A1(new_n910), .A2(new_n911), .B1(new_n878), .B2(new_n879), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n907), .A2(new_n908), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(new_n834), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n914), .A2(new_n874), .A3(new_n909), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n895), .A2(new_n912), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(new_n842), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n895), .B1(new_n912), .B2(new_n915), .ZN(new_n918));
  OAI21_X1  g493(.A(KEYINPUT43), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT107), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n871), .A2(new_n873), .A3(KEYINPUT41), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT41), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n874), .A2(new_n922), .ZN(new_n923));
  AOI22_X1  g498(.A1(new_n921), .A2(new_n923), .B1(new_n914), .B2(new_n909), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n914), .A2(new_n874), .A3(new_n909), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT106), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n912), .A2(new_n927), .A3(new_n915), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n926), .A2(new_n894), .A3(new_n892), .A4(new_n928), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n916), .A2(new_n842), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n933), .B(KEYINPUT43), .C1(new_n917), .C2(new_n918), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n920), .A2(KEYINPUT44), .A3(new_n932), .A4(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n931), .B1(new_n929), .B2(new_n930), .ZN(new_n937));
  NOR3_X1   g512(.A1(new_n917), .A2(KEYINPUT43), .A3(new_n918), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n935), .A2(new_n939), .ZN(G397));
  INV_X1    g515(.A(KEYINPUT110), .ZN(new_n941));
  OR2_X1    g516(.A1(G288), .A2(G1976), .ZN(new_n942));
  INV_X1    g517(.A(G1981), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n597), .A2(new_n943), .A3(new_n605), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n509), .A2(G48), .ZN(new_n945));
  INV_X1    g520(.A(new_n604), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n603), .B1(new_n600), .B2(new_n520), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n945), .B(new_n593), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(G1981), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n944), .A2(new_n949), .A3(KEYINPUT49), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT109), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT109), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n944), .A2(new_n949), .A3(new_n952), .A4(KEYINPUT49), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT49), .B1(new_n944), .B2(new_n949), .ZN(new_n955));
  INV_X1    g530(.A(G8), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n471), .B1(new_n464), .B2(new_n467), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n957), .B(KEYINPUT70), .ZN(new_n958));
  OR2_X1    g533(.A1(new_n474), .A2(new_n466), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n478), .B(KEYINPUT68), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n958), .A2(new_n959), .A3(G40), .A4(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n499), .A2(new_n501), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n493), .A2(new_n496), .ZN(new_n963));
  AOI21_X1  g538(.A(G1384), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n961), .A2(new_n965), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n955), .A2(new_n956), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n942), .B1(new_n954), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n944), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n941), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n966), .A2(new_n956), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NOR3_X1   g547(.A1(new_n968), .A2(new_n941), .A3(new_n969), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT55), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n974), .B1(G166), .B2(new_n956), .ZN(new_n975));
  NAND3_X1  g550(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G40), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n475), .A2(new_n978), .A3(new_n480), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n980), .B1(G164), .B2(G1384), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n500), .B1(new_n485), .B2(G138), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n963), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G1384), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n984), .A2(KEYINPUT45), .A3(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n979), .A2(new_n981), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G1971), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT108), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT50), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n990), .B1(new_n964), .B2(new_n991), .ZN(new_n992));
  OAI211_X1 g567(.A(KEYINPUT108), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n964), .A2(new_n991), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n992), .A2(new_n979), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n989), .B1(G2090), .B2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n977), .A2(G8), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n954), .A2(new_n967), .ZN(new_n998));
  OAI221_X1 g573(.A(G8), .B1(new_n792), .B2(G288), .C1(new_n961), .C2(new_n965), .ZN(new_n999));
  AND2_X1   g574(.A1(new_n999), .A2(KEYINPUT52), .ZN(new_n1000));
  INV_X1    g575(.A(new_n999), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT52), .B1(G288), .B2(new_n792), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1000), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n998), .A2(new_n1003), .ZN(new_n1004));
  OAI22_X1  g579(.A1(new_n972), .A2(new_n973), .B1(new_n997), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT57), .B1(new_n566), .B2(new_n577), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT116), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n575), .A2(new_n1008), .A3(new_n576), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1008), .B1(new_n575), .B2(new_n576), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT115), .B1(new_n563), .B2(new_n565), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT57), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n562), .A2(KEYINPUT9), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n509), .A2(new_n564), .A3(G53), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT115), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1012), .A2(new_n1013), .A3(new_n1017), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1006), .B(new_n1007), .C1(new_n1011), .C2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT57), .B1(new_n1021), .B2(KEYINPUT115), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n1022), .B(new_n1017), .C1(new_n1010), .C2(new_n1009), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1006), .B1(new_n1023), .B2(new_n1007), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT111), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1025), .B1(new_n964), .B2(new_n991), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n961), .B1(new_n1026), .B2(new_n994), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n964), .A2(new_n1025), .A3(new_n991), .ZN(new_n1028));
  AOI21_X1  g603(.A(G1956), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n964), .A2(KEYINPUT45), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1030), .A2(new_n961), .ZN(new_n1031));
  XNOR2_X1  g606(.A(KEYINPUT56), .B(G2072), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1031), .A2(new_n986), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  OAI22_X1  g609(.A1(new_n1020), .A2(new_n1024), .B1(new_n1029), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(KEYINPUT119), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT119), .ZN(new_n1037));
  OAI221_X1 g612(.A(new_n1037), .B1(new_n1029), .B2(new_n1034), .C1(new_n1020), .C2(new_n1024), .ZN(new_n1038));
  AOI22_X1  g613(.A1(new_n995), .A2(new_n735), .B1(new_n747), .B2(new_n966), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1036), .B(new_n1038), .C1(new_n872), .C2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1007), .B1(new_n1011), .B2(new_n1018), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT117), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n991), .B1(new_n984), .B2(new_n985), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n994), .B1(new_n1043), .B2(KEYINPUT111), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1044), .A2(new_n979), .A3(new_n1028), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n776), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1042), .A2(new_n1046), .A3(new_n1019), .A4(new_n1033), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT118), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1029), .A2(new_n1034), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1050), .A2(KEYINPUT118), .A3(new_n1042), .A4(new_n1019), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1040), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT61), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1054), .B1(new_n1055), .B2(new_n1050), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1056), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n995), .A2(new_n735), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n966), .A2(new_n747), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT60), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n872), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT122), .ZN(new_n1063));
  AND4_X1   g638(.A1(new_n1063), .A2(new_n1058), .A3(KEYINPUT60), .A4(new_n1059), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1063), .B1(new_n1039), .B2(KEYINPUT60), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1062), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT122), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n621), .B1(new_n1039), .B2(KEYINPUT60), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1039), .A2(new_n1063), .A3(KEYINPUT60), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1066), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n549), .B1(KEYINPUT121), .B2(KEYINPUT59), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n1073), .B(new_n724), .ZN(new_n1074));
  OAI22_X1  g649(.A1(new_n987), .A2(G1996), .B1(new_n966), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1072), .A2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1077));
  XOR2_X1   g652(.A(new_n1076), .B(new_n1077), .Z(new_n1078));
  NAND3_X1  g653(.A1(new_n1057), .A2(new_n1071), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT61), .B1(new_n1052), .B2(new_n1035), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1053), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT124), .ZN(new_n1082));
  INV_X1    g657(.A(G1961), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n995), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT114), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n964), .A2(new_n1085), .A3(KEYINPUT45), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n986), .A2(KEYINPUT114), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1088), .A2(G2078), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1031), .A2(new_n1086), .A3(new_n1087), .A4(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n979), .A2(new_n729), .A3(new_n981), .A4(new_n986), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n1088), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1084), .A2(new_n1090), .A3(new_n1092), .A4(G301), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT54), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1083), .A2(new_n995), .B1(new_n1091), .B2(new_n1088), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT123), .B1(new_n1030), .B2(new_n961), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT123), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n979), .A2(new_n1097), .A3(new_n981), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1096), .A2(new_n1098), .A3(new_n986), .A4(new_n1089), .ZN(new_n1099));
  AOI21_X1  g674(.A(G301), .B1(new_n1095), .B2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1082), .B1(new_n1094), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1099), .A2(new_n1084), .A3(new_n1092), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(G171), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1103), .A2(KEYINPUT124), .A3(KEYINPUT54), .A4(new_n1093), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1087), .A2(new_n981), .A3(new_n979), .A4(new_n1086), .ZN(new_n1106));
  INV_X1    g681(.A(G1966), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NOR3_X1   g683(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1109), .A2(new_n961), .ZN(new_n1110));
  INV_X1    g685(.A(G2084), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1110), .A2(new_n1111), .A3(new_n993), .A4(new_n992), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1108), .A2(new_n1112), .A3(G168), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(G8), .ZN(new_n1114));
  AOI21_X1  g689(.A(G168), .B1(new_n1108), .B2(new_n1112), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT51), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT51), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1113), .A2(new_n1117), .A3(G8), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT54), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1102), .A2(G171), .ZN(new_n1121));
  AOI21_X1  g696(.A(G301), .B1(new_n1095), .B2(new_n1090), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1120), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1105), .A2(new_n1119), .A3(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1044), .A2(new_n708), .A3(new_n979), .A4(new_n1028), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n1125), .A2(KEYINPUT112), .A3(new_n989), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT112), .B1(new_n1125), .B2(new_n989), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1126), .A2(new_n1127), .A3(new_n956), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT113), .B1(new_n1128), .B2(new_n977), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n998), .A2(new_n997), .A3(new_n1003), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1127), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1125), .A2(KEYINPUT112), .A3(new_n989), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1131), .A2(G8), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT113), .ZN(new_n1134));
  INV_X1    g709(.A(new_n977), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1129), .A2(new_n1130), .A3(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1124), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1005), .B1(new_n1081), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n995), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1140), .A2(new_n1111), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1141));
  NOR3_X1   g716(.A1(new_n1141), .A2(G286), .A3(new_n956), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n996), .A2(G8), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1135), .A2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1130), .A2(KEYINPUT63), .A3(new_n1142), .A4(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1142), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1137), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1145), .B1(new_n1147), .B2(KEYINPUT63), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1119), .A2(KEYINPUT62), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT62), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1116), .A2(new_n1118), .A3(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1150), .A2(new_n1122), .A3(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1149), .B1(new_n1153), .B2(new_n1137), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1137), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n1152), .A2(new_n1122), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1155), .A2(new_n1156), .A3(KEYINPUT125), .A4(new_n1150), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1139), .A2(new_n1148), .A3(new_n1154), .A4(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n961), .A2(new_n981), .ZN(new_n1159));
  INV_X1    g734(.A(G1996), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n758), .B(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n742), .B(new_n747), .ZN(new_n1162));
  OR2_X1    g737(.A1(new_n813), .A2(new_n817), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n813), .A2(new_n817), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(G290), .B(G1986), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1159), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1158), .A2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(G290), .A2(G1986), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1159), .A2(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g745(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  AND2_X1   g747(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1173));
  AOI211_X1 g748(.A(new_n1172), .B(new_n1173), .C1(new_n1159), .C2(new_n1165), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1162), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1159), .B1(new_n1175), .B2(new_n758), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT46), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1177), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1178));
  NOR4_X1   g753(.A1(new_n961), .A2(new_n981), .A3(KEYINPUT46), .A4(G1996), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1176), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  XOR2_X1   g755(.A(new_n1180), .B(KEYINPUT47), .Z(new_n1181));
  NAND2_X1  g756(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1182));
  OAI22_X1  g757(.A1(new_n1182), .A2(new_n1164), .B1(G2067), .B2(new_n742), .ZN(new_n1183));
  AOI211_X1 g758(.A(new_n1174), .B(new_n1181), .C1(new_n1159), .C2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1168), .A2(new_n1184), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g760(.A1(new_n937), .A2(new_n938), .ZN(new_n1187));
  NOR4_X1   g761(.A1(G229), .A2(new_n461), .A3(G401), .A4(G227), .ZN(new_n1188));
  OAI21_X1  g762(.A(new_n1188), .B1(new_n866), .B2(new_n862), .ZN(new_n1189));
  NOR2_X1   g763(.A1(new_n1187), .A2(new_n1189), .ZN(G308));
  OAI221_X1 g764(.A(new_n1188), .B1(new_n866), .B2(new_n862), .C1(new_n937), .C2(new_n938), .ZN(G225));
endmodule


