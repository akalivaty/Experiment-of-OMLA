

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U550 ( .A1(G2104), .A2(n525), .ZN(n885) );
  NOR2_X1 U551 ( .A1(n725), .A2(n946), .ZN(n682) );
  AND2_X1 U552 ( .A1(n685), .A2(n517), .ZN(n691) );
  XNOR2_X1 U553 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X1 U554 ( .A1(G164), .A2(G1384), .ZN(n759) );
  AND2_X1 U555 ( .A1(n787), .A2(n973), .ZN(n515) );
  XOR2_X1 U556 ( .A(n724), .B(KEYINPUT92), .Z(n516) );
  AND2_X1 U557 ( .A1(n684), .A2(n683), .ZN(n517) );
  INV_X1 U558 ( .A(KEYINPUT26), .ZN(n681) );
  INV_X1 U559 ( .A(n709), .ZN(n710) );
  NAND2_X1 U560 ( .A1(n710), .A2(G8), .ZN(n711) );
  OR2_X1 U561 ( .A1(n720), .A2(n711), .ZN(n712) );
  INV_X1 U562 ( .A(KEYINPUT29), .ZN(n704) );
  XNOR2_X1 U563 ( .A(KEYINPUT91), .B(KEYINPUT31), .ZN(n716) );
  XNOR2_X1 U564 ( .A(n717), .B(n716), .ZN(n718) );
  AND2_X1 U565 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U566 ( .A1(n759), .A2(n677), .ZN(n725) );
  NAND2_X1 U567 ( .A1(G8), .A2(n725), .ZN(n789) );
  INV_X1 U568 ( .A(KEYINPUT64), .ZN(n518) );
  NAND2_X1 U569 ( .A1(G160), .A2(G40), .ZN(n758) );
  XNOR2_X1 U570 ( .A(n518), .B(KEYINPUT17), .ZN(n519) );
  INV_X1 U571 ( .A(G2104), .ZN(n524) );
  NOR2_X1 U572 ( .A1(G651), .A2(n614), .ZN(n641) );
  NOR2_X1 U573 ( .A1(G2105), .A2(G2104), .ZN(n520) );
  XNOR2_X2 U574 ( .A(n520), .B(n519), .ZN(n881) );
  NAND2_X1 U575 ( .A1(G138), .A2(n881), .ZN(n522) );
  INV_X1 U576 ( .A(G2105), .ZN(n525) );
  NAND2_X1 U577 ( .A1(n885), .A2(G126), .ZN(n521) );
  AND2_X1 U578 ( .A1(n522), .A2(n521), .ZN(n529) );
  NOR2_X4 U579 ( .A1(G2105), .A2(n524), .ZN(n880) );
  NAND2_X1 U580 ( .A1(G102), .A2(n880), .ZN(n523) );
  XOR2_X1 U581 ( .A(KEYINPUT78), .B(n523), .Z(n527) );
  NOR2_X1 U582 ( .A1(n525), .A2(n524), .ZN(n884) );
  AND2_X1 U583 ( .A1(n884), .A2(G114), .ZN(n526) );
  NOR2_X1 U584 ( .A1(n527), .A2(n526), .ZN(n528) );
  NAND2_X1 U585 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U586 ( .A(n530), .B(KEYINPUT79), .ZN(G164) );
  INV_X1 U587 ( .A(G651), .ZN(n535) );
  NOR2_X1 U588 ( .A1(G543), .A2(n535), .ZN(n531) );
  XOR2_X1 U589 ( .A(KEYINPUT1), .B(n531), .Z(n634) );
  NAND2_X1 U590 ( .A1(G64), .A2(n634), .ZN(n534) );
  XNOR2_X1 U591 ( .A(G543), .B(KEYINPUT0), .ZN(n532) );
  XNOR2_X1 U592 ( .A(n532), .B(KEYINPUT65), .ZN(n614) );
  NAND2_X1 U593 ( .A1(G52), .A2(n641), .ZN(n533) );
  NAND2_X1 U594 ( .A1(n534), .A2(n533), .ZN(n540) );
  NOR2_X1 U595 ( .A1(G651), .A2(G543), .ZN(n635) );
  NAND2_X1 U596 ( .A1(G90), .A2(n635), .ZN(n537) );
  NOR2_X1 U597 ( .A1(n614), .A2(n535), .ZN(n636) );
  NAND2_X1 U598 ( .A1(G77), .A2(n636), .ZN(n536) );
  NAND2_X1 U599 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U600 ( .A(KEYINPUT9), .B(n538), .Z(n539) );
  NOR2_X1 U601 ( .A1(n540), .A2(n539), .ZN(G171) );
  INV_X1 U602 ( .A(G171), .ZN(G301) );
  AND2_X1 U603 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U604 ( .A1(G111), .A2(n884), .ZN(n542) );
  NAND2_X1 U605 ( .A1(G135), .A2(n881), .ZN(n541) );
  NAND2_X1 U606 ( .A1(n542), .A2(n541), .ZN(n545) );
  NAND2_X1 U607 ( .A1(n885), .A2(G123), .ZN(n543) );
  XOR2_X1 U608 ( .A(KEYINPUT18), .B(n543), .Z(n544) );
  NOR2_X1 U609 ( .A1(n545), .A2(n544), .ZN(n547) );
  NAND2_X1 U610 ( .A1(n880), .A2(G99), .ZN(n546) );
  NAND2_X1 U611 ( .A1(n547), .A2(n546), .ZN(n914) );
  XNOR2_X1 U612 ( .A(G2096), .B(n914), .ZN(n548) );
  OR2_X1 U613 ( .A1(G2100), .A2(n548), .ZN(G156) );
  NAND2_X1 U614 ( .A1(n885), .A2(G125), .ZN(n550) );
  NAND2_X1 U615 ( .A1(G137), .A2(n881), .ZN(n549) );
  NAND2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n555) );
  NAND2_X1 U617 ( .A1(n884), .A2(G113), .ZN(n553) );
  NAND2_X1 U618 ( .A1(G101), .A2(n880), .ZN(n551) );
  XOR2_X1 U619 ( .A(KEYINPUT23), .B(n551), .Z(n552) );
  NAND2_X1 U620 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U621 ( .A1(n555), .A2(n554), .ZN(G160) );
  INV_X1 U622 ( .A(G57), .ZN(G237) );
  INV_X1 U623 ( .A(G132), .ZN(G219) );
  INV_X1 U624 ( .A(G82), .ZN(G220) );
  NAND2_X1 U625 ( .A1(G63), .A2(n634), .ZN(n557) );
  NAND2_X1 U626 ( .A1(G51), .A2(n641), .ZN(n556) );
  NAND2_X1 U627 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U628 ( .A(KEYINPUT6), .B(n558), .ZN(n565) );
  NAND2_X1 U629 ( .A1(n635), .A2(G89), .ZN(n559) );
  XNOR2_X1 U630 ( .A(n559), .B(KEYINPUT4), .ZN(n561) );
  NAND2_X1 U631 ( .A1(G76), .A2(n636), .ZN(n560) );
  NAND2_X1 U632 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U633 ( .A(KEYINPUT5), .B(n562), .ZN(n563) );
  XNOR2_X1 U634 ( .A(KEYINPUT69), .B(n563), .ZN(n564) );
  NOR2_X1 U635 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U636 ( .A(KEYINPUT7), .B(n566), .Z(G168) );
  XOR2_X1 U637 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U638 ( .A1(G7), .A2(G661), .ZN(n567) );
  XNOR2_X1 U639 ( .A(n567), .B(KEYINPUT68), .ZN(n568) );
  XOR2_X1 U640 ( .A(KEYINPUT10), .B(n568), .Z(n911) );
  NAND2_X1 U641 ( .A1(n911), .A2(G567), .ZN(n569) );
  XOR2_X1 U642 ( .A(KEYINPUT11), .B(n569), .Z(G234) );
  NAND2_X1 U643 ( .A1(G56), .A2(n634), .ZN(n570) );
  XOR2_X1 U644 ( .A(KEYINPUT14), .B(n570), .Z(n576) );
  NAND2_X1 U645 ( .A1(n635), .A2(G81), .ZN(n571) );
  XNOR2_X1 U646 ( .A(n571), .B(KEYINPUT12), .ZN(n573) );
  NAND2_X1 U647 ( .A1(G68), .A2(n636), .ZN(n572) );
  NAND2_X1 U648 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U649 ( .A(KEYINPUT13), .B(n574), .Z(n575) );
  NOR2_X1 U650 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U651 ( .A1(n641), .A2(G43), .ZN(n577) );
  NAND2_X1 U652 ( .A1(n578), .A2(n577), .ZN(n983) );
  INV_X1 U653 ( .A(G860), .ZN(n611) );
  OR2_X1 U654 ( .A1(n983), .A2(n611), .ZN(G153) );
  NAND2_X1 U655 ( .A1(G868), .A2(G301), .ZN(n587) );
  NAND2_X1 U656 ( .A1(G66), .A2(n634), .ZN(n580) );
  NAND2_X1 U657 ( .A1(G92), .A2(n635), .ZN(n579) );
  NAND2_X1 U658 ( .A1(n580), .A2(n579), .ZN(n584) );
  NAND2_X1 U659 ( .A1(G79), .A2(n636), .ZN(n582) );
  NAND2_X1 U660 ( .A1(G54), .A2(n641), .ZN(n581) );
  NAND2_X1 U661 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U662 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U663 ( .A(KEYINPUT15), .B(n585), .ZN(n898) );
  INV_X1 U664 ( .A(G868), .ZN(n644) );
  NAND2_X1 U665 ( .A1(n898), .A2(n644), .ZN(n586) );
  NAND2_X1 U666 ( .A1(n587), .A2(n586), .ZN(G284) );
  NAND2_X1 U667 ( .A1(G91), .A2(n635), .ZN(n589) );
  NAND2_X1 U668 ( .A1(G78), .A2(n636), .ZN(n588) );
  NAND2_X1 U669 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U670 ( .A(KEYINPUT66), .B(n590), .ZN(n594) );
  NAND2_X1 U671 ( .A1(G65), .A2(n634), .ZN(n592) );
  NAND2_X1 U672 ( .A1(G53), .A2(n641), .ZN(n591) );
  NAND2_X1 U673 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U674 ( .A1(n594), .A2(n593), .ZN(n970) );
  XNOR2_X1 U675 ( .A(n970), .B(KEYINPUT67), .ZN(G299) );
  NOR2_X1 U676 ( .A1(G868), .A2(G299), .ZN(n596) );
  NOR2_X1 U677 ( .A1(G286), .A2(n644), .ZN(n595) );
  NOR2_X1 U678 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U679 ( .A(KEYINPUT70), .B(n597), .ZN(G297) );
  NAND2_X1 U680 ( .A1(n611), .A2(G559), .ZN(n598) );
  INV_X1 U681 ( .A(n898), .ZN(n966) );
  NAND2_X1 U682 ( .A1(n598), .A2(n966), .ZN(n599) );
  XNOR2_X1 U683 ( .A(n599), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U684 ( .A1(G868), .A2(n983), .ZN(n602) );
  NAND2_X1 U685 ( .A1(n966), .A2(G868), .ZN(n600) );
  NOR2_X1 U686 ( .A1(G559), .A2(n600), .ZN(n601) );
  NOR2_X1 U687 ( .A1(n602), .A2(n601), .ZN(G282) );
  NAND2_X1 U688 ( .A1(G67), .A2(n634), .ZN(n604) );
  NAND2_X1 U689 ( .A1(G93), .A2(n635), .ZN(n603) );
  NAND2_X1 U690 ( .A1(n604), .A2(n603), .ZN(n607) );
  NAND2_X1 U691 ( .A1(n636), .A2(G80), .ZN(n605) );
  XOR2_X1 U692 ( .A(KEYINPUT72), .B(n605), .Z(n606) );
  NOR2_X1 U693 ( .A1(n607), .A2(n606), .ZN(n609) );
  NAND2_X1 U694 ( .A1(n641), .A2(G55), .ZN(n608) );
  NAND2_X1 U695 ( .A1(n609), .A2(n608), .ZN(n646) );
  NAND2_X1 U696 ( .A1(G559), .A2(n966), .ZN(n610) );
  XOR2_X1 U697 ( .A(n983), .B(n610), .Z(n652) );
  NAND2_X1 U698 ( .A1(n611), .A2(n652), .ZN(n612) );
  XNOR2_X1 U699 ( .A(n612), .B(KEYINPUT71), .ZN(n613) );
  XOR2_X1 U700 ( .A(n646), .B(n613), .Z(G145) );
  NAND2_X1 U701 ( .A1(G49), .A2(n641), .ZN(n616) );
  NAND2_X1 U702 ( .A1(G87), .A2(n614), .ZN(n615) );
  NAND2_X1 U703 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U704 ( .A1(n634), .A2(n617), .ZN(n619) );
  NAND2_X1 U705 ( .A1(G651), .A2(G74), .ZN(n618) );
  NAND2_X1 U706 ( .A1(n619), .A2(n618), .ZN(G288) );
  NAND2_X1 U707 ( .A1(G62), .A2(n634), .ZN(n621) );
  NAND2_X1 U708 ( .A1(G88), .A2(n635), .ZN(n620) );
  NAND2_X1 U709 ( .A1(n621), .A2(n620), .ZN(n624) );
  NAND2_X1 U710 ( .A1(G75), .A2(n636), .ZN(n622) );
  XNOR2_X1 U711 ( .A(KEYINPUT73), .B(n622), .ZN(n623) );
  NOR2_X1 U712 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U713 ( .A1(n641), .A2(G50), .ZN(n625) );
  NAND2_X1 U714 ( .A1(n626), .A2(n625), .ZN(G303) );
  NAND2_X1 U715 ( .A1(G61), .A2(n634), .ZN(n628) );
  NAND2_X1 U716 ( .A1(G86), .A2(n635), .ZN(n627) );
  NAND2_X1 U717 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U718 ( .A1(n636), .A2(G73), .ZN(n629) );
  XOR2_X1 U719 ( .A(KEYINPUT2), .B(n629), .Z(n630) );
  NOR2_X1 U720 ( .A1(n631), .A2(n630), .ZN(n633) );
  NAND2_X1 U721 ( .A1(n641), .A2(G48), .ZN(n632) );
  NAND2_X1 U722 ( .A1(n633), .A2(n632), .ZN(G305) );
  AND2_X1 U723 ( .A1(n634), .A2(G60), .ZN(n640) );
  NAND2_X1 U724 ( .A1(G85), .A2(n635), .ZN(n638) );
  NAND2_X1 U725 ( .A1(G72), .A2(n636), .ZN(n637) );
  NAND2_X1 U726 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U727 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U728 ( .A1(n641), .A2(G47), .ZN(n642) );
  NAND2_X1 U729 ( .A1(n643), .A2(n642), .ZN(G290) );
  NAND2_X1 U730 ( .A1(n644), .A2(n646), .ZN(n645) );
  XNOR2_X1 U731 ( .A(n645), .B(KEYINPUT74), .ZN(n655) );
  XNOR2_X1 U732 ( .A(KEYINPUT19), .B(G288), .ZN(n651) );
  XOR2_X1 U733 ( .A(n646), .B(G305), .Z(n647) );
  XNOR2_X1 U734 ( .A(n647), .B(G299), .ZN(n648) );
  XOR2_X1 U735 ( .A(G303), .B(n648), .Z(n649) );
  XNOR2_X1 U736 ( .A(n649), .B(G290), .ZN(n650) );
  XNOR2_X1 U737 ( .A(n651), .B(n650), .ZN(n897) );
  XNOR2_X1 U738 ( .A(n897), .B(n652), .ZN(n653) );
  NAND2_X1 U739 ( .A1(G868), .A2(n653), .ZN(n654) );
  NAND2_X1 U740 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U741 ( .A(KEYINPUT75), .B(n656), .Z(G295) );
  NAND2_X1 U742 ( .A1(G2084), .A2(G2078), .ZN(n658) );
  XOR2_X1 U743 ( .A(KEYINPUT76), .B(KEYINPUT20), .Z(n657) );
  XNOR2_X1 U744 ( .A(n658), .B(n657), .ZN(n659) );
  NAND2_X1 U745 ( .A1(G2090), .A2(n659), .ZN(n660) );
  XNOR2_X1 U746 ( .A(KEYINPUT21), .B(n660), .ZN(n661) );
  NAND2_X1 U747 ( .A1(n661), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U748 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U749 ( .A1(G220), .A2(G219), .ZN(n662) );
  XOR2_X1 U750 ( .A(KEYINPUT22), .B(n662), .Z(n663) );
  NOR2_X1 U751 ( .A1(G218), .A2(n663), .ZN(n664) );
  NAND2_X1 U752 ( .A1(G96), .A2(n664), .ZN(n831) );
  NAND2_X1 U753 ( .A1(G2106), .A2(n831), .ZN(n668) );
  NAND2_X1 U754 ( .A1(G69), .A2(G120), .ZN(n665) );
  NOR2_X1 U755 ( .A1(G237), .A2(n665), .ZN(n666) );
  NAND2_X1 U756 ( .A1(G108), .A2(n666), .ZN(n832) );
  NAND2_X1 U757 ( .A1(G567), .A2(n832), .ZN(n667) );
  NAND2_X1 U758 ( .A1(n668), .A2(n667), .ZN(n833) );
  NAND2_X1 U759 ( .A1(G661), .A2(G483), .ZN(n669) );
  XOR2_X1 U760 ( .A(KEYINPUT77), .B(n669), .Z(n670) );
  NOR2_X1 U761 ( .A1(n833), .A2(n670), .ZN(n830) );
  NAND2_X1 U762 ( .A1(n830), .A2(G36), .ZN(G176) );
  INV_X1 U763 ( .A(KEYINPUT86), .ZN(n673) );
  NAND2_X1 U764 ( .A1(n758), .A2(n673), .ZN(n676) );
  INV_X1 U765 ( .A(n758), .ZN(n674) );
  NAND2_X1 U766 ( .A1(KEYINPUT86), .A2(n674), .ZN(n675) );
  NAND2_X1 U767 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U768 ( .A1(G2084), .A2(n725), .ZN(n709) );
  NAND2_X1 U769 ( .A1(G8), .A2(n709), .ZN(n722) );
  NOR2_X1 U770 ( .A1(G1966), .A2(n789), .ZN(n720) );
  XOR2_X1 U771 ( .A(KEYINPUT25), .B(G2078), .Z(n945) );
  NOR2_X1 U772 ( .A1(n945), .A2(n725), .ZN(n678) );
  XOR2_X1 U773 ( .A(KEYINPUT88), .B(n678), .Z(n680) );
  XNOR2_X1 U774 ( .A(G1961), .B(KEYINPUT87), .ZN(n994) );
  NAND2_X1 U775 ( .A1(n725), .A2(n994), .ZN(n679) );
  NAND2_X1 U776 ( .A1(n680), .A2(n679), .ZN(n708) );
  NAND2_X1 U777 ( .A1(n708), .A2(G171), .ZN(n707) );
  XNOR2_X1 U778 ( .A(G1996), .B(KEYINPUT89), .ZN(n946) );
  XNOR2_X1 U779 ( .A(n682), .B(n681), .ZN(n685) );
  NAND2_X1 U780 ( .A1(n725), .A2(G1341), .ZN(n684) );
  INV_X1 U781 ( .A(n983), .ZN(n683) );
  NAND2_X1 U782 ( .A1(n691), .A2(n966), .ZN(n689) );
  INV_X1 U783 ( .A(n725), .ZN(n695) );
  NOR2_X1 U784 ( .A1(n695), .A2(G1348), .ZN(n687) );
  NOR2_X1 U785 ( .A1(G2067), .A2(n725), .ZN(n686) );
  NOR2_X1 U786 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U787 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U788 ( .A(n690), .B(KEYINPUT90), .ZN(n693) );
  OR2_X1 U789 ( .A1(n966), .A2(n691), .ZN(n692) );
  NAND2_X1 U790 ( .A1(n693), .A2(n692), .ZN(n699) );
  NAND2_X1 U791 ( .A1(n695), .A2(G2072), .ZN(n694) );
  XNOR2_X1 U792 ( .A(n694), .B(KEYINPUT27), .ZN(n697) );
  INV_X1 U793 ( .A(G1956), .ZN(n969) );
  NOR2_X1 U794 ( .A1(n969), .A2(n695), .ZN(n696) );
  NOR2_X1 U795 ( .A1(n697), .A2(n696), .ZN(n700) );
  NAND2_X1 U796 ( .A1(n970), .A2(n700), .ZN(n698) );
  NAND2_X1 U797 ( .A1(n699), .A2(n698), .ZN(n703) );
  NOR2_X1 U798 ( .A1(n970), .A2(n700), .ZN(n701) );
  XOR2_X1 U799 ( .A(n701), .B(KEYINPUT28), .Z(n702) );
  NAND2_X1 U800 ( .A1(n703), .A2(n702), .ZN(n705) );
  NAND2_X1 U801 ( .A1(n707), .A2(n706), .ZN(n719) );
  NOR2_X1 U802 ( .A1(G171), .A2(n708), .ZN(n715) );
  XNOR2_X1 U803 ( .A(KEYINPUT30), .B(n712), .ZN(n713) );
  NOR2_X1 U804 ( .A1(G168), .A2(n713), .ZN(n714) );
  NOR2_X1 U805 ( .A1(n715), .A2(n714), .ZN(n717) );
  NAND2_X1 U806 ( .A1(n719), .A2(n718), .ZN(n724) );
  NOR2_X1 U807 ( .A1(n720), .A2(n516), .ZN(n721) );
  NAND2_X1 U808 ( .A1(n722), .A2(n721), .ZN(n735) );
  AND2_X1 U809 ( .A1(G286), .A2(G8), .ZN(n723) );
  NAND2_X1 U810 ( .A1(n724), .A2(n723), .ZN(n732) );
  INV_X1 U811 ( .A(G8), .ZN(n730) );
  NOR2_X1 U812 ( .A1(G1971), .A2(n789), .ZN(n727) );
  NOR2_X1 U813 ( .A1(G2090), .A2(n725), .ZN(n726) );
  NOR2_X1 U814 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U815 ( .A1(n728), .A2(G303), .ZN(n729) );
  OR2_X1 U816 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U817 ( .A(KEYINPUT32), .B(n733), .ZN(n734) );
  NAND2_X1 U818 ( .A1(n735), .A2(n734), .ZN(n787) );
  NOR2_X1 U819 ( .A1(G1976), .A2(G288), .ZN(n743) );
  NOR2_X1 U820 ( .A1(G1971), .A2(G303), .ZN(n736) );
  NOR2_X1 U821 ( .A1(n743), .A2(n736), .ZN(n973) );
  INV_X1 U822 ( .A(KEYINPUT93), .ZN(n737) );
  XNOR2_X1 U823 ( .A(n515), .B(n737), .ZN(n741) );
  NAND2_X1 U824 ( .A1(G288), .A2(G1976), .ZN(n738) );
  XNOR2_X1 U825 ( .A(n738), .B(KEYINPUT94), .ZN(n974) );
  INV_X1 U826 ( .A(n974), .ZN(n739) );
  OR2_X1 U827 ( .A1(n739), .A2(n789), .ZN(n740) );
  NOR2_X1 U828 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U829 ( .A1(n742), .A2(KEYINPUT33), .ZN(n746) );
  NAND2_X1 U830 ( .A1(n743), .A2(KEYINPUT33), .ZN(n744) );
  NOR2_X1 U831 ( .A1(n789), .A2(n744), .ZN(n745) );
  NOR2_X1 U832 ( .A1(n746), .A2(n745), .ZN(n782) );
  XOR2_X1 U833 ( .A(G1981), .B(G305), .Z(n984) );
  XOR2_X1 U834 ( .A(G2067), .B(KEYINPUT37), .Z(n747) );
  XOR2_X1 U835 ( .A(KEYINPUT80), .B(n747), .Z(n800) );
  NAND2_X1 U836 ( .A1(G104), .A2(n880), .ZN(n749) );
  NAND2_X1 U837 ( .A1(G140), .A2(n881), .ZN(n748) );
  NAND2_X1 U838 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U839 ( .A(KEYINPUT34), .B(n750), .ZN(n756) );
  NAND2_X1 U840 ( .A1(G116), .A2(n884), .ZN(n752) );
  NAND2_X1 U841 ( .A1(G128), .A2(n885), .ZN(n751) );
  NAND2_X1 U842 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U843 ( .A(KEYINPUT81), .B(n753), .ZN(n754) );
  XNOR2_X1 U844 ( .A(KEYINPUT35), .B(n754), .ZN(n755) );
  NOR2_X1 U845 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U846 ( .A(KEYINPUT36), .B(n757), .ZN(n875) );
  NOR2_X1 U847 ( .A1(n800), .A2(n875), .ZN(n917) );
  NOR2_X1 U848 ( .A1(n759), .A2(n758), .ZN(n812) );
  NAND2_X1 U849 ( .A1(n917), .A2(n812), .ZN(n760) );
  XOR2_X1 U850 ( .A(KEYINPUT82), .B(n760), .Z(n808) );
  NAND2_X1 U851 ( .A1(G117), .A2(n884), .ZN(n762) );
  NAND2_X1 U852 ( .A1(G129), .A2(n885), .ZN(n761) );
  NAND2_X1 U853 ( .A1(n762), .A2(n761), .ZN(n765) );
  NAND2_X1 U854 ( .A1(n880), .A2(G105), .ZN(n763) );
  XOR2_X1 U855 ( .A(KEYINPUT38), .B(n763), .Z(n764) );
  NOR2_X1 U856 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U857 ( .A(n766), .B(KEYINPUT84), .ZN(n768) );
  NAND2_X1 U858 ( .A1(G141), .A2(n881), .ZN(n767) );
  NAND2_X1 U859 ( .A1(n768), .A2(n767), .ZN(n874) );
  NAND2_X1 U860 ( .A1(n874), .A2(G1996), .ZN(n777) );
  NAND2_X1 U861 ( .A1(G107), .A2(n884), .ZN(n770) );
  NAND2_X1 U862 ( .A1(G119), .A2(n885), .ZN(n769) );
  NAND2_X1 U863 ( .A1(n770), .A2(n769), .ZN(n773) );
  NAND2_X1 U864 ( .A1(G131), .A2(n881), .ZN(n771) );
  XNOR2_X1 U865 ( .A(KEYINPUT83), .B(n771), .ZN(n772) );
  NOR2_X1 U866 ( .A1(n773), .A2(n772), .ZN(n775) );
  NAND2_X1 U867 ( .A1(n880), .A2(G95), .ZN(n774) );
  NAND2_X1 U868 ( .A1(n775), .A2(n774), .ZN(n891) );
  NAND2_X1 U869 ( .A1(G1991), .A2(n891), .ZN(n776) );
  NAND2_X1 U870 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U871 ( .A(n778), .B(KEYINPUT85), .ZN(n922) );
  INV_X1 U872 ( .A(n812), .ZN(n779) );
  NOR2_X1 U873 ( .A1(n922), .A2(n779), .ZN(n803) );
  OR2_X1 U874 ( .A1(n808), .A2(n803), .ZN(n794) );
  INV_X1 U875 ( .A(n794), .ZN(n780) );
  AND2_X1 U876 ( .A1(n984), .A2(n780), .ZN(n781) );
  NAND2_X1 U877 ( .A1(n782), .A2(n781), .ZN(n796) );
  NOR2_X1 U878 ( .A1(G1981), .A2(G305), .ZN(n783) );
  XOR2_X1 U879 ( .A(n783), .B(KEYINPUT24), .Z(n784) );
  OR2_X1 U880 ( .A1(n789), .A2(n784), .ZN(n792) );
  NOR2_X1 U881 ( .A1(G2090), .A2(G303), .ZN(n785) );
  XOR2_X1 U882 ( .A(KEYINPUT95), .B(n785), .Z(n786) );
  NAND2_X1 U883 ( .A1(G8), .A2(n786), .ZN(n788) );
  NAND2_X1 U884 ( .A1(n788), .A2(n787), .ZN(n790) );
  NAND2_X1 U885 ( .A1(n790), .A2(n789), .ZN(n791) );
  AND2_X1 U886 ( .A1(n792), .A2(n791), .ZN(n793) );
  OR2_X1 U887 ( .A1(n794), .A2(n793), .ZN(n795) );
  NAND2_X1 U888 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U889 ( .A(n797), .B(KEYINPUT96), .ZN(n799) );
  XNOR2_X1 U890 ( .A(G1986), .B(G290), .ZN(n968) );
  NAND2_X1 U891 ( .A1(n968), .A2(n812), .ZN(n798) );
  NAND2_X1 U892 ( .A1(n799), .A2(n798), .ZN(n815) );
  AND2_X1 U893 ( .A1(n875), .A2(n800), .ZN(n920) );
  NOR2_X1 U894 ( .A1(G1996), .A2(n874), .ZN(n924) );
  NOR2_X1 U895 ( .A1(G1986), .A2(G290), .ZN(n801) );
  NOR2_X1 U896 ( .A1(G1991), .A2(n891), .ZN(n913) );
  NOR2_X1 U897 ( .A1(n801), .A2(n913), .ZN(n802) );
  NOR2_X1 U898 ( .A1(n803), .A2(n802), .ZN(n804) );
  XOR2_X1 U899 ( .A(KEYINPUT97), .B(n804), .Z(n805) );
  NOR2_X1 U900 ( .A1(n924), .A2(n805), .ZN(n806) );
  XOR2_X1 U901 ( .A(KEYINPUT39), .B(n806), .Z(n807) );
  NOR2_X1 U902 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U903 ( .A(n809), .B(KEYINPUT98), .ZN(n810) );
  NOR2_X1 U904 ( .A1(n920), .A2(n810), .ZN(n811) );
  XNOR2_X1 U905 ( .A(KEYINPUT99), .B(n811), .ZN(n813) );
  NAND2_X1 U906 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U907 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U908 ( .A(n816), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U909 ( .A(G2454), .B(G2446), .ZN(n825) );
  XNOR2_X1 U910 ( .A(G2430), .B(G2443), .ZN(n823) );
  XOR2_X1 U911 ( .A(G2435), .B(KEYINPUT100), .Z(n818) );
  XNOR2_X1 U912 ( .A(G2451), .B(G2438), .ZN(n817) );
  XNOR2_X1 U913 ( .A(n818), .B(n817), .ZN(n819) );
  XOR2_X1 U914 ( .A(n819), .B(G2427), .Z(n821) );
  XNOR2_X1 U915 ( .A(G1341), .B(G1348), .ZN(n820) );
  XNOR2_X1 U916 ( .A(n821), .B(n820), .ZN(n822) );
  XNOR2_X1 U917 ( .A(n823), .B(n822), .ZN(n824) );
  XNOR2_X1 U918 ( .A(n825), .B(n824), .ZN(n826) );
  NAND2_X1 U919 ( .A1(n826), .A2(G14), .ZN(n905) );
  XNOR2_X1 U920 ( .A(KEYINPUT101), .B(n905), .ZN(G401) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n911), .ZN(G217) );
  NAND2_X1 U922 ( .A1(G15), .A2(G2), .ZN(n827) );
  XOR2_X1 U923 ( .A(KEYINPUT102), .B(n827), .Z(n828) );
  NAND2_X1 U924 ( .A1(G661), .A2(n828), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n829) );
  NAND2_X1 U926 ( .A1(n830), .A2(n829), .ZN(G188) );
  INV_X1 U928 ( .A(G120), .ZN(G236) );
  INV_X1 U929 ( .A(G96), .ZN(G221) );
  INV_X1 U930 ( .A(G69), .ZN(G235) );
  NOR2_X1 U931 ( .A1(n832), .A2(n831), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U933 ( .A(KEYINPUT103), .B(n833), .ZN(G319) );
  XOR2_X1 U934 ( .A(G2100), .B(G2096), .Z(n835) );
  XNOR2_X1 U935 ( .A(KEYINPUT42), .B(G2678), .ZN(n834) );
  XNOR2_X1 U936 ( .A(n835), .B(n834), .ZN(n839) );
  XOR2_X1 U937 ( .A(KEYINPUT43), .B(G2090), .Z(n837) );
  XNOR2_X1 U938 ( .A(G2067), .B(G2072), .ZN(n836) );
  XNOR2_X1 U939 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U940 ( .A(n839), .B(n838), .Z(n841) );
  XNOR2_X1 U941 ( .A(G2084), .B(G2078), .ZN(n840) );
  XNOR2_X1 U942 ( .A(n841), .B(n840), .ZN(G227) );
  XOR2_X1 U943 ( .A(KEYINPUT41), .B(KEYINPUT106), .Z(n843) );
  XNOR2_X1 U944 ( .A(KEYINPUT105), .B(G2474), .ZN(n842) );
  XNOR2_X1 U945 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U946 ( .A(n844), .B(KEYINPUT107), .Z(n846) );
  XNOR2_X1 U947 ( .A(G1996), .B(G1991), .ZN(n845) );
  XNOR2_X1 U948 ( .A(n846), .B(n845), .ZN(n854) );
  XNOR2_X1 U949 ( .A(G1971), .B(n969), .ZN(n848) );
  XNOR2_X1 U950 ( .A(G1986), .B(G1961), .ZN(n847) );
  XNOR2_X1 U951 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U952 ( .A(KEYINPUT104), .B(G1976), .Z(n850) );
  XNOR2_X1 U953 ( .A(G1966), .B(G1981), .ZN(n849) );
  XNOR2_X1 U954 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U955 ( .A(n852), .B(n851), .Z(n853) );
  XNOR2_X1 U956 ( .A(n854), .B(n853), .ZN(G229) );
  NAND2_X1 U957 ( .A1(G124), .A2(n885), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n855), .B(KEYINPUT44), .ZN(n857) );
  NAND2_X1 U959 ( .A1(n884), .A2(G112), .ZN(n856) );
  NAND2_X1 U960 ( .A1(n857), .A2(n856), .ZN(n861) );
  NAND2_X1 U961 ( .A1(G100), .A2(n880), .ZN(n859) );
  NAND2_X1 U962 ( .A1(G136), .A2(n881), .ZN(n858) );
  NAND2_X1 U963 ( .A1(n859), .A2(n858), .ZN(n860) );
  NOR2_X1 U964 ( .A1(n861), .A2(n860), .ZN(G162) );
  XOR2_X1 U965 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n862) );
  XNOR2_X1 U966 ( .A(n914), .B(n862), .ZN(n863) );
  XOR2_X1 U967 ( .A(n863), .B(KEYINPUT109), .Z(n865) );
  XNOR2_X1 U968 ( .A(G164), .B(KEYINPUT110), .ZN(n864) );
  XNOR2_X1 U969 ( .A(n865), .B(n864), .ZN(n895) );
  NAND2_X1 U970 ( .A1(G106), .A2(n880), .ZN(n867) );
  NAND2_X1 U971 ( .A1(G142), .A2(n881), .ZN(n866) );
  NAND2_X1 U972 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U973 ( .A(n868), .B(KEYINPUT45), .ZN(n870) );
  NAND2_X1 U974 ( .A1(G118), .A2(n884), .ZN(n869) );
  NAND2_X1 U975 ( .A1(n870), .A2(n869), .ZN(n873) );
  NAND2_X1 U976 ( .A1(n885), .A2(G130), .ZN(n871) );
  XOR2_X1 U977 ( .A(KEYINPUT108), .B(n871), .Z(n872) );
  NOR2_X1 U978 ( .A1(n873), .A2(n872), .ZN(n879) );
  XNOR2_X1 U979 ( .A(n874), .B(G162), .ZN(n877) );
  XOR2_X1 U980 ( .A(G160), .B(n875), .Z(n876) );
  XNOR2_X1 U981 ( .A(n877), .B(n876), .ZN(n878) );
  XNOR2_X1 U982 ( .A(n879), .B(n878), .ZN(n893) );
  NAND2_X1 U983 ( .A1(G103), .A2(n880), .ZN(n883) );
  NAND2_X1 U984 ( .A1(G139), .A2(n881), .ZN(n882) );
  NAND2_X1 U985 ( .A1(n883), .A2(n882), .ZN(n890) );
  NAND2_X1 U986 ( .A1(G115), .A2(n884), .ZN(n887) );
  NAND2_X1 U987 ( .A1(G127), .A2(n885), .ZN(n886) );
  NAND2_X1 U988 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U989 ( .A(KEYINPUT47), .B(n888), .Z(n889) );
  NOR2_X1 U990 ( .A1(n890), .A2(n889), .ZN(n929) );
  XNOR2_X1 U991 ( .A(n891), .B(n929), .ZN(n892) );
  XNOR2_X1 U992 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U993 ( .A(n895), .B(n894), .Z(n896) );
  NOR2_X1 U994 ( .A1(G37), .A2(n896), .ZN(G395) );
  XOR2_X1 U995 ( .A(KEYINPUT111), .B(n897), .Z(n900) );
  XOR2_X1 U996 ( .A(n898), .B(G286), .Z(n899) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n902) );
  XOR2_X1 U998 ( .A(n983), .B(G301), .Z(n901) );
  XNOR2_X1 U999 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n903), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(KEYINPUT112), .B(n904), .ZN(G397) );
  NAND2_X1 U1002 ( .A1(G319), .A2(n905), .ZN(n908) );
  NOR2_X1 U1003 ( .A1(G227), .A2(G229), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(KEYINPUT49), .B(n906), .ZN(n907) );
  NOR2_X1 U1005 ( .A1(n908), .A2(n907), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(G395), .A2(G397), .ZN(n909) );
  NAND2_X1 U1007 ( .A1(n910), .A2(n909), .ZN(G225) );
  INV_X1 U1008 ( .A(G225), .ZN(G308) );
  INV_X1 U1009 ( .A(G108), .ZN(G238) );
  INV_X1 U1010 ( .A(n911), .ZN(G223) );
  XOR2_X1 U1011 ( .A(G160), .B(G2084), .Z(n912) );
  NOR2_X1 U1012 ( .A1(n913), .A2(n912), .ZN(n915) );
  NAND2_X1 U1013 ( .A1(n915), .A2(n914), .ZN(n916) );
  NOR2_X1 U1014 ( .A1(n917), .A2(n916), .ZN(n918) );
  XNOR2_X1 U1015 ( .A(KEYINPUT113), .B(n918), .ZN(n919) );
  NOR2_X1 U1016 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1017 ( .A1(n922), .A2(n921), .ZN(n927) );
  XOR2_X1 U1018 ( .A(G2090), .B(G162), .Z(n923) );
  NOR2_X1 U1019 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1020 ( .A(n925), .B(KEYINPUT51), .ZN(n926) );
  NOR2_X1 U1021 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1022 ( .A(KEYINPUT114), .B(n928), .Z(n936) );
  XNOR2_X1 U1023 ( .A(G164), .B(G2078), .ZN(n932) );
  XOR2_X1 U1024 ( .A(G2072), .B(n929), .Z(n930) );
  XNOR2_X1 U1025 ( .A(KEYINPUT115), .B(n930), .ZN(n931) );
  NAND2_X1 U1026 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1027 ( .A(n933), .B(KEYINPUT50), .ZN(n934) );
  XNOR2_X1 U1028 ( .A(KEYINPUT116), .B(n934), .ZN(n935) );
  NOR2_X1 U1029 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1030 ( .A(KEYINPUT52), .B(n937), .ZN(n938) );
  INV_X1 U1031 ( .A(KEYINPUT55), .ZN(n941) );
  NAND2_X1 U1032 ( .A1(n938), .A2(n941), .ZN(n939) );
  NAND2_X1 U1033 ( .A1(n939), .A2(G29), .ZN(n940) );
  XOR2_X1 U1034 ( .A(KEYINPUT117), .B(n940), .Z(n1026) );
  XNOR2_X1 U1035 ( .A(n941), .B(KEYINPUT120), .ZN(n962) );
  XNOR2_X1 U1036 ( .A(G2090), .B(G35), .ZN(n957) );
  XNOR2_X1 U1037 ( .A(G2067), .B(G26), .ZN(n943) );
  XNOR2_X1 U1038 ( .A(G33), .B(G2072), .ZN(n942) );
  NOR2_X1 U1039 ( .A1(n943), .A2(n942), .ZN(n953) );
  XOR2_X1 U1040 ( .A(G1991), .B(G25), .Z(n944) );
  NAND2_X1 U1041 ( .A1(n944), .A2(G28), .ZN(n951) );
  XOR2_X1 U1042 ( .A(n945), .B(G27), .Z(n948) );
  XNOR2_X1 U1043 ( .A(n946), .B(G32), .ZN(n947) );
  NAND2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1045 ( .A(KEYINPUT118), .B(n949), .ZN(n950) );
  NOR2_X1 U1046 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(KEYINPUT53), .B(n954), .ZN(n955) );
  XNOR2_X1 U1049 ( .A(n955), .B(KEYINPUT119), .ZN(n956) );
  NOR2_X1 U1050 ( .A1(n957), .A2(n956), .ZN(n960) );
  XOR2_X1 U1051 ( .A(G2084), .B(G34), .Z(n958) );
  XNOR2_X1 U1052 ( .A(KEYINPUT54), .B(n958), .ZN(n959) );
  NAND2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1054 ( .A(n962), .B(n961), .ZN(n964) );
  INV_X1 U1055 ( .A(G29), .ZN(n963) );
  NAND2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1057 ( .A1(G11), .A2(n965), .ZN(n1024) );
  INV_X1 U1058 ( .A(G16), .ZN(n1020) );
  XOR2_X1 U1059 ( .A(n1020), .B(KEYINPUT56), .Z(n993) );
  XOR2_X1 U1060 ( .A(G1348), .B(n966), .Z(n967) );
  NOR2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n981) );
  XOR2_X1 U1062 ( .A(n970), .B(n969), .Z(n972) );
  XOR2_X1 U1063 ( .A(G301), .B(G1961), .Z(n971) );
  NAND2_X1 U1064 ( .A1(n972), .A2(n971), .ZN(n979) );
  NAND2_X1 U1065 ( .A1(n974), .A2(n973), .ZN(n976) );
  AND2_X1 U1066 ( .A1(G303), .A2(G1971), .ZN(n975) );
  NOR2_X1 U1067 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1068 ( .A(KEYINPUT122), .B(n977), .Z(n978) );
  NOR2_X1 U1069 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1070 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1071 ( .A(KEYINPUT123), .B(n982), .ZN(n991) );
  XNOR2_X1 U1072 ( .A(n983), .B(G1341), .ZN(n989) );
  XNOR2_X1 U1073 ( .A(G1966), .B(G168), .ZN(n985) );
  NAND2_X1 U1074 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1075 ( .A(n986), .B(KEYINPUT57), .ZN(n987) );
  XNOR2_X1 U1076 ( .A(KEYINPUT121), .B(n987), .ZN(n988) );
  NOR2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1078 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1079 ( .A1(n993), .A2(n992), .ZN(n1022) );
  XNOR2_X1 U1080 ( .A(n994), .B(G5), .ZN(n1016) );
  XOR2_X1 U1081 ( .A(G20), .B(G1956), .Z(n998) );
  XNOR2_X1 U1082 ( .A(G1341), .B(G19), .ZN(n996) );
  XNOR2_X1 U1083 ( .A(G1981), .B(G6), .ZN(n995) );
  NOR2_X1 U1084 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1085 ( .A1(n998), .A2(n997), .ZN(n1001) );
  XOR2_X1 U1086 ( .A(KEYINPUT59), .B(G1348), .Z(n999) );
  XNOR2_X1 U1087 ( .A(G4), .B(n999), .ZN(n1000) );
  NOR2_X1 U1088 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1089 ( .A(KEYINPUT124), .B(n1002), .ZN(n1003) );
  XNOR2_X1 U1090 ( .A(n1003), .B(KEYINPUT60), .ZN(n1011) );
  XOR2_X1 U1091 ( .A(G1976), .B(KEYINPUT126), .Z(n1004) );
  XNOR2_X1 U1092 ( .A(G23), .B(n1004), .ZN(n1008) );
  XNOR2_X1 U1093 ( .A(G1986), .B(G24), .ZN(n1006) );
  XNOR2_X1 U1094 ( .A(G1971), .B(G22), .ZN(n1005) );
  NOR2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1097 ( .A(KEYINPUT58), .B(n1009), .Z(n1010) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1014) );
  XOR2_X1 U1099 ( .A(KEYINPUT125), .B(G1966), .Z(n1012) );
  XNOR2_X1 U1100 ( .A(G21), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1103 ( .A(n1017), .B(KEYINPUT61), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(KEYINPUT127), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1107 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1108 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1027), .ZN(G150) );
  INV_X1 U1110 ( .A(G150), .ZN(G311) );
  INV_X1 U1111 ( .A(G303), .ZN(G166) );
endmodule

