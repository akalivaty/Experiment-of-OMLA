//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 1 0 1 1 0 1 0 0 0 1 1 0 0 1 0 1 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 1 0 0 1 0 1 0 0 1 0 0 0 1 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n789, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n989, new_n990, new_n991,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1018, new_n1019;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(G183gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT27), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT27), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G183gat), .ZN(new_n207));
  INV_X1    g006(.A(G190gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT28), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT27), .B(G183gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n212), .A2(KEYINPUT28), .A3(new_n208), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT26), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NOR3_X1   g018(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n214), .A2(new_n215), .A3(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G169gat), .ZN(new_n223));
  INV_X1    g022(.A(G176gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT23), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(new_n226), .A3(new_n216), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n226), .B1(new_n225), .B2(new_n216), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT23), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n231), .B1(G169gat), .B2(G176gat), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n232), .A2(KEYINPUT25), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n204), .A2(new_n208), .ZN(new_n234));
  NAND3_X1  g033(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n234), .B(new_n235), .C1(new_n236), .C2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT24), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n215), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n240), .A2(KEYINPUT67), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n233), .B1(new_n238), .B2(new_n241), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n230), .A2(new_n242), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT65), .A4(KEYINPUT23), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n244), .A2(new_n216), .A3(new_n232), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT65), .B1(new_n217), .B2(KEYINPUT23), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AND2_X1   g046(.A1(new_n234), .A2(new_n235), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n236), .A2(KEYINPUT64), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT64), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n240), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n248), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT25), .B1(new_n247), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n222), .B1(new_n243), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT29), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n203), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n257));
  OR2_X1    g056(.A1(G197gat), .A2(G204gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(G197gat), .A2(G204gat), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(G211gat), .B(G218gat), .Z(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n263), .B1(new_n260), .B2(new_n261), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n215), .B1(new_n219), .B2(new_n220), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n269), .B1(new_n211), .B2(new_n213), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT25), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n234), .B(new_n235), .C1(new_n236), .C2(KEYINPUT64), .ZN(new_n272));
  INV_X1    g071(.A(new_n249), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT65), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n225), .A2(new_n275), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n276), .A2(new_n244), .A3(new_n216), .A4(new_n232), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n271), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  NOR3_X1   g077(.A1(new_n231), .A2(G169gat), .A3(G176gat), .ZN(new_n279));
  INV_X1    g078(.A(new_n216), .ZN(new_n280));
  OAI21_X1  g079(.A(KEYINPUT66), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(new_n227), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n236), .A2(new_n237), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n240), .A2(KEYINPUT67), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n248), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n282), .A2(new_n285), .A3(new_n233), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n270), .B1(new_n278), .B2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n202), .B(KEYINPUT71), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n268), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(KEYINPUT72), .B1(new_n256), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n288), .B1(new_n254), .B2(new_n255), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n287), .A2(new_n202), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n267), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G8gat), .B(G36gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(G64gat), .B(G92gat), .ZN(new_n296));
  XOR2_X1   g095(.A(new_n295), .B(new_n296), .Z(new_n297));
  OAI21_X1  g096(.A(new_n202), .B1(new_n287), .B2(KEYINPUT29), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n254), .A2(new_n288), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT72), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n298), .A2(new_n299), .A3(new_n300), .A4(new_n268), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n291), .A2(new_n294), .A3(new_n297), .A4(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT30), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n291), .A2(new_n294), .A3(new_n301), .ZN(new_n305));
  INV_X1    g104(.A(new_n297), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n303), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n291), .A2(new_n294), .A3(new_n301), .A4(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n304), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT80), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT80), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n304), .A2(new_n307), .A3(new_n312), .A4(new_n309), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT39), .ZN(new_n314));
  NAND2_X1  g113(.A1(G225gat), .A2(G233gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G113gat), .B(G120gat), .ZN(new_n317));
  OR2_X1    g116(.A1(new_n317), .A2(KEYINPUT1), .ZN(new_n318));
  INV_X1    g117(.A(G134gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G127gat), .ZN(new_n320));
  INV_X1    g119(.A(G127gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(G134gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT1), .ZN(new_n324));
  INV_X1    g123(.A(G120gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n325), .A2(KEYINPUT68), .A3(G113gat), .ZN(new_n326));
  AND4_X1   g125(.A1(new_n324), .A2(new_n326), .A3(new_n320), .A4(new_n322), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT68), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n317), .A2(new_n328), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n318), .A2(new_n323), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G141gat), .A2(G148gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(G141gat), .A2(G148gat), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n332), .A2(new_n333), .A3(KEYINPUT2), .ZN(new_n334));
  XNOR2_X1  g133(.A(G155gat), .B(G162gat), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT73), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(G141gat), .ZN(new_n337));
  INV_X1    g136(.A(G148gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT2), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n339), .A2(new_n340), .A3(new_n331), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT73), .ZN(new_n342));
  INV_X1    g141(.A(G162gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(G155gat), .ZN(new_n344));
  INV_X1    g143(.A(G155gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(G162gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n341), .A2(new_n342), .A3(new_n347), .ZN(new_n348));
  NOR3_X1   g147(.A1(new_n347), .A2(new_n333), .A3(new_n332), .ZN(new_n349));
  XNOR2_X1  g148(.A(KEYINPUT74), .B(G162gat), .ZN(new_n350));
  OAI21_X1  g149(.A(KEYINPUT2), .B1(new_n350), .B2(new_n345), .ZN(new_n351));
  AOI22_X1  g150(.A1(new_n336), .A2(new_n348), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT3), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n330), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n332), .A2(new_n333), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n343), .A2(KEYINPUT74), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT74), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(G162gat), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n345), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n355), .B(new_n335), .C1(new_n359), .C2(new_n340), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n341), .A2(new_n342), .A3(new_n347), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n342), .B1(new_n341), .B2(new_n347), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT3), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT75), .B1(new_n354), .B2(new_n364), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n360), .B(new_n353), .C1(new_n361), .C2(new_n362), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n327), .A2(new_n329), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n323), .B1(new_n317), .B2(KEYINPUT1), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n336), .A2(new_n348), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n353), .B1(new_n371), .B2(new_n360), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT75), .ZN(new_n373));
  NOR3_X1   g172(.A1(new_n370), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n365), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT4), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n376), .B1(new_n363), .B2(new_n369), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n352), .A2(KEYINPUT4), .A3(new_n330), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n314), .B(new_n316), .C1(new_n375), .C2(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n352), .A2(new_n330), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n363), .A2(new_n369), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n314), .B1(new_n383), .B2(new_n315), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n354), .A2(KEYINPUT75), .A3(new_n364), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n373), .B1(new_n370), .B2(new_n372), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n379), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n384), .B1(new_n387), .B2(new_n315), .ZN(new_n388));
  XNOR2_X1  g187(.A(G1gat), .B(G29gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n389), .B(KEYINPUT0), .ZN(new_n390));
  XNOR2_X1  g189(.A(G57gat), .B(G85gat), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n390), .B(new_n391), .Z(new_n392));
  NAND3_X1  g191(.A1(new_n380), .A2(new_n388), .A3(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT40), .ZN(new_n394));
  OR2_X1    g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AND3_X1   g194(.A1(new_n377), .A2(new_n378), .A3(new_n315), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n396), .B1(new_n365), .B2(new_n374), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n316), .B1(new_n381), .B2(new_n382), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT76), .B1(new_n398), .B2(KEYINPUT5), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n352), .A2(new_n330), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n363), .A2(new_n369), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n315), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT76), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT5), .ZN(new_n404));
  NOR3_X1   g203(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n397), .B1(new_n399), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n385), .A2(new_n386), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(new_n404), .A3(new_n396), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n392), .ZN(new_n410));
  AOI22_X1  g209(.A1(new_n393), .A2(new_n394), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n311), .A2(new_n313), .A3(new_n395), .A4(new_n411), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n260), .A2(new_n263), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n260), .A2(new_n263), .ZN(new_n414));
  NOR3_X1   g213(.A1(new_n413), .A2(new_n414), .A3(KEYINPUT29), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n363), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n416), .A2(KEYINPUT77), .A3(new_n364), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT77), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n418), .B(new_n363), .C1(new_n415), .C2(KEYINPUT3), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n268), .B1(new_n255), .B2(new_n366), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n417), .B(new_n419), .C1(new_n420), .C2(KEYINPUT78), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n420), .A2(KEYINPUT78), .ZN(new_n422));
  INV_X1    g221(.A(G228gat), .ZN(new_n423));
  INV_X1    g222(.A(G233gat), .ZN(new_n424));
  OAI22_X1  g223(.A1(new_n421), .A2(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(G78gat), .B(G106gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT31), .B(G50gat), .ZN(new_n427));
  XOR2_X1   g226(.A(new_n426), .B(new_n427), .Z(new_n428));
  NOR2_X1   g227(.A1(new_n428), .A2(KEYINPUT79), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n353), .B1(new_n267), .B2(KEYINPUT29), .ZN(new_n430));
  AOI211_X1 g229(.A(new_n423), .B(new_n424), .C1(new_n430), .C2(new_n363), .ZN(new_n431));
  INV_X1    g230(.A(new_n420), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n429), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n425), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n428), .A2(KEYINPUT79), .ZN(new_n435));
  INV_X1    g234(.A(G22gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n435), .B(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n434), .B(new_n437), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n305), .A2(KEYINPUT37), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n306), .B1(new_n305), .B2(KEYINPUT37), .ZN(new_n440));
  OAI21_X1  g239(.A(KEYINPUT38), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n409), .A2(KEYINPUT6), .A3(new_n410), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n398), .A2(KEYINPUT76), .A3(KEYINPUT5), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n403), .B1(new_n402), .B2(new_n404), .ZN(new_n444));
  AOI22_X1  g243(.A1(new_n443), .A2(new_n444), .B1(new_n407), .B2(new_n396), .ZN(new_n445));
  INV_X1    g244(.A(new_n408), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n410), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT6), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n406), .A2(new_n392), .A3(new_n408), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n441), .A2(new_n442), .A3(new_n450), .A4(new_n302), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT37), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n287), .A2(new_n289), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n267), .B1(new_n256), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT81), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n292), .A2(new_n293), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n454), .A2(new_n455), .B1(new_n456), .B2(new_n268), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n268), .B1(new_n298), .B2(new_n299), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT81), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n452), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT38), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n461), .B(new_n306), .C1(new_n305), .C2(KEYINPUT37), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT82), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n306), .A2(KEYINPUT37), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n307), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT82), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n289), .B1(new_n287), .B2(KEYINPUT29), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n467), .B1(new_n287), .B2(new_n202), .ZN(new_n468));
  OAI22_X1  g267(.A1(new_n458), .A2(KEYINPUT81), .B1(new_n468), .B2(new_n267), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n454), .A2(new_n455), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT37), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n465), .A2(new_n466), .A3(new_n471), .A4(new_n461), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n463), .A2(new_n472), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n412), .B(new_n438), .C1(new_n451), .C2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n450), .A2(new_n442), .ZN(new_n475));
  INV_X1    g274(.A(new_n310), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n437), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n434), .B(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(G227gat), .A2(G233gat), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  AOI211_X1 g281(.A(new_n270), .B(new_n369), .C1(new_n278), .C2(new_n286), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n278), .A2(new_n286), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n330), .B1(new_n484), .B2(new_n222), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n482), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT32), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT33), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  XOR2_X1   g288(.A(G15gat), .B(G43gat), .Z(new_n490));
  XNOR2_X1  g289(.A(G71gat), .B(G99gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n490), .B(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n487), .A2(new_n489), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n254), .A2(new_n369), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n287), .A2(new_n330), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n494), .A2(new_n495), .A3(new_n481), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT34), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n496), .B(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n492), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n486), .B(KEYINPUT32), .C1(new_n488), .C2(new_n499), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n493), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n498), .B1(new_n493), .B2(new_n500), .ZN(new_n502));
  NOR3_X1   g301(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT36), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n493), .A2(new_n500), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT69), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n505), .B1(new_n501), .B2(new_n502), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(KEYINPUT69), .A3(new_n498), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n503), .B1(new_n508), .B2(KEYINPUT36), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n474), .A2(new_n480), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n506), .A2(new_n438), .A3(new_n507), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT35), .B1(new_n511), .B2(new_n477), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n479), .A2(KEYINPUT35), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n311), .A2(new_n313), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n501), .A2(new_n502), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n513), .A2(new_n475), .A3(new_n514), .A4(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n510), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(G232gat), .A2(G233gat), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n520), .A2(KEYINPUT41), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(KEYINPUT88), .ZN(new_n522));
  XNOR2_X1  g321(.A(G134gat), .B(G162gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n522), .B(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n520), .A2(KEYINPUT41), .ZN(new_n526));
  XNOR2_X1  g325(.A(G43gat), .B(G50gat), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n527), .A2(KEYINPUT15), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(KEYINPUT15), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT14), .ZN(new_n530));
  INV_X1    g329(.A(G29gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n533));
  AOI21_X1  g332(.A(G36gat), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(G36gat), .ZN(new_n535));
  NOR3_X1   g334(.A1(new_n530), .A2(new_n535), .A3(G29gat), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n528), .B(new_n529), .C1(new_n534), .C2(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n534), .A2(new_n536), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n538), .A2(KEYINPUT15), .A3(new_n527), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G85gat), .A2(G92gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(KEYINPUT7), .ZN(new_n543));
  NAND2_X1  g342(.A1(G99gat), .A2(G106gat), .ZN(new_n544));
  INV_X1    g343(.A(G85gat), .ZN(new_n545));
  INV_X1    g344(.A(G92gat), .ZN(new_n546));
  AOI22_X1  g345(.A1(KEYINPUT8), .A2(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(G99gat), .B(G106gat), .Z(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n549), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n551), .A2(new_n543), .A3(new_n547), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n526), .B1(new_n541), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT90), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT90), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n556), .B(new_n526), .C1(new_n541), .C2(new_n553), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT91), .ZN(new_n558));
  XNOR2_X1  g357(.A(G190gat), .B(G218gat), .ZN(new_n559));
  AOI22_X1  g358(.A1(new_n555), .A2(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT17), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n540), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n537), .A2(KEYINPUT17), .A3(new_n539), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(new_n563), .A3(new_n553), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT89), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n559), .A2(new_n558), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(KEYINPUT92), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n560), .A2(new_n565), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n568), .B1(new_n560), .B2(new_n565), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n525), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n560), .A2(new_n565), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(new_n567), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n574), .A2(new_n524), .A3(new_n569), .ZN(new_n575));
  AND2_X1   g374(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(G71gat), .B(G78gat), .Z(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT9), .ZN(new_n579));
  INV_X1    g378(.A(G71gat), .ZN(new_n580));
  INV_X1    g379(.A(G78gat), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(G57gat), .B(G64gat), .Z(new_n583));
  NAND3_X1  g382(.A1(new_n578), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n582), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(new_n577), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT21), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G231gat), .A2(G233gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(new_n321), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n436), .A2(G15gat), .ZN(new_n593));
  INV_X1    g392(.A(G15gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(G22gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT16), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n597), .A2(G1gat), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G15gat), .B(G22gat), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n600), .A2(G1gat), .ZN(new_n601));
  OAI21_X1  g400(.A(G8gat), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT84), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT84), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n604), .B(G8gat), .C1(new_n599), .C2(new_n601), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n600), .A2(G1gat), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n600), .B(KEYINPUT85), .C1(new_n597), .C2(G1gat), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT85), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n608), .B1(new_n596), .B2(new_n598), .ZN(new_n609));
  INV_X1    g408(.A(G8gat), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n606), .A2(new_n607), .A3(new_n609), .A4(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n603), .A2(new_n605), .A3(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n587), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n612), .B1(KEYINPUT21), .B2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n592), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(new_n345), .ZN(new_n617));
  XNOR2_X1  g416(.A(G183gat), .B(G211gat), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n617), .B(new_n618), .Z(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n615), .A2(new_n620), .ZN(new_n621));
  OR2_X1    g420(.A1(new_n592), .A2(new_n614), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n592), .A2(new_n614), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n622), .A2(new_n623), .A3(new_n619), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G230gat), .A2(G233gat), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n553), .A2(new_n587), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT10), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT93), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n550), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n551), .A2(new_n630), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n584), .A2(new_n552), .A3(new_n586), .A4(new_n632), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n628), .B(new_n629), .C1(new_n631), .C2(new_n633), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n613), .A2(KEYINPUT10), .A3(new_n552), .A4(new_n550), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n627), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n628), .B1(new_n631), .B2(new_n633), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n636), .B1(new_n627), .B2(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(G120gat), .B(G148gat), .Z(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT94), .ZN(new_n640));
  XNOR2_X1  g439(.A(G176gat), .B(G204gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n634), .A2(new_n635), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(new_n626), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n637), .A2(new_n627), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n645), .A2(new_n646), .A3(new_n642), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n576), .A2(new_n625), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n612), .A2(new_n540), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT87), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n653), .B1(new_n612), .B2(new_n540), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(G229gat), .A2(G233gat), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n656), .B(KEYINPUT13), .Z(new_n657));
  NAND2_X1  g456(.A1(new_n652), .A2(new_n654), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n655), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n612), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n660), .A2(new_n563), .A3(new_n562), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n661), .A2(new_n656), .A3(new_n651), .ZN(new_n662));
  AND3_X1   g461(.A1(new_n662), .A2(KEYINPUT86), .A3(KEYINPUT18), .ZN(new_n663));
  AOI21_X1  g462(.A(KEYINPUT18), .B1(new_n662), .B2(KEYINPUT86), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n659), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(G113gat), .B(G141gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(G197gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT11), .B(G169gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT83), .B(KEYINPUT12), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n665), .A2(new_n672), .ZN(new_n673));
  OAI211_X1 g472(.A(new_n659), .B(new_n671), .C1(new_n663), .C2(new_n664), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n650), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n518), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n678), .A2(new_n475), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT95), .B(G1gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1324gat));
  XNOR2_X1  g480(.A(KEYINPUT16), .B(G8gat), .ZN(new_n682));
  NOR2_X1   g481(.A1(KEYINPUT97), .A2(KEYINPUT42), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n678), .A2(new_n514), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT42), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT96), .ZN(new_n688));
  OAI22_X1  g487(.A1(new_n685), .A2(new_n688), .B1(new_n686), .B2(G8gat), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n678), .A2(KEYINPUT96), .A3(new_n514), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n687), .B1(new_n689), .B2(new_n690), .ZN(G1325gat));
  OAI21_X1  g490(.A(G15gat), .B1(new_n678), .B2(new_n509), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n515), .A2(new_n594), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n692), .B1(new_n678), .B2(new_n693), .ZN(G1326gat));
  NOR2_X1   g493(.A1(new_n678), .A2(new_n438), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT98), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT43), .B(G22gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1327gat));
  AOI21_X1  g497(.A(new_n576), .B1(new_n510), .B2(new_n517), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n676), .A2(new_n625), .A3(new_n648), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n475), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n701), .A2(new_n531), .A3(new_n702), .ZN(new_n703));
  XOR2_X1   g502(.A(KEYINPUT99), .B(KEYINPUT45), .Z(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n477), .A2(KEYINPUT100), .A3(new_n479), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT100), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n310), .B1(new_n450), .B2(new_n442), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n707), .B1(new_n708), .B2(new_n438), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n474), .A2(new_n509), .A3(new_n706), .A4(new_n709), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n710), .A2(new_n517), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n572), .A2(new_n575), .ZN(new_n712));
  XNOR2_X1  g511(.A(KEYINPUT101), .B(KEYINPUT44), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n715));
  OAI22_X1  g514(.A1(new_n711), .A2(new_n714), .B1(new_n699), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n700), .ZN(new_n717));
  OAI21_X1  g516(.A(G29gat), .B1(new_n717), .B2(new_n475), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n705), .A2(new_n718), .ZN(G1328gat));
  INV_X1    g518(.A(new_n514), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n701), .A2(new_n535), .A3(new_n720), .ZN(new_n721));
  XOR2_X1   g520(.A(KEYINPUT102), .B(KEYINPUT46), .Z(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(G36gat), .B1(new_n717), .B2(new_n514), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(G1329gat));
  NAND2_X1  g524(.A1(new_n699), .A2(new_n700), .ZN(new_n726));
  INV_X1    g525(.A(new_n515), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n726), .A2(G43gat), .A3(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT47), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n509), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n716), .A2(new_n731), .A3(new_n700), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT103), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(G43gat), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n732), .A2(new_n733), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n730), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n732), .A2(G43gat), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n729), .B1(new_n738), .B2(new_n728), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(G1330gat));
  INV_X1    g539(.A(KEYINPUT48), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n715), .B1(new_n518), .B2(new_n712), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n714), .B1(new_n710), .B2(new_n517), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n479), .B(new_n700), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n744), .A2(G50gat), .ZN(new_n745));
  INV_X1    g544(.A(G50gat), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n699), .A2(new_n746), .A3(new_n479), .A4(new_n700), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n741), .B1(new_n745), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(KEYINPUT48), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n746), .B1(new_n744), .B2(KEYINPUT104), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT104), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n716), .A2(new_n752), .A3(new_n479), .A4(new_n700), .ZN(new_n753));
  AOI211_X1 g552(.A(KEYINPUT105), .B(new_n750), .C1(new_n751), .C2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT105), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n744), .A2(KEYINPUT104), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n756), .A2(G50gat), .A3(new_n753), .ZN(new_n757));
  INV_X1    g556(.A(new_n750), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n755), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n749), .B1(new_n754), .B2(new_n759), .ZN(G1331gat));
  NAND2_X1  g559(.A1(new_n710), .A2(new_n517), .ZN(new_n761));
  INV_X1    g560(.A(new_n625), .ZN(new_n762));
  NOR4_X1   g561(.A1(new_n762), .A2(new_n675), .A3(new_n712), .A4(new_n649), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT106), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(KEYINPUT106), .B1(new_n761), .B2(new_n763), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n702), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g569(.A(new_n764), .B(new_n765), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n514), .B(KEYINPUT107), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n774));
  AND2_X1   g573(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(new_n773), .B2(new_n774), .ZN(G1333gat));
  OAI21_X1  g576(.A(new_n580), .B1(new_n771), .B2(new_n727), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n509), .A2(new_n580), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT108), .B1(new_n768), .B2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT108), .ZN(new_n781));
  INV_X1    g580(.A(new_n779), .ZN(new_n782));
  NOR4_X1   g581(.A1(new_n766), .A2(new_n767), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n778), .B1(new_n780), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT50), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT50), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n778), .B(new_n786), .C1(new_n780), .C2(new_n783), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(G1334gat));
  NAND2_X1  g587(.A1(new_n768), .A2(new_n479), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g589(.A1(new_n625), .A2(new_n675), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n792), .A2(new_n649), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n716), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n702), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT109), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT109), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n794), .A2(new_n797), .A3(new_n702), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n796), .A2(G85gat), .A3(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT110), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n761), .A2(new_n801), .A3(new_n712), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n791), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n576), .B1(new_n710), .B2(new_n517), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n804), .A2(new_n801), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n800), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT110), .B1(new_n711), .B2(new_n576), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n792), .B1(new_n804), .B2(new_n801), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT111), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n807), .A2(new_n808), .A3(new_n809), .A4(KEYINPUT51), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n806), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n807), .A2(new_n808), .A3(KEYINPUT51), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(KEYINPUT111), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n702), .A2(new_n545), .A3(new_n648), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n799), .B1(new_n814), .B2(new_n815), .ZN(G1336gat));
  XOR2_X1   g615(.A(new_n514), .B(KEYINPUT107), .Z(new_n817));
  NAND3_X1  g616(.A1(new_n817), .A2(new_n546), .A3(new_n648), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(KEYINPUT112), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n819), .B1(new_n806), .B2(new_n812), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n546), .B1(new_n794), .B2(new_n720), .ZN(new_n821));
  OAI21_X1  g620(.A(KEYINPUT52), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n819), .B1(new_n811), .B2(new_n813), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n794), .A2(new_n817), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(G92gat), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n822), .B1(new_n823), .B2(new_n827), .ZN(G1337gat));
  NAND2_X1  g627(.A1(new_n794), .A2(new_n731), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(G99gat), .ZN(new_n830));
  OR3_X1    g629(.A1(new_n727), .A2(G99gat), .A3(new_n649), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n830), .B1(new_n814), .B2(new_n831), .ZN(G1338gat));
  NOR3_X1   g631(.A1(new_n438), .A2(new_n649), .A3(G106gat), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT114), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n834), .B1(new_n806), .B2(new_n812), .ZN(new_n835));
  XOR2_X1   g634(.A(KEYINPUT113), .B(G106gat), .Z(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n837), .B1(new_n794), .B2(new_n479), .ZN(new_n838));
  OAI21_X1  g637(.A(KEYINPUT53), .B1(new_n835), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n834), .B1(new_n811), .B2(new_n813), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n794), .A2(new_n479), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n836), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT53), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n839), .B1(new_n840), .B2(new_n844), .ZN(G1339gat));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n634), .A2(new_n627), .A3(new_n635), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n645), .A2(KEYINPUT54), .A3(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n642), .B1(new_n636), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT55), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n848), .A2(KEYINPUT55), .A3(new_n850), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n647), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n851), .B1(new_n853), .B2(KEYINPUT115), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT115), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n852), .A2(new_n855), .A3(new_n647), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n675), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n669), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n657), .B1(new_n655), .B2(new_n658), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n656), .B1(new_n661), .B2(new_n651), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n674), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n648), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n712), .B1(new_n857), .B2(new_n863), .ZN(new_n864));
  AND4_X1   g663(.A1(new_n712), .A2(new_n862), .A3(new_n854), .A4(new_n856), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n762), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n650), .A2(new_n675), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n479), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n817), .A2(new_n727), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n868), .A2(new_n702), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(G113gat), .B1(new_n870), .B2(new_n676), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n871), .B(KEYINPUT116), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n676), .A2(G113gat), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n508), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n868), .A2(new_n702), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(KEYINPUT117), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT117), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n868), .A2(new_n878), .A3(new_n702), .A4(new_n875), .ZN(new_n879));
  AOI211_X1 g678(.A(new_n817), .B(new_n874), .C1(new_n877), .C2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n846), .B1(new_n872), .B2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT116), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n871), .B(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n877), .ZN(new_n884));
  INV_X1    g683(.A(new_n879), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n772), .B(new_n873), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n883), .A2(KEYINPUT118), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n881), .A2(new_n887), .ZN(G1340gat));
  NOR3_X1   g687(.A1(new_n870), .A2(new_n325), .A3(new_n649), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n772), .B1(new_n884), .B2(new_n885), .ZN(new_n890));
  OR2_X1    g689(.A1(new_n890), .A2(new_n649), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n889), .B1(new_n891), .B2(new_n325), .ZN(G1341gat));
  OAI21_X1  g691(.A(G127gat), .B1(new_n870), .B2(new_n762), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n625), .A2(new_n321), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n893), .B1(new_n890), .B2(new_n894), .ZN(G1342gat));
  NOR2_X1   g694(.A1(new_n720), .A2(new_n576), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n319), .B(new_n896), .C1(new_n884), .C2(new_n885), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n897), .A2(KEYINPUT56), .ZN(new_n898));
  OAI21_X1  g697(.A(G134gat), .B1(new_n870), .B2(new_n576), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(KEYINPUT56), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(G1343gat));
  NAND2_X1  g700(.A1(new_n866), .A2(new_n867), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n479), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n772), .A2(new_n702), .A3(new_n509), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n676), .A2(G141gat), .ZN(new_n906));
  AOI21_X1  g705(.A(KEYINPUT58), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n438), .B1(new_n866), .B2(new_n867), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT57), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n904), .A2(KEYINPUT119), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT119), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n772), .A2(new_n913), .A3(new_n702), .A4(new_n509), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n853), .A2(new_n851), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n675), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n712), .B1(new_n916), .B2(new_n863), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n762), .B1(new_n917), .B2(new_n865), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n438), .B1(new_n918), .B2(new_n867), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n912), .B(new_n914), .C1(new_n919), .C2(new_n909), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n911), .A2(new_n920), .A3(new_n676), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n907), .B1(new_n921), .B2(new_n337), .ZN(new_n922));
  OAI21_X1  g721(.A(KEYINPUT120), .B1(new_n911), .B2(new_n920), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n919), .A2(new_n909), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT120), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n912), .A2(new_n914), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n924), .A2(new_n925), .A3(new_n926), .A4(new_n910), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n923), .A2(new_n927), .A3(new_n675), .ZN(new_n928));
  AOI22_X1  g727(.A1(new_n928), .A2(G141gat), .B1(new_n905), .B2(new_n906), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT58), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n922), .B1(new_n929), .B2(new_n930), .ZN(G1344gat));
  NAND3_X1  g730(.A1(new_n905), .A2(new_n338), .A3(new_n648), .ZN(new_n932));
  OR2_X1    g731(.A1(new_n338), .A2(KEYINPUT59), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n923), .A2(new_n927), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n933), .B1(new_n934), .B2(new_n648), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n912), .A2(new_n648), .A3(new_n914), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n903), .A2(KEYINPUT57), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n848), .A2(new_n850), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT55), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n941), .A2(new_n647), .A3(new_n852), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n942), .B1(new_n673), .B2(new_n674), .ZN(new_n943));
  AND3_X1   g742(.A1(new_n648), .A2(new_n674), .A3(new_n861), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n576), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n712), .A2(new_n862), .A3(new_n854), .A4(new_n856), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n625), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n650), .A2(new_n675), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n909), .B(new_n479), .C1(new_n947), .C2(new_n948), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n937), .A2(new_n938), .A3(KEYINPUT121), .A4(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT121), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n949), .B1(new_n908), .B2(new_n909), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n952), .B2(new_n936), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n950), .A2(new_n953), .A3(G148gat), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n954), .A2(KEYINPUT59), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n932), .B1(new_n935), .B2(new_n955), .ZN(G1345gat));
  AOI21_X1  g755(.A(G155gat), .B1(new_n905), .B2(new_n625), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n625), .A2(G155gat), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n958), .B(KEYINPUT122), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n957), .B1(new_n934), .B2(new_n959), .ZN(G1346gat));
  NAND2_X1  g759(.A1(new_n934), .A2(new_n712), .ZN(new_n961));
  INV_X1    g760(.A(new_n350), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n475), .A2(new_n962), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n908), .A2(new_n509), .A3(new_n896), .A4(new_n964), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n963), .A2(new_n965), .ZN(G1347gat));
  OR2_X1    g765(.A1(new_n772), .A2(new_n511), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT123), .ZN(new_n968));
  OR2_X1    g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n702), .B1(new_n866), .B2(new_n867), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n967), .A2(new_n968), .ZN(new_n971));
  AND3_X1   g770(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g771(.A(G169gat), .B1(new_n972), .B2(new_n675), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n702), .A2(new_n514), .ZN(new_n974));
  AND3_X1   g773(.A1(new_n868), .A2(new_n515), .A3(new_n974), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n676), .A2(new_n223), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(G1348gat));
  AOI21_X1  g776(.A(G176gat), .B1(new_n972), .B2(new_n648), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n649), .A2(new_n224), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n978), .B1(new_n975), .B2(new_n979), .ZN(G1349gat));
  NAND3_X1  g779(.A1(new_n972), .A2(new_n212), .A3(new_n625), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n975), .A2(new_n625), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(G183gat), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT124), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n984), .A2(KEYINPUT60), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n981), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  OR2_X1    g785(.A1(new_n984), .A2(KEYINPUT60), .ZN(new_n987));
  XNOR2_X1  g786(.A(new_n986), .B(new_n987), .ZN(G1350gat));
  AOI21_X1  g787(.A(new_n208), .B1(new_n975), .B2(new_n712), .ZN(new_n989));
  XOR2_X1   g788(.A(new_n989), .B(KEYINPUT61), .Z(new_n990));
  NAND3_X1  g789(.A1(new_n972), .A2(new_n208), .A3(new_n712), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(G1351gat));
  NAND4_X1  g791(.A1(new_n970), .A2(new_n479), .A3(new_n509), .A4(new_n817), .ZN(new_n993));
  NOR2_X1   g792(.A1(new_n993), .A2(new_n676), .ZN(new_n994));
  AND2_X1   g793(.A1(new_n509), .A2(new_n974), .ZN(new_n995));
  OAI211_X1 g794(.A(new_n949), .B(new_n995), .C1(new_n908), .C2(new_n909), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n675), .A2(G197gat), .ZN(new_n997));
  OAI22_X1  g796(.A1(new_n994), .A2(G197gat), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g797(.A(new_n998), .ZN(G1352gat));
  NOR3_X1   g798(.A1(new_n993), .A2(G204gat), .A3(new_n649), .ZN(new_n1000));
  XNOR2_X1  g799(.A(new_n1000), .B(KEYINPUT62), .ZN(new_n1001));
  OAI21_X1  g800(.A(G204gat), .B1(new_n996), .B2(new_n649), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1001), .A2(new_n1002), .ZN(G1353gat));
  INV_X1    g802(.A(G211gat), .ZN(new_n1004));
  INV_X1    g803(.A(KEYINPUT63), .ZN(new_n1005));
  AOI21_X1  g804(.A(new_n1004), .B1(KEYINPUT127), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g805(.A(KEYINPUT126), .ZN(new_n1007));
  INV_X1    g806(.A(new_n996), .ZN(new_n1008));
  AOI21_X1  g807(.A(new_n1007), .B1(new_n1008), .B2(new_n625), .ZN(new_n1009));
  NOR3_X1   g808(.A1(new_n996), .A2(KEYINPUT126), .A3(new_n762), .ZN(new_n1010));
  OAI21_X1  g809(.A(new_n1006), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g810(.A1(new_n1005), .A2(KEYINPUT127), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI221_X1 g812(.A(new_n1006), .B1(KEYINPUT127), .B2(new_n1005), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1014));
  NOR3_X1   g813(.A1(new_n993), .A2(G211gat), .A3(new_n762), .ZN(new_n1015));
  XNOR2_X1  g814(.A(new_n1015), .B(KEYINPUT125), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n1013), .A2(new_n1014), .A3(new_n1016), .ZN(G1354gat));
  OAI21_X1  g816(.A(G218gat), .B1(new_n996), .B2(new_n576), .ZN(new_n1018));
  OR2_X1    g817(.A1(new_n576), .A2(G218gat), .ZN(new_n1019));
  OAI21_X1  g818(.A(new_n1018), .B1(new_n993), .B2(new_n1019), .ZN(G1355gat));
endmodule


