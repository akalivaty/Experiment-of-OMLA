//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 0 0 1 0 1 0 1 0 0 1 1 1 0 0 1 0 0 1 0 1 0 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G210), .B1(G237), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  OAI21_X1  g005(.A(KEYINPUT3), .B1(new_n191), .B2(G107), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(new_n194), .A3(G104), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n191), .A2(G107), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n192), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  AND2_X1   g011(.A1(new_n197), .A2(G101), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT4), .ZN(new_n199));
  XOR2_X1   g013(.A(KEYINPUT2), .B(G113), .Z(new_n200));
  INV_X1    g014(.A(G116), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT65), .B1(new_n201), .B2(G119), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT65), .ZN(new_n203));
  INV_X1    g017(.A(G119), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(new_n204), .A3(G116), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n201), .A2(G119), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n200), .A2(new_n202), .A3(new_n205), .A4(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n202), .A2(new_n205), .A3(new_n206), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT2), .B(G113), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AOI22_X1  g024(.A1(new_n198), .A2(new_n199), .B1(new_n207), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(G101), .B1(new_n191), .B2(G107), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n192), .A2(new_n212), .A3(new_n195), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT72), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT72), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n192), .A2(new_n212), .A3(new_n195), .A4(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n199), .B1(new_n197), .B2(G101), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n191), .A2(G107), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n194), .A2(G104), .ZN(new_n221));
  OAI21_X1  g035(.A(G101), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n223), .B1(new_n214), .B2(new_n216), .ZN(new_n224));
  INV_X1    g038(.A(new_n208), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n202), .A2(new_n205), .A3(KEYINPUT5), .A4(new_n206), .ZN(new_n226));
  NOR3_X1   g040(.A1(new_n201), .A2(KEYINPUT5), .A3(G119), .ZN(new_n227));
  INV_X1    g041(.A(G113), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n225), .A2(new_n200), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n211), .A2(new_n219), .B1(new_n224), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(G110), .B(G122), .ZN(new_n232));
  NOR3_X1   g046(.A1(new_n231), .A2(KEYINPUT6), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G143), .ZN(new_n234));
  OAI21_X1  g048(.A(KEYINPUT1), .B1(new_n234), .B2(G146), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n234), .A2(G146), .ZN(new_n236));
  INV_X1    g050(.A(G146), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(G143), .ZN(new_n238));
  OAI211_X1 g052(.A(G128), .B(new_n235), .C1(new_n236), .C2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G125), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n237), .A2(G143), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n234), .A2(G146), .ZN(new_n242));
  INV_X1    g056(.A(G128), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n241), .B(new_n242), .C1(KEYINPUT1), .C2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n239), .A2(new_n240), .A3(new_n244), .ZN(new_n245));
  AND2_X1   g059(.A1(KEYINPUT0), .A2(G128), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n241), .A2(new_n242), .A3(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(G143), .B(G146), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT0), .B(G128), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n247), .B(G125), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n245), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G953), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G224), .ZN(new_n253));
  XOR2_X1   g067(.A(new_n253), .B(KEYINPUT76), .Z(new_n254));
  XNOR2_X1  g068(.A(new_n251), .B(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n224), .A2(new_n230), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n217), .A2(new_n218), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n207), .A2(new_n210), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n197), .A2(new_n199), .A3(G101), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n256), .B(new_n232), .C1(new_n257), .C2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT75), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT75), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n231), .A2(new_n263), .A3(new_n232), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n231), .A2(new_n232), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI211_X1 g082(.A(new_n233), .B(new_n255), .C1(new_n265), .C2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT78), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT7), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n271), .A2(KEYINPUT77), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n272), .B1(new_n245), .B2(new_n250), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n253), .A2(KEYINPUT7), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n273), .B(new_n275), .ZN(new_n276));
  XOR2_X1   g090(.A(new_n232), .B(KEYINPUT8), .Z(new_n277));
  NAND2_X1  g091(.A1(new_n217), .A2(new_n222), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n226), .A2(new_n229), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n207), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n277), .B1(new_n281), .B2(new_n256), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n270), .B1(new_n276), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n277), .ZN(new_n284));
  INV_X1    g098(.A(new_n256), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n224), .A2(new_n230), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n273), .B(new_n274), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n287), .A2(new_n288), .A3(KEYINPUT78), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n265), .A2(new_n283), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G902), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n190), .B1(new_n269), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n265), .A2(new_n268), .ZN(new_n294));
  INV_X1    g108(.A(new_n233), .ZN(new_n295));
  INV_X1    g109(.A(new_n255), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n297), .A2(new_n291), .A3(new_n290), .A4(new_n189), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n188), .B1(new_n293), .B2(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(KEYINPUT9), .B(G234), .ZN(new_n300));
  OAI21_X1  g114(.A(G221), .B1(new_n300), .B2(G902), .ZN(new_n301));
  INV_X1    g115(.A(G469), .ZN(new_n302));
  XNOR2_X1  g116(.A(G110), .B(G140), .ZN(new_n303));
  INV_X1    g117(.A(G227), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n304), .A2(G953), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n303), .B(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT11), .ZN(new_n308));
  INV_X1    g122(.A(G134), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n308), .B1(new_n309), .B2(G137), .ZN(new_n310));
  INV_X1    g124(.A(G137), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(KEYINPUT11), .A3(G134), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n309), .A2(G137), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n310), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G131), .ZN(new_n315));
  INV_X1    g129(.A(G131), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n310), .A2(new_n312), .A3(new_n316), .A4(new_n313), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n219), .A2(new_n320), .A3(new_n259), .ZN(new_n321));
  AND3_X1   g135(.A1(new_n239), .A2(new_n244), .A3(new_n222), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n217), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT10), .ZN(new_n324));
  AOI21_X1  g138(.A(KEYINPUT73), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT73), .ZN(new_n326));
  AOI211_X1 g140(.A(new_n326), .B(KEYINPUT10), .C1(new_n322), .C2(new_n217), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n321), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n322), .A2(new_n217), .A3(KEYINPUT10), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT74), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n322), .A2(new_n217), .A3(KEYINPUT74), .A4(KEYINPUT10), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n318), .B1(new_n328), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n239), .A2(new_n244), .A3(new_n222), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n336), .B1(new_n216), .B2(new_n214), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n326), .B1(new_n337), .B2(KEYINPUT10), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n323), .A2(KEYINPUT73), .A3(new_n324), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n318), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n340), .A2(new_n341), .A3(new_n333), .A4(new_n321), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n307), .B1(new_n335), .B2(new_n342), .ZN(new_n343));
  AOI22_X1  g157(.A1(new_n217), .A2(new_n222), .B1(new_n244), .B2(new_n239), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n318), .B1(new_n344), .B2(new_n337), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT12), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI211_X1 g161(.A(KEYINPUT12), .B(new_n318), .C1(new_n344), .C2(new_n337), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n342), .A2(new_n349), .A3(new_n307), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n302), .B(new_n291), .C1(new_n343), .C2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(G469), .A2(G902), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n342), .A2(new_n349), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n306), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n335), .A2(new_n342), .A3(new_n307), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n355), .A3(G469), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n351), .A2(new_n352), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n299), .A2(new_n301), .A3(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(G113), .B(G122), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n359), .B(new_n191), .ZN(new_n360));
  NOR3_X1   g174(.A1(new_n240), .A2(KEYINPUT16), .A3(G140), .ZN(new_n361));
  XNOR2_X1  g175(.A(G125), .B(G140), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n361), .B1(new_n362), .B2(KEYINPUT16), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n363), .A2(G146), .ZN(new_n364));
  AOI211_X1 g178(.A(new_n237), .B(new_n361), .C1(KEYINPUT16), .C2(new_n362), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AND2_X1   g180(.A1(KEYINPUT66), .A2(G237), .ZN(new_n367));
  NOR2_X1   g181(.A1(KEYINPUT66), .A2(G237), .ZN(new_n368));
  OAI211_X1 g182(.A(G214), .B(new_n252), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n234), .ZN(new_n370));
  XNOR2_X1  g184(.A(KEYINPUT66), .B(G237), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n371), .A2(G143), .A3(G214), .A4(new_n252), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(KEYINPUT17), .A3(G131), .ZN(new_n374));
  OR2_X1    g188(.A1(KEYINPUT66), .A2(G237), .ZN(new_n375));
  NAND2_X1  g189(.A1(KEYINPUT66), .A2(G237), .ZN(new_n376));
  AOI21_X1  g190(.A(G953), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(G143), .B1(new_n377), .B2(G214), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n369), .A2(new_n234), .ZN(new_n379));
  OAI21_X1  g193(.A(G131), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n370), .A2(new_n372), .A3(new_n316), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n366), .B(new_n374), .C1(new_n382), .C2(KEYINPUT17), .ZN(new_n383));
  NAND2_X1  g197(.A1(KEYINPUT18), .A2(G131), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n370), .A2(new_n372), .A3(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n362), .B(new_n237), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n384), .ZN(new_n388));
  AOI21_X1  g202(.A(KEYINPUT79), .B1(new_n373), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT79), .ZN(new_n390));
  AOI211_X1 g204(.A(new_n390), .B(new_n384), .C1(new_n370), .C2(new_n372), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n387), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n360), .B1(new_n383), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n383), .A2(new_n360), .A3(new_n392), .ZN(new_n395));
  AOI21_X1  g209(.A(G902), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G475), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT81), .ZN(new_n399));
  NOR2_X1   g213(.A1(KEYINPUT80), .A2(KEYINPUT19), .ZN(new_n400));
  AND2_X1   g214(.A1(KEYINPUT80), .A2(KEYINPUT19), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n362), .B(new_n399), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G140), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G125), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n240), .A2(G140), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n404), .B(new_n405), .C1(new_n401), .C2(new_n400), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT81), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT19), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n362), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n402), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n365), .B1(new_n410), .B2(new_n237), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n382), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT82), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n392), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n360), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n413), .B1(new_n392), .B2(new_n412), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n395), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(G475), .A2(G902), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT20), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT20), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n418), .A2(new_n422), .A3(new_n419), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n398), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(G122), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT83), .B1(new_n425), .B2(G116), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT83), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(new_n201), .A3(G122), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  OR2_X1    g243(.A1(new_n201), .A2(G122), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n429), .A2(new_n194), .A3(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT85), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n234), .A2(G128), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n243), .A2(G143), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(new_n434), .A3(new_n309), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n433), .A2(new_n434), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(G134), .ZN(new_n437));
  AOI22_X1  g251(.A1(new_n431), .A2(new_n432), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n429), .A2(KEYINPUT14), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT14), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n426), .A2(new_n428), .A3(new_n440), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n439), .A2(new_n430), .A3(new_n441), .ZN(new_n442));
  OAI221_X1 g256(.A(new_n438), .B1(new_n432), .B2(new_n431), .C1(new_n442), .C2(new_n194), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n234), .A2(KEYINPUT13), .A3(G128), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n434), .ZN(new_n445));
  AOI21_X1  g259(.A(KEYINPUT13), .B1(new_n234), .B2(G128), .ZN(new_n446));
  OAI21_X1  g260(.A(G134), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n447), .B(KEYINPUT84), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n429), .A2(new_n430), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G107), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n431), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n448), .A2(new_n435), .A3(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(G217), .ZN(new_n453));
  NOR3_X1   g267(.A1(new_n300), .A2(new_n453), .A3(G953), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n443), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n454), .B1(new_n443), .B2(new_n452), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n291), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G478), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n459), .A2(KEYINPUT15), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n458), .B(new_n460), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n252), .A2(G952), .ZN(new_n462));
  INV_X1    g276(.A(G234), .ZN(new_n463));
  INV_X1    g277(.A(G237), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  AOI211_X1 g280(.A(new_n291), .B(new_n252), .C1(G234), .C2(G237), .ZN(new_n467));
  XNOR2_X1  g281(.A(KEYINPUT21), .B(G898), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n461), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n424), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(KEYINPUT86), .B1(new_n358), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n471), .ZN(new_n473));
  INV_X1    g287(.A(new_n301), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n342), .A2(new_n307), .ZN(new_n475));
  AOI22_X1  g289(.A1(new_n475), .A2(new_n335), .B1(new_n353), .B2(new_n306), .ZN(new_n476));
  OAI21_X1  g290(.A(G469), .B1(new_n476), .B2(G902), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n474), .B1(new_n477), .B2(new_n351), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT86), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n473), .A2(new_n478), .A3(new_n479), .A4(new_n299), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n472), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n453), .B1(G234), .B2(new_n291), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n243), .A2(G119), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n204), .A2(G128), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  XOR2_X1   g299(.A(KEYINPUT24), .B(G110), .Z(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(new_n486), .A3(KEYINPUT69), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT69), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n483), .A2(new_n484), .ZN(new_n489));
  XNOR2_X1  g303(.A(KEYINPUT24), .B(G110), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT23), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n493), .B1(new_n204), .B2(G128), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n243), .A2(KEYINPUT23), .A3(G119), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n494), .A2(new_n495), .A3(new_n484), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(G110), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n492), .B(new_n497), .C1(new_n364), .C2(new_n365), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n363), .A2(G146), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n362), .A2(new_n237), .ZN(new_n500));
  INV_X1    g314(.A(G110), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n494), .A2(new_n495), .A3(new_n501), .A4(new_n484), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT70), .ZN(new_n503));
  OAI22_X1  g317(.A1(new_n502), .A2(new_n503), .B1(new_n485), .B2(new_n486), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n502), .A2(new_n503), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n499), .B(new_n500), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n498), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(KEYINPUT22), .B(G137), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n252), .A2(G221), .A3(G234), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n498), .A2(new_n506), .A3(new_n510), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(new_n291), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT71), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n515), .A2(KEYINPUT25), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n514), .A2(new_n516), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n482), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n512), .A2(new_n513), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n482), .A2(G902), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n519), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n239), .A2(new_n317), .A3(new_n244), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT64), .B1(new_n309), .B2(G137), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT64), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(new_n311), .A3(G134), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n527), .A2(new_n529), .A3(new_n313), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n530), .A2(G131), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n319), .B1(new_n317), .B2(new_n315), .ZN(new_n533));
  NOR3_X1   g347(.A1(new_n532), .A2(new_n533), .A3(new_n258), .ZN(new_n534));
  AND2_X1   g348(.A1(new_n207), .A2(new_n210), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n318), .A2(new_n320), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n530), .A2(G131), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n537), .A2(new_n317), .A3(new_n244), .A4(new_n239), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n535), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT28), .B1(new_n534), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g354(.A(G210), .B(new_n252), .C1(new_n367), .C2(new_n368), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT27), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT27), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n371), .A2(new_n543), .A3(G210), .A4(new_n252), .ZN(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT26), .B(G101), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n542), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n545), .B1(new_n542), .B2(new_n544), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n536), .A2(new_n535), .A3(new_n538), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT28), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n540), .A2(new_n548), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n548), .ZN(new_n553));
  OAI21_X1  g367(.A(KEYINPUT30), .B1(new_n532), .B2(new_n533), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT30), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n536), .A2(new_n555), .A3(new_n538), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n535), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n553), .B1(new_n557), .B2(new_n534), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT29), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n552), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n291), .B1(new_n552), .B2(new_n559), .ZN(new_n561));
  OAI21_X1  g375(.A(G472), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT68), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI211_X1 g378(.A(KEYINPUT68), .B(G472), .C1(new_n560), .C2(new_n561), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(G472), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT31), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT67), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n549), .A2(new_n569), .A3(new_n548), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(new_n557), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n549), .A2(new_n548), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(KEYINPUT67), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n568), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n532), .A2(new_n533), .A3(KEYINPUT30), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n555), .B1(new_n536), .B2(new_n538), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n258), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n578), .A2(new_n574), .A3(new_n568), .A4(new_n570), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n258), .B1(new_n532), .B2(new_n533), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n550), .B1(new_n580), .B2(new_n549), .ZN(new_n581));
  INV_X1    g395(.A(new_n551), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n553), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n567), .B(new_n291), .C1(new_n575), .C2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT32), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n578), .A2(new_n574), .A3(new_n570), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT31), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n588), .A2(new_n583), .A3(new_n579), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT32), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n589), .A2(new_n590), .A3(new_n567), .A4(new_n291), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n586), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n525), .B1(new_n566), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n481), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g409(.A(new_n595), .B(G101), .Z(G3));
  NAND2_X1  g410(.A1(new_n357), .A2(new_n301), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n589), .A2(new_n291), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(G472), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n514), .B(new_n516), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n523), .B1(new_n600), .B2(new_n482), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n599), .A2(new_n585), .A3(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT87), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n597), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n585), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n567), .B1(new_n589), .B2(new_n291), .ZN(new_n606));
  NOR3_X1   g420(.A1(new_n605), .A2(new_n606), .A3(new_n525), .ZN(new_n607));
  AOI21_X1  g421(.A(KEYINPUT87), .B1(new_n478), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n293), .A2(new_n298), .ZN(new_n610));
  INV_X1    g424(.A(new_n469), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n610), .A2(new_n187), .A3(new_n611), .ZN(new_n612));
  OR2_X1    g426(.A1(new_n396), .A2(new_n397), .ZN(new_n613));
  INV_X1    g427(.A(new_n423), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n422), .B1(new_n418), .B2(new_n419), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT33), .ZN(new_n617));
  OAI22_X1  g431(.A1(new_n456), .A2(new_n457), .B1(KEYINPUT88), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n457), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT88), .B(KEYINPUT33), .Z(new_n620));
  NAND3_X1  g434(.A1(new_n619), .A2(new_n455), .A3(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n459), .A2(G902), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n618), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n458), .A2(new_n459), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n616), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n612), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n609), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(KEYINPUT89), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT34), .B(G104), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G6));
  INV_X1    g446(.A(new_n612), .ZN(new_n633));
  INV_X1    g447(.A(new_n460), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n458), .B(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(new_n398), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT90), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n421), .A2(new_n637), .A3(new_n423), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n615), .A2(KEYINPUT90), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n636), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n609), .A2(new_n633), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT35), .B(G107), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G9));
  NAND2_X1  g457(.A1(new_n507), .A2(KEYINPUT91), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT91), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n498), .A2(new_n506), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n511), .A2(KEYINPUT36), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n644), .A2(new_n648), .A3(new_n646), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n522), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n652), .B1(new_n600), .B2(new_n482), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n654), .A2(new_n599), .A3(new_n585), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n481), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT37), .B(G110), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G12));
  INV_X1    g472(.A(new_n358), .ZN(new_n659));
  INV_X1    g473(.A(G900), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n467), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n465), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n636), .A2(new_n638), .A3(new_n639), .A4(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n653), .B1(new_n566), .B2(new_n592), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n659), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G128), .ZN(G30));
  XNOR2_X1  g481(.A(KEYINPUT93), .B(KEYINPUT39), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n662), .B(new_n668), .ZN(new_n669));
  AND2_X1   g483(.A1(new_n478), .A2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT40), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n610), .B(KEYINPUT38), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n616), .A2(new_n461), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n674), .A2(new_n188), .A3(new_n654), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n672), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n548), .B1(new_n580), .B2(new_n549), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n677), .B1(new_n572), .B2(new_n574), .ZN(new_n678));
  OAI21_X1  g492(.A(G472), .B1(new_n678), .B2(G902), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n592), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT92), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n670), .A2(new_n671), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n676), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT94), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G143), .ZN(G45));
  NAND3_X1  g499(.A1(new_n616), .A2(new_n626), .A3(new_n662), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n659), .A2(new_n687), .A3(new_n665), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G146), .ZN(G48));
  NAND2_X1  g503(.A1(new_n566), .A2(new_n592), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n291), .B1(new_n343), .B2(new_n350), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(G469), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n692), .A2(new_n301), .A3(new_n351), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n690), .A2(new_n693), .A3(new_n601), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n421), .A2(new_n423), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n625), .B1(new_n695), .B2(new_n613), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n696), .A2(new_n299), .A3(new_n611), .ZN(new_n697));
  OAI21_X1  g511(.A(KEYINPUT95), .B1(new_n694), .B2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT95), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n628), .A2(new_n699), .A3(new_n593), .A4(new_n693), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT41), .B(G113), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G15));
  NAND4_X1  g517(.A1(new_n593), .A2(new_n633), .A3(new_n640), .A4(new_n693), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G116), .ZN(G18));
  NAND2_X1  g519(.A1(new_n610), .A2(new_n187), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n692), .A2(new_n301), .A3(new_n351), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(new_n665), .A3(new_n473), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT96), .B(G119), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G21));
  INV_X1    g525(.A(new_n674), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n602), .A2(new_n469), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n708), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G122), .ZN(G24));
  NOR2_X1   g529(.A1(new_n686), .A2(new_n655), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n708), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G125), .ZN(G27));
  NAND3_X1  g532(.A1(new_n293), .A2(new_n187), .A3(new_n298), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT97), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n293), .A2(new_n298), .A3(KEYINPUT97), .A4(new_n187), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n593), .A2(new_n478), .A3(new_n721), .A4(new_n722), .ZN(new_n723));
  AND2_X1   g537(.A1(KEYINPUT98), .A2(KEYINPUT42), .ZN(new_n724));
  NOR2_X1   g538(.A1(KEYINPUT98), .A2(KEYINPUT42), .ZN(new_n725));
  OAI22_X1  g539(.A1(new_n723), .A2(new_n686), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n721), .A2(new_n478), .A3(new_n722), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(new_n593), .A3(new_n687), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n726), .B1(new_n728), .B2(new_n725), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G131), .ZN(G33));
  INV_X1    g544(.A(KEYINPUT99), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n663), .A2(new_n731), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n638), .A2(new_n639), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n733), .A2(KEYINPUT99), .A3(new_n636), .A4(new_n662), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n727), .A2(new_n593), .A3(new_n732), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G134), .ZN(G36));
  NAND2_X1  g550(.A1(new_n354), .A2(new_n355), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT45), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n302), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n739), .B1(new_n738), .B2(new_n737), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n740), .A2(new_n352), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT46), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n351), .ZN(new_n743));
  OR2_X1    g557(.A1(new_n743), .A2(KEYINPUT100), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n741), .A2(KEYINPUT46), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n745), .B1(new_n743), .B2(KEYINPUT100), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n474), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n747), .A2(new_n669), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n424), .B(KEYINPUT102), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(KEYINPUT43), .A3(new_n626), .ZN(new_n750));
  XNOR2_X1  g564(.A(KEYINPUT101), .B(KEYINPUT43), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n751), .B1(new_n616), .B2(new_n625), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n653), .B1(new_n599), .B2(new_n585), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT44), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n721), .A2(new_n722), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n753), .A2(KEYINPUT44), .A3(new_n754), .ZN(new_n759));
  AND3_X1   g573(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n748), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G137), .ZN(G39));
  OR2_X1    g576(.A1(new_n747), .A2(KEYINPUT47), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n747), .A2(KEYINPUT47), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n758), .A2(new_n687), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n766), .A2(new_n690), .A3(new_n601), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G140), .ZN(G42));
  NAND3_X1  g583(.A1(new_n626), .A2(new_n187), .A3(new_n301), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n673), .A2(new_n525), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n692), .A2(new_n351), .ZN(new_n772));
  XOR2_X1   g586(.A(new_n772), .B(KEYINPUT49), .Z(new_n773));
  NAND4_X1  g587(.A1(new_n771), .A2(new_n681), .A3(new_n749), .A4(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n662), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n674), .A2(new_n654), .A3(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n776), .A2(new_n659), .A3(new_n680), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n777), .A2(new_n666), .A3(new_n688), .A4(new_n717), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(KEYINPUT106), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n778), .B(new_n780), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n781), .B1(new_n782), .B2(new_n779), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n461), .A2(new_n398), .A3(new_n775), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n727), .A2(new_n733), .A3(new_n665), .A4(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT105), .B1(new_n727), .B2(new_n716), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n721), .A2(new_n478), .A3(new_n722), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n605), .A2(new_n606), .A3(new_n653), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(new_n696), .A3(new_n662), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT105), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n788), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n735), .B(new_n786), .C1(new_n787), .C2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT104), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n613), .B(new_n461), .C1(new_n614), .C2(new_n615), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n794), .B1(new_n612), .B2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n795), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n797), .A2(new_n299), .A3(KEYINPUT104), .A4(new_n611), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n796), .A2(new_n697), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n609), .A2(new_n799), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n472), .B(new_n480), .C1(new_n593), .C2(new_n789), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n793), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT103), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n698), .A2(new_n700), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n704), .A2(new_n709), .A3(new_n714), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n806), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n808), .A2(KEYINPUT103), .A3(new_n701), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n803), .A2(new_n807), .A3(new_n729), .A4(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n810), .A2(KEYINPUT53), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n784), .A2(new_n811), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n805), .A2(new_n804), .A3(new_n806), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT103), .B1(new_n808), .B2(new_n701), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n815), .A2(new_n782), .A3(new_n729), .A4(new_n803), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT53), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n812), .A2(new_n817), .A3(KEYINPUT54), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(KEYINPUT107), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT53), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n778), .B(KEYINPUT52), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n820), .B1(new_n810), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(KEYINPUT108), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT108), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n824), .B(new_n820), .C1(new_n810), .C2(new_n821), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(KEYINPUT110), .B(KEYINPUT54), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n793), .A2(new_n802), .A3(new_n820), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n806), .B1(new_n700), .B2(new_n698), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n829), .A2(KEYINPUT109), .A3(new_n729), .ZN(new_n830));
  AOI21_X1  g644(.A(KEYINPUT109), .B1(new_n829), .B2(new_n729), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n828), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(new_n783), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n826), .A2(new_n827), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT111), .B1(new_n819), .B2(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n812), .A2(new_n817), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(KEYINPUT107), .A3(KEYINPUT54), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT107), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n818), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n838), .A2(new_n835), .A3(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT111), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n836), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n465), .B1(new_n750), .B2(new_n752), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(KEYINPUT112), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n758), .A2(new_n693), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(new_n789), .A3(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n847), .A2(new_n601), .A3(new_n466), .A4(new_n681), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n424), .A2(new_n625), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n763), .B(new_n764), .C1(new_n301), .C2(new_n772), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n846), .A2(new_n607), .A3(new_n758), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n851), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n673), .A2(new_n187), .A3(new_n707), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n846), .A2(new_n607), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT113), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT114), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT50), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n862), .B1(new_n857), .B2(KEYINPUT114), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n859), .A2(new_n860), .A3(new_n862), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n855), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT51), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n866), .A2(new_n867), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n846), .A2(new_n593), .A3(new_n847), .ZN(new_n870));
  XOR2_X1   g684(.A(new_n870), .B(KEYINPUT48), .Z(new_n871));
  NAND3_X1  g685(.A1(new_n846), .A2(new_n607), .A3(new_n708), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n872), .B(new_n462), .C1(new_n627), .C2(new_n849), .ZN(new_n873));
  OR2_X1    g687(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n868), .A2(new_n869), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT115), .B1(new_n844), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n819), .A2(KEYINPUT111), .A3(new_n835), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n841), .A2(new_n842), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n875), .A2(new_n877), .A3(new_n878), .A4(KEYINPUT115), .ZN(new_n879));
  NOR2_X1   g693(.A1(G952), .A2(G953), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT116), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n774), .B1(new_n876), .B2(new_n882), .ZN(G75));
  NOR2_X1   g697(.A1(new_n252), .A2(G952), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n291), .B1(new_n826), .B2(new_n834), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT56), .B1(new_n886), .B2(G210), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n233), .B1(new_n265), .B2(new_n268), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n888), .A2(new_n296), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n889), .A2(new_n269), .ZN(new_n890));
  XNOR2_X1  g704(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n890), .B(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n885), .B1(new_n887), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n893), .B1(new_n887), .B2(new_n892), .ZN(G51));
  INV_X1    g708(.A(new_n886), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n895), .A2(new_n740), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n343), .A2(new_n350), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n352), .B(KEYINPUT57), .Z(new_n898));
  INV_X1    g712(.A(new_n827), .ZN(new_n899));
  AOI211_X1 g713(.A(new_n899), .B(new_n833), .C1(new_n825), .C2(new_n823), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n827), .B1(new_n826), .B2(new_n834), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n897), .B1(new_n902), .B2(KEYINPUT118), .ZN(new_n903));
  INV_X1    g717(.A(new_n898), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n824), .B1(new_n816), .B2(new_n820), .ZN(new_n905));
  INV_X1    g719(.A(new_n825), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n834), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n899), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n904), .B1(new_n908), .B2(new_n835), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT118), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n896), .B1(new_n903), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(KEYINPUT119), .B1(new_n912), .B2(new_n884), .ZN(new_n913));
  INV_X1    g727(.A(new_n896), .ZN(new_n914));
  INV_X1    g728(.A(new_n897), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n915), .B1(new_n909), .B2(new_n910), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n902), .A2(KEYINPUT118), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT119), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n918), .A2(new_n919), .A3(new_n885), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n913), .A2(new_n920), .ZN(G54));
  NAND3_X1  g735(.A1(new_n886), .A2(KEYINPUT58), .A3(G475), .ZN(new_n922));
  INV_X1    g736(.A(new_n418), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n884), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n924), .B1(new_n923), .B2(new_n922), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT120), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(G60));
  NAND2_X1  g741(.A1(new_n618), .A2(new_n621), .ZN(new_n928));
  NAND2_X1  g742(.A1(G478), .A2(G902), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT59), .Z(new_n930));
  AOI211_X1 g744(.A(new_n928), .B(new_n930), .C1(new_n908), .C2(new_n835), .ZN(new_n931));
  INV_X1    g745(.A(new_n930), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n932), .B1(new_n836), .B2(new_n843), .ZN(new_n933));
  AOI211_X1 g747(.A(new_n884), .B(new_n931), .C1(new_n933), .C2(new_n928), .ZN(G63));
  NAND2_X1  g748(.A1(G217), .A2(G902), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT60), .Z(new_n936));
  NAND2_X1  g750(.A1(new_n907), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n884), .B1(new_n937), .B2(new_n520), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n650), .A2(new_n651), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n938), .B1(new_n939), .B2(new_n937), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT61), .Z(G66));
  INV_X1    g755(.A(new_n468), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n252), .B1(new_n942), .B2(G224), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n815), .A2(new_n800), .A3(new_n801), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n943), .B1(new_n944), .B2(new_n252), .ZN(new_n945));
  INV_X1    g759(.A(G898), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n888), .B1(new_n946), .B2(G953), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n945), .B(new_n947), .ZN(G69));
  INV_X1    g762(.A(KEYINPUT122), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n627), .A2(new_n795), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n758), .A2(new_n670), .A3(new_n593), .A4(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n761), .A2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT121), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n761), .A2(KEYINPUT121), .A3(new_n951), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n666), .A2(new_n717), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n957), .A2(new_n688), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n684), .A2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT62), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n684), .A2(KEYINPUT62), .A3(new_n958), .ZN(new_n962));
  AOI22_X1  g776(.A1(new_n961), .A2(new_n962), .B1(new_n765), .B2(new_n767), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n956), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n576), .A2(new_n577), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(new_n410), .Z(new_n966));
  NOR2_X1   g780(.A1(new_n966), .A2(G953), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n660), .A2(G953), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n594), .A2(new_n706), .A3(new_n674), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n748), .B1(new_n760), .B2(new_n971), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n958), .A2(new_n729), .A3(new_n735), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n768), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n970), .B1(new_n974), .B2(new_n252), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n949), .B1(new_n968), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n967), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n978), .B1(new_n956), .B2(new_n963), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n979), .A2(KEYINPUT122), .A3(new_n975), .ZN(new_n980));
  OAI21_X1  g794(.A(KEYINPUT123), .B1(new_n977), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(G953), .B1(new_n304), .B2(new_n660), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n968), .A2(new_n949), .A3(new_n976), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT123), .ZN(new_n984));
  OAI21_X1  g798(.A(KEYINPUT122), .B1(new_n979), .B2(new_n975), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n983), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n981), .A2(new_n982), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n982), .B1(new_n981), .B2(new_n986), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n987), .A2(new_n988), .ZN(G72));
  XOR2_X1   g803(.A(KEYINPUT124), .B(KEYINPUT63), .Z(new_n990));
  NOR2_X1   g804(.A1(new_n567), .A2(new_n291), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n990), .B(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n587), .A2(new_n558), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n837), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT126), .Z(new_n995));
  OAI21_X1  g809(.A(new_n992), .B1(new_n974), .B2(new_n944), .ZN(new_n996));
  NOR3_X1   g810(.A1(new_n557), .A2(new_n534), .A3(new_n548), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n884), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n992), .B1(new_n964), .B2(new_n944), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n1000), .B(KEYINPUT125), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n553), .B1(new_n578), .B2(new_n549), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n999), .B1(new_n1001), .B2(new_n1002), .ZN(G57));
endmodule


