

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771;

  AND2_X1 U371 ( .A1(n364), .A2(n398), .ZN(n354) );
  NAND2_X1 U372 ( .A1(n373), .A2(n428), .ZN(n372) );
  NAND2_X1 U373 ( .A1(n381), .A2(n436), .ZN(n595) );
  NOR2_X1 U374 ( .A1(n617), .A2(n681), .ZN(n628) );
  NOR2_X1 U375 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U376 ( .A1(n583), .A2(n582), .ZN(n584) );
  BUF_X1 U377 ( .A(n703), .Z(n374) );
  AND2_X1 U378 ( .A1(n703), .A2(n375), .ZN(n581) );
  XNOR2_X1 U379 ( .A(n389), .B(n351), .ZN(n703) );
  XNOR2_X1 U380 ( .A(n760), .B(n503), .ZN(n521) );
  XNOR2_X1 U381 ( .A(n501), .B(n500), .ZN(n760) );
  BUF_X2 U382 ( .A(G125), .Z(n348) );
  XNOR2_X2 U383 ( .A(n659), .B(n661), .ZN(n662) );
  NOR2_X1 U384 ( .A1(n605), .A2(n587), .ZN(n388) );
  XNOR2_X2 U385 ( .A(n642), .B(n641), .ZN(n741) );
  XOR2_X2 U386 ( .A(KEYINPUT62), .B(n652), .Z(n653) );
  XNOR2_X2 U387 ( .A(n365), .B(n356), .ZN(n381) );
  XNOR2_X2 U388 ( .A(n372), .B(KEYINPUT87), .ZN(n364) );
  NOR2_X2 U389 ( .A1(n622), .A2(n621), .ZN(n647) );
  NAND2_X1 U390 ( .A1(n423), .A2(n425), .ZN(n737) );
  NAND2_X1 U391 ( .A1(n390), .A2(n426), .ZN(n423) );
  XNOR2_X2 U392 ( .A(n637), .B(KEYINPUT59), .ZN(n638) );
  XNOR2_X2 U393 ( .A(KEYINPUT15), .B(G902), .ZN(n634) );
  XNOR2_X1 U394 ( .A(G137), .B(G128), .ZN(n510) );
  XNOR2_X1 U395 ( .A(G113), .B(G143), .ZN(n477) );
  NAND2_X2 U396 ( .A1(n423), .A2(n425), .ZN(n391) );
  XNOR2_X1 U397 ( .A(n526), .B(n405), .ZN(n404) );
  XNOR2_X2 U398 ( .A(n386), .B(G146), .ZN(n471) );
  NOR2_X2 U399 ( .A1(n585), .A2(n625), .ZN(n430) );
  NOR2_X1 U400 ( .A1(G953), .A2(G237), .ZN(n516) );
  NAND2_X1 U401 ( .A1(n552), .A2(n550), .ZN(n690) );
  XNOR2_X1 U402 ( .A(n735), .B(n734), .ZN(n347) );
  AND2_X1 U403 ( .A1(n624), .A2(n416), .ZN(n363) );
  NAND2_X1 U404 ( .A1(n555), .A2(n529), .ZN(n530) );
  XNOR2_X1 U405 ( .A(n401), .B(n400), .ZN(n535) );
  XNOR2_X1 U406 ( .A(n385), .B(n384), .ZN(n717) );
  XNOR2_X1 U407 ( .A(n586), .B(KEYINPUT38), .ZN(n688) );
  XNOR2_X1 U408 ( .A(n463), .B(n462), .ZN(n585) );
  XNOR2_X1 U409 ( .A(n437), .B(n350), .ZN(n700) );
  NOR2_X1 U410 ( .A1(n347), .A2(n736), .ZN(G63) );
  INV_X2 U411 ( .A(G125), .ZN(n386) );
  XNOR2_X1 U412 ( .A(n595), .B(n594), .ZN(n624) );
  INV_X1 U413 ( .A(KEYINPUT46), .ZN(n594) );
  NAND2_X1 U414 ( .A1(n635), .A2(n633), .ZN(n431) );
  AND2_X1 U415 ( .A1(n700), .A2(n438), .ZN(n579) );
  XNOR2_X1 U416 ( .A(n597), .B(n378), .ZN(n697) );
  INV_X1 U417 ( .A(KEYINPUT1), .ZN(n378) );
  NOR2_X1 U418 ( .A1(n647), .A2(n429), .ZN(n415) );
  INV_X1 U419 ( .A(KEYINPUT0), .ZN(n400) );
  AND2_X1 U420 ( .A1(n545), .A2(n556), .ZN(n534) );
  INV_X1 U421 ( .A(KEYINPUT41), .ZN(n384) );
  NOR2_X1 U422 ( .A1(n690), .A2(n625), .ZN(n383) );
  INV_X1 U423 ( .A(KEYINPUT39), .ZN(n387) );
  NAND2_X1 U424 ( .A1(n614), .A2(n366), .ZN(n522) );
  INV_X1 U425 ( .A(n374), .ZN(n376) );
  NAND2_X1 U426 ( .A1(n408), .A2(n461), .ZN(n379) );
  NOR2_X1 U427 ( .A1(n738), .A2(G902), .ZN(n437) );
  INV_X1 U428 ( .A(n697), .ZN(n626) );
  INV_X1 U429 ( .A(KEYINPUT48), .ZN(n429) );
  NOR2_X1 U430 ( .A1(n433), .A2(n411), .ZN(n410) );
  OR2_X1 U431 ( .A1(n434), .A2(n633), .ZN(n433) );
  NOR2_X1 U432 ( .A1(n634), .A2(KEYINPUT86), .ZN(n434) );
  NAND2_X1 U433 ( .A1(n634), .A2(KEYINPUT86), .ZN(n432) );
  XOR2_X1 U434 ( .A(KEYINPUT80), .B(KEYINPUT96), .Z(n448) );
  XNOR2_X1 U435 ( .A(G113), .B(KEYINPUT71), .ZN(n454) );
  XNOR2_X1 U436 ( .A(G119), .B(G116), .ZN(n453) );
  XOR2_X1 U437 ( .A(KEYINPUT11), .B(KEYINPUT99), .Z(n473) );
  XOR2_X1 U438 ( .A(KEYINPUT100), .B(KEYINPUT12), .Z(n476) );
  NAND2_X1 U439 ( .A1(n688), .A2(n375), .ZN(n692) );
  INV_X1 U440 ( .A(G237), .ZN(n460) );
  NOR2_X1 U441 ( .A1(n353), .A2(n700), .ZN(n590) );
  NOR2_X1 U442 ( .A1(n697), .A2(n698), .ZN(n545) );
  XNOR2_X1 U443 ( .A(n441), .B(n440), .ZN(n512) );
  XNOR2_X1 U444 ( .A(KEYINPUT68), .B(KEYINPUT8), .ZN(n440) );
  XNOR2_X1 U445 ( .A(n442), .B(KEYINPUT67), .ZN(n441) );
  NAND2_X1 U446 ( .A1(n749), .A2(G234), .ZN(n442) );
  XNOR2_X1 U447 ( .A(n397), .B(n368), .ZN(n758) );
  XNOR2_X1 U448 ( .A(KEYINPUT10), .B(G140), .ZN(n368) );
  XNOR2_X1 U449 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n370) );
  INV_X1 U450 ( .A(KEYINPUT102), .ZN(n421) );
  XNOR2_X1 U451 ( .A(KEYINPUT105), .B(KEYINPUT9), .ZN(n487) );
  NAND2_X1 U452 ( .A1(G237), .A2(G234), .ZN(n465) );
  INV_X1 U453 ( .A(KEYINPUT6), .ZN(n377) );
  XNOR2_X1 U454 ( .A(n371), .B(n367), .ZN(n738) );
  NAND2_X1 U455 ( .A1(n512), .A2(G221), .ZN(n371) );
  XNOR2_X1 U456 ( .A(n369), .B(n758), .ZN(n367) );
  XNOR2_X1 U457 ( .A(n511), .B(n370), .ZN(n369) );
  XNOR2_X1 U458 ( .A(n422), .B(n419), .ZN(n734) );
  XNOR2_X1 U459 ( .A(n491), .B(n420), .ZN(n419) );
  XNOR2_X1 U460 ( .A(n490), .B(n488), .ZN(n422) );
  XNOR2_X1 U461 ( .A(n489), .B(n421), .ZN(n420) );
  XNOR2_X1 U462 ( .A(n593), .B(n418), .ZN(n436) );
  INV_X1 U463 ( .A(KEYINPUT42), .ZN(n418) );
  NOR2_X1 U464 ( .A1(n717), .A2(n592), .ZN(n593) );
  NAND2_X1 U465 ( .A1(n376), .A2(n366), .ZN(n528) );
  XNOR2_X1 U466 ( .A(n530), .B(G110), .ZN(G12) );
  AND2_X1 U467 ( .A1(n364), .A2(n355), .ZN(n349) );
  INV_X1 U468 ( .A(n625), .ZN(n375) );
  XOR2_X1 U469 ( .A(n515), .B(n514), .Z(n350) );
  INV_X1 U470 ( .A(n701), .ZN(n439) );
  XNOR2_X1 U471 ( .A(G472), .B(KEYINPUT73), .ZN(n351) );
  XOR2_X1 U472 ( .A(G119), .B(G110), .Z(n352) );
  OR2_X1 U473 ( .A1(n589), .A2(n439), .ZN(n353) );
  XNOR2_X1 U474 ( .A(n613), .B(n612), .ZN(n623) );
  INV_X1 U475 ( .A(n623), .ZN(n362) );
  AND2_X1 U476 ( .A1(n646), .A2(n432), .ZN(n355) );
  XOR2_X1 U477 ( .A(n588), .B(KEYINPUT112), .Z(n356) );
  XOR2_X1 U478 ( .A(n497), .B(KEYINPUT22), .Z(n357) );
  INV_X1 U479 ( .A(G902), .ZN(n461) );
  NAND2_X1 U480 ( .A1(n432), .A2(KEYINPUT64), .ZN(n424) );
  INV_X1 U481 ( .A(n634), .ZN(n635) );
  INV_X1 U482 ( .A(G146), .ZN(n679) );
  NAND2_X1 U483 ( .A1(n360), .A2(n358), .ZN(n373) );
  NAND2_X1 U484 ( .A1(n362), .A2(n359), .ZN(n358) );
  AND2_X1 U485 ( .A1(n415), .A2(n624), .ZN(n359) );
  NAND2_X1 U486 ( .A1(n361), .A2(n429), .ZN(n360) );
  NAND2_X1 U487 ( .A1(n363), .A2(n362), .ZN(n361) );
  AND2_X1 U488 ( .A1(n364), .A2(n646), .ZN(n382) );
  NAND2_X1 U489 ( .A1(n632), .A2(n678), .ZN(n365) );
  XNOR2_X1 U490 ( .A(n388), .B(n387), .ZN(n632) );
  INV_X1 U491 ( .A(n700), .ZN(n366) );
  NOR2_X1 U492 ( .A1(n615), .A2(n376), .ZN(n591) );
  XNOR2_X1 U493 ( .A(n374), .B(n377), .ZN(n556) );
  XNOR2_X2 U494 ( .A(n379), .B(n509), .ZN(n597) );
  XNOR2_X1 U495 ( .A(n380), .B(G134), .ZN(n501) );
  XNOR2_X1 U496 ( .A(n380), .B(n443), .ZN(n444) );
  XNOR2_X2 U497 ( .A(G143), .B(G128), .ZN(n380) );
  XNOR2_X1 U498 ( .A(n381), .B(G131), .ZN(G33) );
  NAND2_X1 U499 ( .A1(n750), .A2(n382), .ZN(n435) );
  XNOR2_X1 U500 ( .A(n382), .B(n761), .ZN(n762) );
  NAND2_X1 U501 ( .A1(n688), .A2(n383), .ZN(n385) );
  NOR2_X1 U502 ( .A1(n414), .A2(n424), .ZN(n390) );
  AND2_X2 U503 ( .A1(n402), .A2(n354), .ZN(n414) );
  XNOR2_X1 U504 ( .A(n436), .B(G137), .ZN(G39) );
  NOR2_X1 U505 ( .A1(n652), .A2(G902), .ZN(n389) );
  NAND2_X1 U506 ( .A1(n750), .A2(n349), .ZN(n412) );
  BUF_X1 U507 ( .A(n404), .Z(n392) );
  NAND2_X1 U508 ( .A1(n445), .A2(n444), .ZN(n395) );
  NAND2_X1 U509 ( .A1(n393), .A2(n394), .ZN(n396) );
  NAND2_X1 U510 ( .A1(n396), .A2(n395), .ZN(n450) );
  INV_X1 U511 ( .A(n445), .ZN(n393) );
  INV_X1 U512 ( .A(n444), .ZN(n394) );
  XNOR2_X1 U513 ( .A(n679), .B(n348), .ZN(n397) );
  XNOR2_X1 U514 ( .A(n399), .B(n602), .ZN(n427) );
  AND2_X1 U515 ( .A1(n646), .A2(n431), .ZN(n398) );
  NAND2_X1 U516 ( .A1(n600), .A2(n601), .ZN(n399) );
  NOR2_X1 U517 ( .A1(n596), .A2(n470), .ZN(n401) );
  XNOR2_X1 U518 ( .A(n571), .B(KEYINPUT45), .ZN(n402) );
  BUF_X1 U519 ( .A(n770), .Z(n403) );
  XNOR2_X1 U520 ( .A(n571), .B(KEYINPUT45), .ZN(n750) );
  XNOR2_X1 U521 ( .A(n539), .B(n538), .ZN(n770) );
  INV_X1 U522 ( .A(n392), .ZN(n650) );
  XOR2_X1 U523 ( .A(n525), .B(KEYINPUT65), .Z(n405) );
  NOR2_X1 U524 ( .A1(n410), .A2(KEYINPUT64), .ZN(n409) );
  AND2_X2 U525 ( .A1(n413), .A2(n406), .ZN(n425) );
  NAND2_X1 U526 ( .A1(n412), .A2(n409), .ZN(n406) );
  XNOR2_X1 U527 ( .A(n407), .B(KEYINPUT34), .ZN(n536) );
  NOR2_X2 U528 ( .A1(n549), .A2(n718), .ZN(n407) );
  INV_X1 U529 ( .A(n729), .ZN(n408) );
  NAND2_X1 U530 ( .A1(n435), .A2(n433), .ZN(n426) );
  INV_X1 U531 ( .A(n432), .ZN(n411) );
  NAND2_X1 U532 ( .A1(n414), .A2(n636), .ZN(n413) );
  INV_X1 U533 ( .A(n647), .ZN(n416) );
  XNOR2_X1 U534 ( .A(n417), .B(n603), .ZN(n611) );
  NAND2_X1 U535 ( .A1(n427), .A2(n691), .ZN(n417) );
  NAND2_X1 U536 ( .A1(n427), .A2(n674), .ZN(n675) );
  NAND2_X1 U537 ( .A1(n427), .A2(n678), .ZN(n680) );
  INV_X1 U538 ( .A(n649), .ZN(n428) );
  XNOR2_X1 U539 ( .A(n430), .B(KEYINPUT92), .ZN(n618) );
  XNOR2_X1 U540 ( .A(n435), .B(n633), .ZN(n723) );
  NAND2_X1 U541 ( .A1(n700), .A2(n701), .ZN(n698) );
  NOR2_X1 U542 ( .A1(n589), .A2(n439), .ZN(n438) );
  INV_X4 U543 ( .A(G953), .ZN(n749) );
  BUF_X1 U544 ( .A(n527), .Z(n555) );
  INV_X1 U545 ( .A(KEYINPUT77), .ZN(n612) );
  XNOR2_X1 U546 ( .A(n532), .B(n531), .ZN(n563) );
  XNOR2_X1 U547 ( .A(n534), .B(n533), .ZN(n718) );
  INV_X1 U548 ( .A(KEYINPUT84), .ZN(n602) );
  XNOR2_X1 U549 ( .A(n537), .B(KEYINPUT81), .ZN(n538) );
  INV_X1 U550 ( .A(KEYINPUT60), .ZN(n644) );
  XNOR2_X2 U551 ( .A(KEYINPUT66), .B(G101), .ZN(n502) );
  XNOR2_X1 U552 ( .A(n471), .B(n502), .ZN(n445) );
  XNOR2_X1 U553 ( .A(KEYINPUT17), .B(KEYINPUT4), .ZN(n443) );
  NAND2_X1 U554 ( .A1(G224), .A2(n749), .ZN(n446) );
  XNOR2_X1 U555 ( .A(n446), .B(KEYINPUT18), .ZN(n447) );
  XNOR2_X1 U556 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U557 ( .A(n450), .B(n449), .ZN(n452) );
  XOR2_X1 U558 ( .A(G110), .B(G104), .Z(n451) );
  XNOR2_X1 U559 ( .A(n451), .B(G107), .ZN(n744) );
  XNOR2_X1 U560 ( .A(n744), .B(KEYINPUT72), .ZN(n506) );
  XNOR2_X1 U561 ( .A(n452), .B(n506), .ZN(n459) );
  XNOR2_X1 U562 ( .A(n453), .B(KEYINPUT3), .ZN(n455) );
  XNOR2_X1 U563 ( .A(n455), .B(n454), .ZN(n519) );
  XNOR2_X1 U564 ( .A(KEYINPUT76), .B(KEYINPUT16), .ZN(n457) );
  XNOR2_X1 U565 ( .A(G122), .B(KEYINPUT75), .ZN(n456) );
  XNOR2_X1 U566 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U567 ( .A(n519), .B(n458), .ZN(n745) );
  XNOR2_X1 U568 ( .A(n459), .B(n745), .ZN(n658) );
  NAND2_X1 U569 ( .A1(n658), .A2(n634), .ZN(n463) );
  NAND2_X1 U570 ( .A1(n461), .A2(n460), .ZN(n464) );
  NAND2_X1 U571 ( .A1(n464), .A2(G210), .ZN(n462) );
  AND2_X1 U572 ( .A1(n464), .A2(G214), .ZN(n625) );
  XNOR2_X1 U573 ( .A(n618), .B(KEYINPUT19), .ZN(n596) );
  XNOR2_X1 U574 ( .A(n465), .B(KEYINPUT14), .ZN(n714) );
  NAND2_X1 U575 ( .A1(n749), .A2(G952), .ZN(n575) );
  INV_X1 U576 ( .A(G898), .ZN(n467) );
  NAND2_X1 U577 ( .A1(G953), .A2(G902), .ZN(n572) );
  INV_X1 U578 ( .A(n572), .ZN(n466) );
  NAND2_X1 U579 ( .A1(n467), .A2(n466), .ZN(n468) );
  NAND2_X1 U580 ( .A1(n575), .A2(n468), .ZN(n469) );
  NAND2_X1 U581 ( .A1(n714), .A2(n469), .ZN(n470) );
  XNOR2_X1 U582 ( .A(KEYINPUT101), .B(KEYINPUT13), .ZN(n483) );
  NAND2_X1 U583 ( .A1(n516), .A2(G214), .ZN(n472) );
  XNOR2_X1 U584 ( .A(n473), .B(n472), .ZN(n474) );
  XOR2_X1 U585 ( .A(n474), .B(G131), .Z(n480) );
  XNOR2_X1 U586 ( .A(G104), .B(G122), .ZN(n475) );
  XNOR2_X1 U587 ( .A(n476), .B(n475), .ZN(n478) );
  XNOR2_X1 U588 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U589 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U590 ( .A(n758), .B(n481), .ZN(n637) );
  NOR2_X1 U591 ( .A1(G902), .A2(n637), .ZN(n482) );
  XNOR2_X1 U592 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U593 ( .A(n484), .B(G475), .ZN(n552) );
  XOR2_X1 U594 ( .A(KEYINPUT7), .B(KEYINPUT103), .Z(n486) );
  XNOR2_X1 U595 ( .A(G107), .B(KEYINPUT104), .ZN(n485) );
  XNOR2_X1 U596 ( .A(n486), .B(n485), .ZN(n491) );
  NAND2_X1 U597 ( .A1(G217), .A2(n512), .ZN(n490) );
  XNOR2_X1 U598 ( .A(n501), .B(n487), .ZN(n488) );
  XNOR2_X1 U599 ( .A(G116), .B(G122), .ZN(n489) );
  NOR2_X1 U600 ( .A1(G902), .A2(n734), .ZN(n492) );
  XNOR2_X1 U601 ( .A(G478), .B(n492), .ZN(n550) );
  XOR2_X1 U602 ( .A(KEYINPUT20), .B(KEYINPUT97), .Z(n494) );
  NAND2_X1 U603 ( .A1(G234), .A2(n634), .ZN(n493) );
  XNOR2_X1 U604 ( .A(n494), .B(n493), .ZN(n513) );
  AND2_X1 U605 ( .A1(n513), .A2(G221), .ZN(n495) );
  XNOR2_X1 U606 ( .A(n495), .B(KEYINPUT21), .ZN(n701) );
  OR2_X1 U607 ( .A1(n690), .A2(n439), .ZN(n496) );
  NOR2_X2 U608 ( .A1(n535), .A2(n496), .ZN(n498) );
  INV_X1 U609 ( .A(KEYINPUT74), .ZN(n497) );
  XNOR2_X1 U610 ( .A(n498), .B(n357), .ZN(n527) );
  XNOR2_X1 U611 ( .A(KEYINPUT4), .B(G137), .ZN(n499) );
  XNOR2_X1 U612 ( .A(n499), .B(G131), .ZN(n500) );
  XNOR2_X1 U613 ( .A(n502), .B(n679), .ZN(n503) );
  INV_X1 U614 ( .A(n521), .ZN(n508) );
  NAND2_X1 U615 ( .A1(n749), .A2(G227), .ZN(n504) );
  XNOR2_X1 U616 ( .A(n504), .B(G140), .ZN(n505) );
  XNOR2_X1 U617 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U618 ( .A(n508), .B(n507), .ZN(n729) );
  XNOR2_X1 U619 ( .A(KEYINPUT70), .B(G469), .ZN(n509) );
  XNOR2_X1 U620 ( .A(n697), .B(KEYINPUT94), .ZN(n621) );
  XNOR2_X1 U621 ( .A(n352), .B(n510), .ZN(n511) );
  XOR2_X1 U622 ( .A(KEYINPUT25), .B(KEYINPUT98), .Z(n515) );
  NAND2_X1 U623 ( .A1(n513), .A2(G217), .ZN(n514) );
  NAND2_X1 U624 ( .A1(n516), .A2(G210), .ZN(n517) );
  XNOR2_X1 U625 ( .A(n517), .B(KEYINPUT5), .ZN(n518) );
  XNOR2_X1 U626 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U627 ( .A(n521), .B(n520), .ZN(n652) );
  INV_X1 U628 ( .A(n556), .ZN(n614) );
  OR2_X1 U629 ( .A1(n621), .A2(n522), .ZN(n523) );
  XNOR2_X1 U630 ( .A(n523), .B(KEYINPUT83), .ZN(n524) );
  NAND2_X1 U631 ( .A1(n527), .A2(n524), .ZN(n526) );
  XNOR2_X1 U632 ( .A(KEYINPUT82), .B(KEYINPUT32), .ZN(n525) );
  NOR2_X1 U633 ( .A1(n528), .A2(n626), .ZN(n529) );
  NAND2_X1 U634 ( .A1(n404), .A2(n530), .ZN(n532) );
  INV_X1 U635 ( .A(KEYINPUT91), .ZN(n531) );
  XOR2_X1 U636 ( .A(KEYINPUT107), .B(KEYINPUT33), .Z(n533) );
  BUF_X2 U637 ( .A(n535), .Z(n549) );
  NOR2_X1 U638 ( .A1(n552), .A2(n550), .ZN(n606) );
  NAND2_X1 U639 ( .A1(n536), .A2(n606), .ZN(n539) );
  INV_X1 U640 ( .A(KEYINPUT35), .ZN(n537) );
  NAND2_X1 U641 ( .A1(n770), .A2(KEYINPUT90), .ZN(n540) );
  NAND2_X1 U642 ( .A1(n540), .A2(KEYINPUT44), .ZN(n541) );
  NOR2_X1 U643 ( .A1(n563), .A2(n541), .ZN(n544) );
  INV_X1 U644 ( .A(KEYINPUT90), .ZN(n542) );
  NOR2_X1 U645 ( .A1(n542), .A2(KEYINPUT44), .ZN(n543) );
  NOR2_X1 U646 ( .A1(n544), .A2(n543), .ZN(n562) );
  NAND2_X1 U647 ( .A1(n545), .A2(n374), .ZN(n707) );
  NOR2_X1 U648 ( .A1(n549), .A2(n707), .ZN(n546) );
  XNOR2_X1 U649 ( .A(n546), .B(KEYINPUT31), .ZN(n685) );
  NOR2_X1 U650 ( .A1(n698), .A2(n374), .ZN(n547) );
  NAND2_X1 U651 ( .A1(n547), .A2(n597), .ZN(n548) );
  OR2_X1 U652 ( .A1(n549), .A2(n548), .ZN(n670) );
  NAND2_X1 U653 ( .A1(n685), .A2(n670), .ZN(n553) );
  INV_X1 U654 ( .A(n550), .ZN(n551) );
  AND2_X1 U655 ( .A1(n552), .A2(n551), .ZN(n674) );
  INV_X1 U656 ( .A(n674), .ZN(n686) );
  OR2_X1 U657 ( .A1(n552), .A2(n551), .ZN(n681) );
  NAND2_X1 U658 ( .A1(n686), .A2(n681), .ZN(n691) );
  NAND2_X1 U659 ( .A1(n553), .A2(n691), .ZN(n554) );
  XNOR2_X1 U660 ( .A(n554), .B(KEYINPUT106), .ZN(n560) );
  NOR2_X1 U661 ( .A1(n626), .A2(n556), .ZN(n557) );
  NAND2_X1 U662 ( .A1(n555), .A2(n557), .ZN(n558) );
  XNOR2_X1 U663 ( .A(n558), .B(KEYINPUT89), .ZN(n559) );
  NAND2_X1 U664 ( .A1(n559), .A2(n700), .ZN(n668) );
  NAND2_X1 U665 ( .A1(n560), .A2(n668), .ZN(n561) );
  NOR2_X1 U666 ( .A1(n562), .A2(n561), .ZN(n570) );
  INV_X1 U667 ( .A(n563), .ZN(n565) );
  INV_X1 U668 ( .A(KEYINPUT44), .ZN(n564) );
  NAND2_X1 U669 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U670 ( .A1(n566), .A2(KEYINPUT90), .ZN(n568) );
  INV_X1 U671 ( .A(n403), .ZN(n567) );
  NAND2_X1 U672 ( .A1(n568), .A2(n567), .ZN(n569) );
  NAND2_X1 U673 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U674 ( .A1(G900), .A2(n572), .ZN(n573) );
  NAND2_X1 U675 ( .A1(n714), .A2(n573), .ZN(n574) );
  XOR2_X1 U676 ( .A(KEYINPUT108), .B(n574), .Z(n578) );
  INV_X1 U677 ( .A(n714), .ZN(n576) );
  NOR2_X1 U678 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U679 ( .A1(n578), .A2(n577), .ZN(n589) );
  NAND2_X1 U680 ( .A1(n579), .A2(n597), .ZN(n583) );
  XOR2_X1 U681 ( .A(KEYINPUT110), .B(KEYINPUT30), .Z(n580) );
  XNOR2_X1 U682 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U683 ( .A(n584), .B(KEYINPUT79), .ZN(n605) );
  BUF_X1 U684 ( .A(n585), .Z(n586) );
  INV_X1 U685 ( .A(n688), .ZN(n587) );
  INV_X1 U686 ( .A(n681), .ZN(n678) );
  XNOR2_X1 U687 ( .A(KEYINPUT113), .B(KEYINPUT40), .ZN(n588) );
  XNOR2_X1 U688 ( .A(n590), .B(KEYINPUT69), .ZN(n615) );
  XNOR2_X1 U689 ( .A(n591), .B(KEYINPUT28), .ZN(n601) );
  NAND2_X1 U690 ( .A1(n601), .A2(n597), .ZN(n592) );
  BUF_X1 U691 ( .A(n596), .Z(n599) );
  INV_X1 U692 ( .A(n597), .ZN(n598) );
  NOR2_X1 U693 ( .A1(n599), .A2(n598), .ZN(n600) );
  INV_X1 U694 ( .A(KEYINPUT78), .ZN(n604) );
  NOR2_X1 U695 ( .A1(n604), .A2(KEYINPUT47), .ZN(n603) );
  NAND2_X1 U696 ( .A1(n604), .A2(KEYINPUT47), .ZN(n609) );
  INV_X1 U697 ( .A(n586), .ZN(n630) );
  NAND2_X1 U698 ( .A1(n606), .A2(n630), .ZN(n607) );
  NOR2_X1 U699 ( .A1(n605), .A2(n607), .ZN(n608) );
  XNOR2_X1 U700 ( .A(n608), .B(KEYINPUT111), .ZN(n771) );
  AND2_X1 U701 ( .A1(n609), .A2(n771), .ZN(n610) );
  NAND2_X1 U702 ( .A1(n611), .A2(n610), .ZN(n613) );
  XNOR2_X1 U703 ( .A(n616), .B(KEYINPUT109), .ZN(n617) );
  BUF_X1 U704 ( .A(n618), .Z(n619) );
  NAND2_X1 U705 ( .A1(n628), .A2(n619), .ZN(n620) );
  XNOR2_X1 U706 ( .A(n620), .B(KEYINPUT36), .ZN(n622) );
  NOR2_X1 U707 ( .A1(n626), .A2(n625), .ZN(n627) );
  NAND2_X1 U708 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U709 ( .A(KEYINPUT43), .B(n629), .Z(n631) );
  NOR2_X1 U710 ( .A1(n631), .A2(n630), .ZN(n649) );
  NAND2_X1 U711 ( .A1(n632), .A2(n674), .ZN(n646) );
  INV_X1 U712 ( .A(KEYINPUT2), .ZN(n633) );
  INV_X1 U713 ( .A(KEYINPUT64), .ZN(n636) );
  NAND2_X1 U714 ( .A1(n737), .A2(G475), .ZN(n639) );
  XNOR2_X1 U715 ( .A(n639), .B(n638), .ZN(n643) );
  INV_X1 U716 ( .A(G952), .ZN(n640) );
  NAND2_X1 U717 ( .A1(n640), .A2(G953), .ZN(n642) );
  INV_X1 U718 ( .A(KEYINPUT95), .ZN(n641) );
  NAND2_X1 U719 ( .A1(n643), .A2(n741), .ZN(n645) );
  XNOR2_X1 U720 ( .A(n645), .B(n644), .ZN(G60) );
  XNOR2_X1 U721 ( .A(n646), .B(G134), .ZN(G36) );
  XOR2_X1 U722 ( .A(n348), .B(KEYINPUT37), .Z(n648) );
  XOR2_X1 U723 ( .A(n648), .B(n647), .Z(G27) );
  XOR2_X1 U724 ( .A(G140), .B(n649), .Z(G42) );
  XNOR2_X1 U725 ( .A(G119), .B(KEYINPUT127), .ZN(n651) );
  XNOR2_X1 U726 ( .A(n650), .B(n651), .ZN(G21) );
  NAND2_X1 U727 ( .A1(n391), .A2(G472), .ZN(n654) );
  XNOR2_X1 U728 ( .A(n654), .B(n653), .ZN(n655) );
  NAND2_X1 U729 ( .A1(n655), .A2(n741), .ZN(n657) );
  XOR2_X1 U730 ( .A(KEYINPUT93), .B(KEYINPUT63), .Z(n656) );
  XNOR2_X1 U731 ( .A(n657), .B(n656), .ZN(G57) );
  NAND2_X1 U732 ( .A1(n391), .A2(G210), .ZN(n663) );
  BUF_X1 U733 ( .A(n658), .Z(n659) );
  XNOR2_X1 U734 ( .A(KEYINPUT85), .B(KEYINPUT54), .ZN(n660) );
  XNOR2_X1 U735 ( .A(n660), .B(KEYINPUT55), .ZN(n661) );
  XNOR2_X1 U736 ( .A(n663), .B(n662), .ZN(n664) );
  NAND2_X1 U737 ( .A1(n664), .A2(n741), .ZN(n667) );
  XOR2_X1 U738 ( .A(KEYINPUT118), .B(KEYINPUT56), .Z(n665) );
  XNOR2_X1 U739 ( .A(n665), .B(KEYINPUT88), .ZN(n666) );
  XNOR2_X1 U740 ( .A(n667), .B(n666), .ZN(G51) );
  XNOR2_X1 U741 ( .A(G101), .B(n668), .ZN(G3) );
  NOR2_X1 U742 ( .A1(n681), .A2(n670), .ZN(n669) );
  XOR2_X1 U743 ( .A(G104), .B(n669), .Z(G6) );
  NOR2_X1 U744 ( .A1(n686), .A2(n670), .ZN(n672) );
  XNOR2_X1 U745 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n671) );
  XNOR2_X1 U746 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U747 ( .A(G107), .B(n673), .ZN(G9) );
  XOR2_X1 U748 ( .A(KEYINPUT29), .B(KEYINPUT114), .Z(n676) );
  XNOR2_X1 U749 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U750 ( .A(G128), .B(n677), .ZN(G30) );
  XNOR2_X1 U751 ( .A(n680), .B(G146), .ZN(G48) );
  NOR2_X1 U752 ( .A1(n681), .A2(n685), .ZN(n683) );
  XNOR2_X1 U753 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n682) );
  XNOR2_X1 U754 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U755 ( .A(G113), .B(n684), .ZN(G15) );
  NOR2_X1 U756 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U757 ( .A(G116), .B(n687), .Z(G18) );
  NOR2_X1 U758 ( .A1(n688), .A2(n375), .ZN(n689) );
  NOR2_X1 U759 ( .A1(n690), .A2(n689), .ZN(n695) );
  INV_X1 U760 ( .A(n691), .ZN(n693) );
  NOR2_X1 U761 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U762 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U763 ( .A1(n696), .A2(n718), .ZN(n712) );
  NAND2_X1 U764 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U765 ( .A(n699), .B(KEYINPUT50), .ZN(n706) );
  NOR2_X1 U766 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U767 ( .A(KEYINPUT49), .B(n702), .Z(n704) );
  NOR2_X1 U768 ( .A1(n704), .A2(n374), .ZN(n705) );
  NAND2_X1 U769 ( .A1(n706), .A2(n705), .ZN(n708) );
  NAND2_X1 U770 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U771 ( .A(KEYINPUT51), .B(n709), .ZN(n710) );
  NOR2_X1 U772 ( .A1(n717), .A2(n710), .ZN(n711) );
  NOR2_X1 U773 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U774 ( .A(KEYINPUT52), .B(n713), .ZN(n716) );
  NAND2_X1 U775 ( .A1(n714), .A2(G952), .ZN(n715) );
  NOR2_X1 U776 ( .A1(n716), .A2(n715), .ZN(n721) );
  NOR2_X1 U777 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U778 ( .A(n719), .B(KEYINPUT117), .Z(n720) );
  NOR2_X1 U779 ( .A1(n721), .A2(n720), .ZN(n722) );
  AND2_X1 U780 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U781 ( .A1(n749), .A2(n724), .ZN(n725) );
  XOR2_X1 U782 ( .A(KEYINPUT53), .B(n725), .Z(G75) );
  INV_X1 U783 ( .A(n741), .ZN(n736) );
  BUF_X1 U784 ( .A(n391), .Z(n726) );
  NAND2_X1 U785 ( .A1(n726), .A2(G469), .ZN(n732) );
  XOR2_X1 U786 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n728) );
  XNOR2_X1 U787 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n727) );
  XNOR2_X1 U788 ( .A(n728), .B(n727), .ZN(n730) );
  XOR2_X1 U789 ( .A(n730), .B(n729), .Z(n731) );
  XNOR2_X1 U790 ( .A(n732), .B(n731), .ZN(n733) );
  NOR2_X1 U791 ( .A1(n733), .A2(n736), .ZN(G54) );
  NAND2_X1 U792 ( .A1(n726), .A2(G478), .ZN(n735) );
  NAND2_X1 U793 ( .A1(n737), .A2(G217), .ZN(n740) );
  INV_X1 U794 ( .A(n738), .ZN(n739) );
  XNOR2_X1 U795 ( .A(n740), .B(n739), .ZN(n742) );
  NAND2_X1 U796 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U797 ( .A(n743), .B(KEYINPUT121), .ZN(G66) );
  XOR2_X1 U798 ( .A(n744), .B(G101), .Z(n746) );
  XNOR2_X1 U799 ( .A(n746), .B(n745), .ZN(n748) );
  NOR2_X1 U800 ( .A1(G898), .A2(n749), .ZN(n747) );
  NOR2_X1 U801 ( .A1(n748), .A2(n747), .ZN(n757) );
  AND2_X1 U802 ( .A1(n402), .A2(n749), .ZN(n754) );
  NAND2_X1 U803 ( .A1(G953), .A2(G224), .ZN(n751) );
  XOR2_X1 U804 ( .A(KEYINPUT61), .B(n751), .Z(n752) );
  NOR2_X1 U805 ( .A1(n467), .A2(n752), .ZN(n753) );
  NOR2_X1 U806 ( .A1(n754), .A2(n753), .ZN(n755) );
  XOR2_X1 U807 ( .A(n755), .B(KEYINPUT122), .Z(n756) );
  XNOR2_X1 U808 ( .A(n757), .B(n756), .ZN(G69) );
  XNOR2_X1 U809 ( .A(n758), .B(KEYINPUT123), .ZN(n759) );
  XOR2_X1 U810 ( .A(n760), .B(n759), .Z(n764) );
  XNOR2_X1 U811 ( .A(n764), .B(KEYINPUT124), .ZN(n761) );
  NOR2_X1 U812 ( .A1(n762), .A2(G953), .ZN(n763) );
  XNOR2_X1 U813 ( .A(KEYINPUT125), .B(n763), .ZN(n768) );
  XNOR2_X1 U814 ( .A(G227), .B(n764), .ZN(n765) );
  NAND2_X1 U815 ( .A1(n765), .A2(G900), .ZN(n766) );
  NAND2_X1 U816 ( .A1(n766), .A2(G953), .ZN(n767) );
  NAND2_X1 U817 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U818 ( .A(n769), .B(KEYINPUT126), .ZN(G72) );
  XOR2_X1 U819 ( .A(n403), .B(G122), .Z(G24) );
  XNOR2_X1 U820 ( .A(G143), .B(n771), .ZN(G45) );
endmodule

