//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 1 1 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n560, new_n562, new_n563, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n614, new_n617, new_n619,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT64), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n464));
  XNOR2_X1  g039(.A(new_n463), .B(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(G2105), .B1(new_n465), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  AND2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  OAI211_X1 g050(.A(G137), .B(new_n473), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT66), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n468), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G101), .ZN(new_n479));
  AND3_X1   g054(.A1(new_n476), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n477), .B1(new_n476), .B2(new_n479), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n472), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  AOI21_X1  g058(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT67), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n473), .B1(new_n469), .B2(new_n470), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT68), .ZN(new_n489));
  INV_X1    g064(.A(G100), .ZN(new_n490));
  AND3_X1   g065(.A1(new_n490), .A2(new_n473), .A3(KEYINPUT69), .ZN(new_n491));
  AOI21_X1  g066(.A(KEYINPUT69), .B1(new_n490), .B2(new_n473), .ZN(new_n492));
  OAI221_X1 g067(.A(G2104), .B1(G112), .B2(new_n473), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  AND3_X1   g068(.A1(new_n486), .A2(new_n489), .A3(new_n493), .ZN(G162));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n496), .B1(new_n474), .B2(new_n475), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n497), .A2(KEYINPUT70), .A3(new_n498), .ZN(new_n499));
  OAI211_X1 g074(.A(G126), .B(G2105), .C1(new_n474), .C2(new_n475), .ZN(new_n500));
  OR2_X1    g075(.A1(G102), .A2(G2105), .ZN(new_n501));
  INV_X1    g076(.A(G114), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G2105), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n501), .A2(new_n503), .A3(G2104), .ZN(new_n504));
  AND2_X1   g079(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n473), .A2(G138), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n506), .B1(new_n469), .B2(new_n470), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT4), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI211_X1 g084(.A(new_n496), .B(new_n508), .C1(new_n475), .C2(new_n474), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  OAI211_X1 g086(.A(new_n499), .B(new_n505), .C1(new_n509), .C2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  OR2_X1    g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT72), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n519), .B(new_n520), .ZN(new_n521));
  OAI21_X1  g096(.A(KEYINPUT71), .B1(new_n518), .B2(KEYINPUT6), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT71), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT6), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(new_n524), .A3(G651), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n522), .A2(new_n525), .B1(KEYINPUT6), .B2(new_n518), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(new_n516), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n526), .A2(G543), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n528), .A2(G88), .B1(new_n529), .B2(G50), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n521), .A2(new_n530), .ZN(G303));
  INV_X1    g106(.A(G303), .ZN(G166));
  XNOR2_X1  g107(.A(KEYINPUT73), .B(KEYINPUT7), .ZN(new_n533));
  AND3_X1   g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n534), .ZN(new_n536));
  AND2_X1   g111(.A1(G63), .A2(G651), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n535), .A2(new_n536), .B1(new_n516), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n526), .A2(G51), .A3(G543), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n526), .A2(G89), .A3(new_n516), .ZN(new_n540));
  AND3_X1   g115(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(G168));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n514), .A2(new_n515), .ZN(new_n543));
  INV_X1    g118(.A(G64), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G651), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n526), .A2(G90), .A3(new_n516), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n526), .A2(G52), .A3(G543), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G56), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n543), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G651), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n526), .A2(G81), .A3(new_n516), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n526), .A2(G43), .A3(G543), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n560));
  XOR2_X1   g135(.A(new_n560), .B(KEYINPUT74), .Z(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n529), .A2(new_n565), .A3(G53), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n526), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G53), .ZN(new_n568));
  OAI21_X1  g143(.A(KEYINPUT9), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n516), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n571), .A2(new_n518), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n572), .B1(G91), .B2(new_n528), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n570), .A2(new_n573), .ZN(G299));
  NAND3_X1  g149(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(G286));
  OAI21_X1  g150(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(KEYINPUT75), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n578));
  OAI211_X1 g153(.A(new_n578), .B(G651), .C1(new_n516), .C2(G74), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n526), .A2(G49), .A3(G543), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n526), .A2(G87), .A3(new_n516), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(G288));
  NAND3_X1  g158(.A1(new_n526), .A2(G48), .A3(G543), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(KEYINPUT77), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n526), .A2(G86), .A3(new_n516), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  XOR2_X1   g162(.A(new_n587), .B(KEYINPUT76), .Z(new_n588));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n589), .B1(new_n514), .B2(new_n515), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT77), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n526), .A2(new_n592), .A3(G48), .A4(G543), .ZN(new_n593));
  NAND4_X1  g168(.A1(new_n585), .A2(new_n586), .A3(new_n591), .A4(new_n593), .ZN(G305));
  NAND2_X1  g169(.A1(new_n528), .A2(G85), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n529), .A2(G47), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  OAI211_X1 g172(.A(new_n595), .B(new_n596), .C1(new_n518), .C2(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n528), .A2(KEYINPUT10), .A3(G92), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  INV_X1    g176(.A(G92), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n527), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n543), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n529), .A2(G54), .B1(new_n607), .B2(G651), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n599), .B1(new_n610), .B2(G868), .ZN(G284));
  OAI21_X1  g186(.A(new_n599), .B1(new_n610), .B2(G868), .ZN(G321));
  INV_X1    g187(.A(G868), .ZN(new_n613));
  NAND2_X1  g188(.A1(G299), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(new_n613), .B2(G168), .ZN(G297));
  OAI21_X1  g190(.A(new_n614), .B1(new_n613), .B2(G168), .ZN(G280));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n610), .B1(new_n617), .B2(G860), .ZN(G148));
  NOR2_X1   g193(.A1(new_n558), .A2(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n610), .A2(new_n617), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G868), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT78), .Z(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n469), .A2(new_n470), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(new_n478), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT79), .B(G2100), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n484), .A2(G135), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n487), .A2(G123), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n473), .A2(G111), .ZN(new_n632));
  OAI21_X1  g207(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n633));
  OAI211_X1 g208(.A(new_n630), .B(new_n631), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT80), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2096), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n629), .A2(new_n636), .ZN(G156));
  XNOR2_X1  g212(.A(G2427), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(KEYINPUT14), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2443), .B(G2446), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2451), .B(G2454), .Z(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n645), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(G14), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n649), .A2(new_n650), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(KEYINPUT82), .ZN(new_n654));
  INV_X1    g229(.A(KEYINPUT82), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n655), .B1(new_n649), .B2(new_n650), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n652), .B1(new_n654), .B2(new_n656), .ZN(G401));
  XOR2_X1   g232(.A(KEYINPUT83), .B(KEYINPUT18), .Z(new_n658));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(KEYINPUT17), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n659), .A2(new_n660), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n658), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  INV_X1    g240(.A(new_n658), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n665), .B1(new_n661), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n664), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2096), .B(G2100), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT84), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n668), .B(new_n670), .ZN(G227));
  XOR2_X1   g246(.A(KEYINPUT85), .B(KEYINPUT19), .Z(new_n672));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1956), .B(G2474), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1961), .B(G1966), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT20), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n675), .A2(new_n676), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n680), .A2(new_n677), .ZN(new_n682));
  OAI211_X1 g257(.A(new_n679), .B(new_n681), .C1(new_n674), .C2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1991), .B(G1996), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1981), .B(G1986), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(G229));
  INV_X1    g265(.A(G29), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G32), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n478), .A2(G105), .ZN(new_n693));
  NAND3_X1  g268(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT26), .ZN(new_n695));
  AOI211_X1 g270(.A(new_n693), .B(new_n695), .C1(G141), .C2(new_n484), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n487), .A2(G129), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT91), .ZN(new_n698));
  AND2_X1   g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n692), .B1(new_n699), .B2(new_n691), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT27), .B(G1996), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G5), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G171), .B2(new_n704), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n703), .B1(G1961), .B2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(G2084), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT24), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n691), .B1(new_n709), .B2(G34), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n710), .A2(KEYINPUT90), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n709), .A2(G34), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(new_n710), .B2(KEYINPUT90), .ZN(new_n713));
  OAI22_X1  g288(.A1(new_n482), .A2(new_n691), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n707), .B1(new_n708), .B2(new_n714), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT94), .Z(new_n716));
  NAND2_X1  g291(.A1(new_n691), .A2(G26), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT28), .Z(new_n718));
  NAND2_X1  g293(.A1(new_n487), .A2(G128), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT88), .ZN(new_n720));
  OAI21_X1  g295(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n721));
  INV_X1    g296(.A(G116), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(G2105), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n484), .B2(G140), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n718), .B1(new_n725), .B2(G29), .ZN(new_n726));
  INV_X1    g301(.A(G2067), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(G29), .A2(G33), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT25), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n624), .A2(G127), .ZN(new_n732));
  NAND2_X1  g307(.A1(G115), .A2(G2104), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n473), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AOI211_X1 g309(.A(new_n731), .B(new_n734), .C1(G139), .C2(new_n484), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n729), .B1(new_n735), .B2(G29), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT89), .B(G2072), .Z(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT31), .B(G11), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n634), .B2(new_n691), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT92), .B(G28), .ZN(new_n741));
  AOI21_X1  g316(.A(G29), .B1(new_n741), .B2(KEYINPUT30), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n742), .A2(KEYINPUT93), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n741), .A2(KEYINPUT30), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n742), .B2(KEYINPUT93), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n740), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n738), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n736), .A2(new_n737), .ZN(new_n748));
  NOR3_X1   g323(.A1(new_n728), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n704), .A2(G20), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT23), .Z(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G299), .B2(G16), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G1956), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n704), .A2(G21), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G168), .B2(new_n704), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G1966), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n558), .A2(G16), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G16), .B2(G19), .ZN(new_n758));
  INV_X1    g333(.A(G1341), .ZN(new_n759));
  OAI22_X1  g334(.A1(new_n758), .A2(new_n759), .B1(new_n708), .B2(new_n714), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n758), .A2(new_n759), .B1(G1961), .B2(new_n706), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n749), .A2(new_n753), .A3(new_n761), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n691), .A2(G35), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G162), .B2(new_n691), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT29), .ZN(new_n766));
  INV_X1    g341(.A(G2090), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n610), .A2(G16), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G4), .B2(G16), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT87), .B(G1348), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n700), .A2(new_n702), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n691), .A2(G27), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G164), .B2(new_n691), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G2078), .ZN(new_n777));
  NOR3_X1   g352(.A1(new_n773), .A2(new_n774), .A3(new_n777), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n768), .A2(new_n772), .A3(new_n778), .ZN(new_n779));
  NOR3_X1   g354(.A1(new_n716), .A2(new_n763), .A3(new_n779), .ZN(new_n780));
  OR2_X1    g355(.A1(G16), .A2(G22), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G303), .B2(new_n704), .ZN(new_n782));
  INV_X1    g357(.A(G1971), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n704), .A2(G23), .ZN(new_n785));
  INV_X1    g360(.A(G288), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n785), .B1(new_n786), .B2(new_n704), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT33), .B(G1976), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  OR2_X1    g364(.A1(G6), .A2(G16), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G305), .B2(new_n704), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT32), .B(G1981), .Z(new_n792));
  AOI22_X1  g367(.A1(new_n782), .A2(new_n783), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n784), .A2(new_n789), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(KEYINPUT34), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(KEYINPUT34), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n484), .A2(G131), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n487), .A2(G119), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n473), .A2(G107), .ZN(new_n800));
  OAI21_X1  g375(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n798), .B(new_n799), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  MUX2_X1   g377(.A(G25), .B(new_n802), .S(G29), .Z(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT35), .B(G1991), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n803), .B(new_n804), .Z(new_n805));
  INV_X1    g380(.A(G1986), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n704), .A2(G24), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G290), .B2(G16), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n805), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n806), .B2(new_n808), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n796), .A2(new_n797), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(KEYINPUT86), .A2(KEYINPUT36), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OR2_X1    g388(.A1(KEYINPUT86), .A2(KEYINPUT36), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n811), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n780), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(G311));
  INV_X1    g392(.A(KEYINPUT95), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n816), .B(new_n818), .ZN(G150));
  NOR2_X1   g394(.A1(new_n609), .A2(new_n617), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n526), .A2(G93), .A3(new_n516), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n824));
  INV_X1    g399(.A(G55), .ZN(new_n825));
  OAI221_X1 g400(.A(new_n823), .B1(new_n824), .B2(new_n518), .C1(new_n567), .C2(new_n825), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n826), .A2(new_n557), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n826), .A2(new_n557), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n822), .B(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(KEYINPUT39), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT97), .ZN(new_n832));
  INV_X1    g407(.A(G860), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(new_n830), .B2(KEYINPUT39), .ZN(new_n834));
  AOI21_X1  g409(.A(KEYINPUT37), .B1(new_n826), .B2(G860), .ZN(new_n835));
  AND3_X1   g410(.A1(new_n826), .A2(KEYINPUT37), .A3(G860), .ZN(new_n836));
  OAI22_X1  g411(.A1(new_n832), .A2(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT98), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(G145));
  XNOR2_X1  g414(.A(new_n482), .B(new_n634), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(G162), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n725), .B(G164), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(new_n699), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n735), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n802), .B(KEYINPUT100), .Z(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(new_n626), .ZN(new_n846));
  OAI21_X1  g421(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n847));
  INV_X1    g422(.A(G118), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n847), .B1(new_n848), .B2(G2105), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n487), .A2(G130), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT99), .ZN(new_n851));
  AOI211_X1 g426(.A(new_n849), .B(new_n851), .C1(G142), .C2(new_n484), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n846), .B(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n841), .B1(new_n844), .B2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n853), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n843), .A2(new_n735), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n843), .A2(new_n735), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(G37), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n853), .A2(KEYINPUT101), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n844), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n856), .A2(KEYINPUT101), .A3(new_n853), .A4(new_n857), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(new_n841), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n859), .A2(new_n860), .A3(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g441(.A1(new_n609), .A2(G299), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n604), .A2(new_n570), .A3(new_n573), .A4(new_n608), .ZN(new_n868));
  AND3_X1   g443(.A1(new_n867), .A2(KEYINPUT41), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(KEYINPUT41), .B1(new_n867), .B2(new_n868), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n620), .B(new_n829), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n867), .A2(new_n868), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n874), .B1(new_n876), .B2(new_n873), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n877), .A2(KEYINPUT42), .ZN(new_n878));
  XNOR2_X1  g453(.A(G303), .B(G305), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n786), .B(G290), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n879), .B(new_n880), .Z(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n877), .A2(KEYINPUT42), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n878), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n882), .B1(new_n878), .B2(new_n883), .ZN(new_n885));
  OAI21_X1  g460(.A(G868), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n826), .A2(new_n613), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(G295));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n887), .ZN(G331));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n890));
  NAND2_X1  g465(.A1(G286), .A2(G301), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(G286), .A2(G301), .ZN(new_n893));
  OAI22_X1  g468(.A1(new_n892), .A2(new_n893), .B1(new_n827), .B2(new_n828), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n826), .A2(new_n557), .ZN(new_n895));
  NAND2_X1  g470(.A1(G171), .A2(G168), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n826), .A2(new_n557), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n895), .A2(new_n896), .A3(new_n897), .A4(new_n891), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT103), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n894), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n892), .A2(new_n893), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n901), .A2(new_n829), .A3(KEYINPUT103), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n898), .A2(KEYINPUT102), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT102), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n901), .A2(new_n829), .A3(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n904), .A2(new_n906), .A3(new_n894), .ZN(new_n907));
  OAI22_X1  g482(.A1(new_n872), .A2(new_n903), .B1(new_n907), .B2(new_n875), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n882), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n875), .B1(new_n900), .B2(new_n902), .ZN(new_n910));
  AOI22_X1  g485(.A1(new_n910), .A2(KEYINPUT104), .B1(new_n871), .B2(new_n907), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n903), .A2(new_n876), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT104), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n911), .A2(new_n914), .A3(new_n881), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n909), .A2(new_n860), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n890), .B1(new_n916), .B2(KEYINPUT43), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n860), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n881), .B1(new_n911), .B2(new_n914), .ZN(new_n919));
  OR2_X1    g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n917), .B1(new_n920), .B2(KEYINPUT43), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT105), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT43), .B1(new_n918), .B2(new_n919), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n909), .A2(new_n915), .A3(new_n924), .A4(new_n860), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n922), .B1(new_n926), .B2(new_n890), .ZN(new_n927));
  AOI211_X1 g502(.A(KEYINPUT105), .B(KEYINPUT44), .C1(new_n923), .C2(new_n925), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n921), .B1(new_n927), .B2(new_n928), .ZN(G397));
  INV_X1    g504(.A(KEYINPUT47), .ZN(new_n930));
  XNOR2_X1  g505(.A(KEYINPUT106), .B(G1384), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n500), .A2(new_n504), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n508), .B1(new_n624), .B2(new_n496), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n932), .B1(new_n498), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n497), .A2(KEYINPUT70), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n935), .A2(KEYINPUT4), .A3(new_n510), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n931), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  OAI211_X1 g512(.A(G40), .B(new_n472), .C1(new_n480), .C2(new_n481), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n937), .A2(KEYINPUT45), .A3(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n725), .A2(G2067), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n727), .B1(new_n720), .B2(new_n724), .ZN(new_n943));
  OR3_X1    g518(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n942), .B1(new_n941), .B2(new_n943), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n940), .B1(new_n946), .B2(new_n699), .ZN(new_n947));
  INV_X1    g522(.A(G1996), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n939), .A2(new_n948), .ZN(new_n949));
  XOR2_X1   g524(.A(new_n949), .B(KEYINPUT46), .Z(new_n950));
  OAI21_X1  g525(.A(new_n930), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NOR3_X1   g527(.A1(new_n947), .A2(new_n950), .A3(new_n930), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT125), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n953), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT125), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n955), .A2(new_n956), .A3(new_n951), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n946), .A2(new_n948), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n947), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n699), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n949), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n802), .A2(new_n804), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n960), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n939), .B1(new_n965), .B2(new_n941), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n802), .B(new_n804), .ZN(new_n967));
  XOR2_X1   g542(.A(new_n967), .B(KEYINPUT108), .Z(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n939), .ZN(new_n969));
  NOR2_X1   g544(.A1(G290), .A2(G1986), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n939), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n971), .B(KEYINPUT48), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n960), .A2(new_n963), .A3(new_n969), .A4(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n958), .A2(KEYINPUT126), .A3(new_n966), .A4(new_n973), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n966), .A2(new_n954), .A3(new_n973), .A4(new_n957), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT126), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  XOR2_X1   g553(.A(KEYINPUT111), .B(G8), .Z(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G1384), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n935), .A2(KEYINPUT4), .A3(new_n510), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n499), .A2(new_n504), .A3(new_n500), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT50), .ZN(new_n985));
  INV_X1    g560(.A(new_n938), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT50), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n512), .A2(new_n987), .A3(new_n981), .ZN(new_n988));
  AND4_X1   g563(.A1(new_n708), .A2(new_n985), .A3(new_n986), .A4(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n938), .B1(new_n984), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(G1384), .B1(new_n934), .B2(new_n936), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(KEYINPUT45), .ZN(new_n993));
  AOI21_X1  g568(.A(G1966), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n980), .B1(new_n989), .B2(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(G168), .A2(new_n979), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n996), .A2(KEYINPUT51), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G8), .ZN(new_n999));
  INV_X1    g574(.A(G1966), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n986), .B1(new_n992), .B2(KEYINPUT45), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n984), .A2(new_n990), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1000), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n938), .B1(new_n984), .B2(KEYINPUT50), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1004), .A2(new_n708), .A3(new_n988), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n999), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT51), .B1(new_n1006), .B2(new_n996), .ZN(new_n1007));
  OAI211_X1 g582(.A(G286), .B(new_n980), .C1(new_n989), .C2(new_n994), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n998), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT62), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(G1961), .B1(new_n1004), .B2(new_n988), .ZN(new_n1013));
  INV_X1    g588(.A(G2078), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT109), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1015), .B1(new_n937), .B2(KEYINPUT45), .ZN(new_n1016));
  INV_X1    g591(.A(new_n931), .ZN(new_n1017));
  AND4_X1   g592(.A1(new_n1015), .A2(new_n512), .A3(KEYINPUT45), .A4(new_n1017), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1014), .B(new_n991), .C1(new_n1016), .C2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1013), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n991), .A2(KEYINPUT53), .A3(new_n1014), .A4(new_n993), .ZN(new_n1022));
  AOI21_X1  g597(.A(G301), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g598(.A(KEYINPUT110), .B(KEYINPUT55), .ZN(new_n1024));
  AND3_X1   g599(.A1(G303), .A2(G8), .A3(new_n1024), .ZN(new_n1025));
  AND2_X1   g600(.A1(KEYINPUT110), .A2(KEYINPUT55), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1026), .B1(G303), .B2(G8), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n991), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1029));
  AOI211_X1 g604(.A(KEYINPUT50), .B(G1384), .C1(new_n934), .C2(new_n936), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n987), .B1(new_n512), .B2(new_n981), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n1030), .A2(new_n1031), .A3(new_n938), .ZN(new_n1032));
  AOI22_X1  g607(.A1(new_n1029), .A2(new_n783), .B1(new_n1032), .B2(new_n767), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1028), .B1(new_n1033), .B2(new_n979), .ZN(new_n1034));
  NAND3_X1  g609(.A1(G303), .A2(G8), .A3(new_n1024), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n999), .B1(new_n521), .B2(new_n530), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1035), .B1(new_n1036), .B2(new_n1026), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n512), .A2(new_n1017), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT109), .B1(new_n1038), .B2(new_n990), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n937), .A2(new_n1015), .A3(KEYINPUT45), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(G1971), .B1(new_n1041), .B2(new_n991), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n985), .A2(new_n986), .A3(new_n988), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1043), .A2(G2090), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1037), .B(G8), .C1(new_n1042), .C2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n580), .A2(G1976), .A3(new_n581), .A4(new_n582), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1046), .B(new_n980), .C1(new_n984), .C2(new_n938), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(KEYINPUT52), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1049), .B1(new_n786), .B2(G1976), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1048), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n591), .A2(new_n586), .ZN(new_n1052));
  INV_X1    g627(.A(G1981), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1052), .A2(new_n1053), .A3(new_n585), .A4(new_n593), .ZN(new_n1054));
  NAND2_X1  g629(.A1(G305), .A2(G1981), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1054), .A2(new_n1055), .A3(KEYINPUT49), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT112), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1054), .A2(new_n1055), .A3(KEYINPUT112), .A4(KEYINPUT49), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT49), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n986), .A2(new_n992), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n980), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1051), .B1(new_n1060), .B2(new_n1064), .ZN(new_n1065));
  AND4_X1   g640(.A1(new_n1023), .A2(new_n1034), .A3(new_n1045), .A4(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT123), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1012), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1008), .B(KEYINPUT51), .C1(new_n996), .C2(new_n1006), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT62), .B1(new_n1069), .B2(new_n998), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1023), .A2(new_n1034), .A3(new_n1045), .A4(new_n1065), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT123), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT124), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT124), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1069), .A2(new_n1074), .A3(KEYINPUT62), .A4(new_n998), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1068), .A2(new_n1072), .A3(new_n1073), .A4(new_n1075), .ZN(new_n1076));
  XOR2_X1   g651(.A(new_n1054), .B(KEYINPUT113), .Z(new_n1077));
  NAND2_X1  g652(.A1(new_n1060), .A2(new_n1064), .ZN(new_n1078));
  NOR2_X1   g653(.A1(G288), .A2(G1976), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1077), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1065), .ZN(new_n1081));
  OAI22_X1  g656(.A1(new_n1080), .A2(new_n1063), .B1(new_n1081), .B2(new_n1045), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n1065), .A2(new_n1045), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n995), .A2(G286), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1028), .B1(new_n1033), .B2(new_n999), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1083), .A2(KEYINPUT63), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1034), .A2(new_n1065), .A3(new_n1045), .A4(new_n1084), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT63), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1082), .B1(new_n1086), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1076), .A2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT56), .B(G2072), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1041), .A2(new_n991), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT114), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1001), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT114), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1095), .A2(new_n1096), .A3(new_n1092), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(G1956), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1043), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g676(.A(G299), .B(KEYINPUT57), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1102), .B(KEYINPUT118), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(G1348), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1043), .A2(new_n1105), .ZN(new_n1106));
  OR4_X1    g681(.A1(KEYINPUT116), .A2(new_n984), .A3(G2067), .A4(new_n938), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n986), .A2(new_n992), .A3(new_n727), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT116), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1106), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT117), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n1043), .A2(new_n1105), .B1(KEYINPUT116), .B2(new_n1108), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT117), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1112), .A2(new_n1113), .A3(new_n1107), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1104), .B1(new_n609), .B2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1032), .A2(G1956), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1117), .A2(new_n1102), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1093), .A2(KEYINPUT114), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1096), .B1(new_n1095), .B2(new_n1092), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1118), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(KEYINPUT115), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT115), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1098), .A2(new_n1123), .A3(new_n1118), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1116), .A2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1115), .A2(KEYINPUT60), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT60), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1128), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT120), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n610), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1112), .A2(new_n1113), .A3(new_n1107), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1113), .B1(new_n1112), .B2(new_n1107), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT60), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1134), .A2(KEYINPUT120), .A3(new_n609), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1131), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1127), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1139), .B1(new_n1098), .B2(new_n1118), .ZN(new_n1140));
  XNOR2_X1  g715(.A(KEYINPUT119), .B(G1996), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1041), .A2(new_n991), .A3(new_n1141), .ZN(new_n1142));
  XOR2_X1   g717(.A(KEYINPUT58), .B(G1341), .Z(new_n1143));
  NAND2_X1  g718(.A1(new_n1062), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n557), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT59), .ZN(new_n1146));
  OR2_X1    g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1104), .A2(new_n1140), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1122), .A2(new_n1124), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1149), .B1(new_n1150), .B2(KEYINPUT61), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1126), .B1(new_n1138), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT54), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n938), .A2(new_n1020), .A3(G2078), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1041), .B(new_n1154), .C1(KEYINPUT45), .C2(new_n937), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(KEYINPUT121), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(new_n1021), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1153), .B1(new_n1157), .B2(G171), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1021), .A2(G301), .A3(new_n1022), .ZN(new_n1159));
  XOR2_X1   g734(.A(new_n1159), .B(KEYINPUT122), .Z(new_n1160));
  NAND2_X1  g735(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n1156), .A2(G301), .A3(new_n1021), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1153), .B1(new_n1162), .B2(new_n1023), .ZN(new_n1163));
  AND4_X1   g738(.A1(new_n1069), .A2(new_n1083), .A3(new_n998), .A4(new_n1034), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1161), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1091), .B1(new_n1152), .B2(new_n1165), .ZN(new_n1166));
  AND2_X1   g741(.A1(G290), .A2(G1986), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n939), .B1(new_n1167), .B2(new_n970), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n960), .A2(new_n1168), .A3(new_n963), .A4(new_n969), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n978), .B1(new_n1166), .B2(new_n1169), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g745(.A(G401), .ZN(new_n1172));
  INV_X1    g746(.A(KEYINPUT127), .ZN(new_n1173));
  NOR2_X1   g747(.A1(G227), .A2(new_n461), .ZN(new_n1174));
  NAND3_X1  g748(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  INV_X1    g749(.A(new_n1174), .ZN(new_n1176));
  OAI21_X1  g750(.A(KEYINPUT127), .B1(G401), .B2(new_n1176), .ZN(new_n1177));
  AND4_X1   g751(.A1(new_n689), .A2(new_n865), .A3(new_n1175), .A4(new_n1177), .ZN(new_n1178));
  AND2_X1   g752(.A1(new_n1178), .A2(new_n926), .ZN(G308));
  NAND2_X1  g753(.A1(new_n1178), .A2(new_n926), .ZN(G225));
endmodule


