//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 0 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979;
  INV_X1    g000(.A(G43gat), .ZN(new_n202));
  INV_X1    g001(.A(G50gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G43gat), .A2(G50gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n206), .A2(KEYINPUT15), .ZN(new_n207));
  NAND2_X1  g006(.A1(G29gat), .A2(G36gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT83), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n206), .A2(KEYINPUT81), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT81), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n204), .A2(new_n213), .A3(new_n205), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(KEYINPUT15), .A3(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G29gat), .ZN(new_n216));
  INV_X1    g015(.A(G36gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(new_n217), .A3(KEYINPUT14), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT14), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(G29gat), .B2(G36gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  OR2_X1    g020(.A1(new_n221), .A2(KEYINPUT82), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(KEYINPUT82), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n211), .A2(new_n215), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n218), .A2(new_n220), .A3(new_n208), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n212), .A2(KEYINPUT15), .A3(new_n225), .A4(new_n214), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT17), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G15gat), .B(G22gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT16), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n230), .B1(new_n231), .B2(G1gat), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(G1gat), .B2(new_n230), .ZN(new_n233));
  INV_X1    g032(.A(G8gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n224), .A2(KEYINPUT17), .A3(new_n226), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n229), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n235), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(new_n227), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G229gat), .A2(G233gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n240), .A2(KEYINPUT18), .A3(new_n241), .ZN(new_n242));
  XOR2_X1   g041(.A(new_n235), .B(new_n227), .Z(new_n243));
  XOR2_X1   g042(.A(new_n241), .B(KEYINPUT13), .Z(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n237), .A2(new_n241), .A3(new_n239), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT18), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n242), .A2(new_n245), .A3(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G113gat), .B(G141gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(G197gat), .ZN(new_n251));
  XOR2_X1   g050(.A(KEYINPUT11), .B(G169gat), .Z(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(KEYINPUT12), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n249), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n242), .A2(new_n254), .A3(new_n245), .A4(new_n248), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(G228gat), .A2(G233gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(G211gat), .B(G218gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(G197gat), .B(G204gat), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT22), .ZN(new_n263));
  INV_X1    g062(.A(G211gat), .ZN(new_n264));
  INV_X1    g063(.A(G218gat), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n261), .A2(new_n262), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n261), .B1(new_n266), .B2(new_n262), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  XOR2_X1   g069(.A(G155gat), .B(G162gat), .Z(new_n271));
  OR2_X1    g070(.A1(G141gat), .A2(G148gat), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT2), .ZN(new_n273));
  NAND2_X1  g072(.A1(G141gat), .A2(G148gat), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(KEYINPUT72), .B(KEYINPUT3), .ZN(new_n277));
  INV_X1    g076(.A(G162gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT71), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(G162gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n273), .B1(new_n282), .B2(G155gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(G155gat), .B(G162gat), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n284), .A2(new_n272), .A3(new_n274), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n276), .B(new_n277), .C1(new_n283), .C2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT73), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AND2_X1   g087(.A1(new_n272), .A2(new_n274), .ZN(new_n289));
  INV_X1    g088(.A(G155gat), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n290), .B1(new_n279), .B2(new_n281), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n289), .B(new_n284), .C1(new_n291), .C2(new_n273), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n292), .A2(KEYINPUT73), .A3(new_n276), .A4(new_n277), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n288), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT29), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n270), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n284), .A2(new_n272), .A3(new_n274), .ZN(new_n297));
  XNOR2_X1  g096(.A(KEYINPUT71), .B(G162gat), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT2), .B1(new_n298), .B2(new_n290), .ZN(new_n299));
  AOI22_X1  g098(.A1(new_n297), .A2(new_n299), .B1(new_n271), .B2(new_n275), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n270), .A2(new_n295), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n300), .B1(new_n301), .B2(new_n277), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n260), .B1(new_n296), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G22gat), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT3), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n305), .B1(new_n269), .B2(KEYINPUT29), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n276), .B1(new_n283), .B2(new_n285), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n260), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT29), .B1(new_n288), .B2(new_n293), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n308), .B1(new_n309), .B2(new_n270), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n303), .A2(new_n304), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT77), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT77), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n303), .A2(new_n313), .A3(new_n304), .A4(new_n310), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n303), .A2(new_n310), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G22gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n312), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G78gat), .B(G106gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n318), .B(new_n203), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n319), .B(KEYINPUT75), .ZN(new_n320));
  XOR2_X1   g119(.A(KEYINPUT74), .B(KEYINPUT31), .Z(new_n321));
  XOR2_X1   g120(.A(new_n320), .B(new_n321), .Z(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n317), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT78), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT76), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n303), .A2(KEYINPUT76), .A3(new_n304), .A4(new_n310), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n327), .A2(new_n316), .A3(new_n322), .A4(new_n328), .ZN(new_n329));
  AND3_X1   g128(.A1(new_n324), .A2(new_n325), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n325), .B1(new_n324), .B2(new_n329), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(G169gat), .ZN(new_n333));
  INV_X1    g132(.A(G176gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n333), .A2(new_n334), .A3(KEYINPUT23), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT23), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n336), .B1(G169gat), .B2(G176gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(G169gat), .A2(G176gat), .ZN(new_n338));
  AND3_X1   g137(.A1(new_n335), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(KEYINPUT65), .B(G183gat), .ZN(new_n340));
  INV_X1    g139(.A(G190gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(G183gat), .A2(G190gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT24), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT24), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n344), .A2(G183gat), .A3(G190gat), .ZN(new_n345));
  AOI22_X1  g144(.A1(new_n340), .A2(new_n341), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT66), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n339), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(G183gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT65), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT65), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(G183gat), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n350), .A2(new_n352), .A3(new_n341), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n343), .A2(new_n345), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n355), .A2(KEYINPUT66), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT25), .B1(new_n348), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n333), .A2(new_n334), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT26), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n342), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n360), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT27), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(new_n349), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n364), .B1(new_n340), .B2(new_n363), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT28), .B1(new_n365), .B2(new_n341), .ZN(new_n366));
  XOR2_X1   g165(.A(KEYINPUT27), .B(G183gat), .Z(new_n367));
  INV_X1    g166(.A(KEYINPUT28), .ZN(new_n368));
  NOR3_X1   g167(.A1(new_n367), .A2(new_n368), .A3(G190gat), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n362), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n354), .B1(G183gat), .B2(G190gat), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT25), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n371), .A2(new_n372), .A3(new_n339), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n370), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(G120gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(G113gat), .ZN(new_n376));
  INV_X1    g175(.A(G113gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(G120gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT1), .ZN(new_n380));
  INV_X1    g179(.A(G134gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(G127gat), .ZN(new_n382));
  INV_X1    g181(.A(G127gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(G134gat), .ZN(new_n384));
  AOI22_X1  g183(.A1(new_n379), .A2(new_n380), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT67), .ZN(new_n386));
  AND3_X1   g185(.A1(new_n376), .A2(new_n378), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n375), .A2(KEYINPUT67), .A3(G113gat), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n388), .A2(new_n382), .A3(new_n384), .A4(new_n380), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT68), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  AND3_X1   g189(.A1(new_n382), .A2(new_n384), .A3(new_n380), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT68), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n376), .A2(new_n378), .A3(new_n386), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n391), .A2(new_n392), .A3(new_n393), .A4(new_n388), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n385), .B1(new_n390), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n374), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n373), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n346), .A2(new_n347), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n355), .A2(KEYINPUT66), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(new_n399), .A3(new_n339), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n397), .B1(new_n400), .B2(KEYINPUT25), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n390), .A2(new_n394), .ZN(new_n402));
  INV_X1    g201(.A(new_n385), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n401), .A2(new_n404), .A3(new_n370), .ZN(new_n405));
  NAND2_X1  g204(.A1(G227gat), .A2(G233gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n406), .B(KEYINPUT64), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n396), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT32), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT33), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  XOR2_X1   g210(.A(G15gat), .B(G43gat), .Z(new_n412));
  XNOR2_X1  g211(.A(G71gat), .B(G99gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n409), .A2(new_n411), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n414), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n408), .B(KEYINPUT32), .C1(new_n410), .C2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT69), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT69), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n415), .A2(new_n420), .A3(new_n417), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n396), .A2(new_n405), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(new_n406), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT34), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n407), .A2(KEYINPUT34), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n419), .A2(new_n421), .A3(new_n428), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n427), .A2(new_n420), .A3(new_n415), .A4(new_n417), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(G225gat), .A2(G233gat), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n402), .A2(new_n300), .A3(new_n403), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n395), .A2(new_n300), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT5), .ZN(new_n437));
  AOI22_X1  g236(.A1(new_n402), .A2(new_n403), .B1(new_n307), .B2(KEYINPUT3), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n294), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT4), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n440), .B1(new_n404), .B2(new_n307), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n395), .A2(KEYINPUT4), .A3(new_n300), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n439), .A2(new_n441), .A3(new_n432), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n437), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n442), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT4), .B1(new_n395), .B2(new_n300), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n447), .A2(KEYINPUT5), .A3(new_n432), .A4(new_n439), .ZN(new_n448));
  XNOR2_X1  g247(.A(G1gat), .B(G29gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n449), .B(KEYINPUT0), .ZN(new_n450));
  XNOR2_X1  g249(.A(G57gat), .B(G85gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  AND4_X1   g251(.A1(KEYINPUT6), .A2(new_n444), .A3(new_n448), .A4(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n444), .A2(new_n448), .ZN(new_n454));
  INV_X1    g253(.A(new_n452), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT6), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n452), .B(KEYINPUT79), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n444), .A2(new_n448), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n453), .B1(new_n456), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(G226gat), .A2(G233gat), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n462), .B1(new_n374), .B2(new_n295), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n461), .B1(new_n401), .B2(new_n370), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n269), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n374), .A2(new_n462), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT29), .B1(new_n401), .B2(new_n370), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n466), .B(new_n270), .C1(new_n467), .C2(new_n462), .ZN(new_n468));
  XOR2_X1   g267(.A(G8gat), .B(G36gat), .Z(new_n469));
  XNOR2_X1  g268(.A(new_n469), .B(KEYINPUT70), .ZN(new_n470));
  XNOR2_X1  g269(.A(G64gat), .B(G92gat), .ZN(new_n471));
  XOR2_X1   g270(.A(new_n470), .B(new_n471), .Z(new_n472));
  NAND3_X1  g271(.A1(new_n465), .A2(new_n468), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT30), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n465), .A2(new_n468), .A3(KEYINPUT30), .A4(new_n472), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n465), .A2(new_n468), .ZN(new_n477));
  INV_X1    g276(.A(new_n472), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n475), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  NOR3_X1   g279(.A1(new_n460), .A2(new_n480), .A3(KEYINPUT35), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n332), .A2(KEYINPUT80), .A3(new_n431), .A4(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n304), .B1(new_n303), .B2(new_n310), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n483), .B1(KEYINPUT77), .B2(new_n311), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n322), .B1(new_n484), .B2(new_n314), .ZN(new_n485));
  INV_X1    g284(.A(new_n329), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT78), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n324), .A2(new_n325), .A3(new_n329), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n431), .A2(new_n481), .A3(new_n487), .A4(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT80), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n444), .A2(new_n448), .A3(new_n452), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n453), .B1(new_n456), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n493), .A2(new_n480), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n431), .A2(new_n487), .A3(new_n488), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT35), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n482), .A2(new_n491), .A3(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n459), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n447), .A2(new_n439), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n433), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n457), .B1(new_n500), .B2(KEYINPUT39), .ZN(new_n501));
  OR2_X1    g300(.A1(new_n434), .A2(new_n435), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT39), .B1(new_n502), .B2(new_n433), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n503), .B1(new_n433), .B2(new_n499), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n498), .B1(new_n505), .B2(KEYINPUT40), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n506), .B(new_n480), .C1(KEYINPUT40), .C2(new_n505), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n477), .A2(KEYINPUT37), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT37), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n465), .A2(new_n468), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n508), .A2(new_n478), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT38), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT38), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n508), .A2(new_n513), .A3(new_n478), .A4(new_n510), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n512), .A2(new_n460), .A3(new_n473), .A4(new_n514), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n507), .A2(new_n515), .A3(new_n487), .A4(new_n488), .ZN(new_n516));
  INV_X1    g315(.A(new_n431), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT36), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT36), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n431), .A2(new_n519), .ZN(new_n520));
  OAI22_X1  g319(.A1(new_n330), .A2(new_n331), .B1(new_n493), .B2(new_n480), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n516), .A2(new_n518), .A3(new_n520), .A4(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n259), .B1(new_n497), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT92), .ZN(new_n524));
  XOR2_X1   g323(.A(G134gat), .B(G162gat), .Z(new_n525));
  AND2_X1   g324(.A1(G232gat), .A2(G233gat), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n526), .A2(KEYINPUT41), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n525), .B(new_n527), .ZN(new_n528));
  XOR2_X1   g327(.A(new_n528), .B(KEYINPUT91), .Z(new_n529));
  INV_X1    g328(.A(G85gat), .ZN(new_n530));
  INV_X1    g329(.A(G92gat), .ZN(new_n531));
  OAI211_X1 g330(.A(KEYINPUT87), .B(KEYINPUT7), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(KEYINPUT87), .A2(KEYINPUT7), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n533), .A2(G85gat), .A3(G92gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(G99gat), .A2(G106gat), .ZN(new_n536));
  AOI22_X1  g335(.A1(KEYINPUT8), .A2(new_n536), .B1(new_n530), .B2(new_n531), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  OR2_X1    g337(.A1(G99gat), .A2(G106gat), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n538), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n536), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n535), .A2(new_n541), .A3(new_n537), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n229), .A2(KEYINPUT88), .A3(new_n236), .A4(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n526), .A2(KEYINPUT41), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n543), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n546), .B1(new_n227), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT89), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n543), .B1(new_n226), .B2(new_n224), .ZN(new_n551));
  NOR3_X1   g350(.A1(new_n551), .A2(KEYINPUT89), .A3(new_n546), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n544), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n229), .A2(new_n236), .A3(new_n543), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT88), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(KEYINPUT90), .B1(new_n553), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G190gat), .B(G218gat), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n548), .A2(new_n549), .ZN(new_n561));
  OAI21_X1  g360(.A(KEYINPUT89), .B1(new_n551), .B2(new_n546), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT90), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n563), .A2(new_n556), .A3(new_n564), .A4(new_n544), .ZN(new_n565));
  AND3_X1   g364(.A1(new_n558), .A2(new_n560), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n560), .B1(new_n558), .B2(new_n565), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n529), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n558), .A2(new_n565), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(new_n559), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n528), .A2(KEYINPUT91), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n558), .A2(new_n560), .A3(new_n565), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(new_n290), .ZN(new_n577));
  XNOR2_X1  g376(.A(G183gat), .B(G211gat), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n577), .B(new_n578), .Z(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(G57gat), .ZN(new_n581));
  OAI21_X1  g380(.A(KEYINPUT85), .B1(new_n581), .B2(G64gat), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT85), .ZN(new_n583));
  INV_X1    g382(.A(G64gat), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n583), .A2(new_n584), .A3(G57gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n581), .A2(G64gat), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n582), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(G71gat), .A2(G78gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT9), .ZN(new_n589));
  NAND2_X1  g388(.A1(G71gat), .A2(G78gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT86), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n587), .A2(new_n591), .A3(KEYINPUT86), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n588), .B1(KEYINPUT84), .B2(new_n590), .ZN(new_n597));
  XNOR2_X1  g396(.A(G57gat), .B(G64gat), .ZN(new_n598));
  NOR2_X1   g397(.A1(KEYINPUT84), .A2(KEYINPUT9), .ZN(new_n599));
  OAI221_X1 g398(.A(new_n597), .B1(KEYINPUT84), .B2(new_n590), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT21), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G231gat), .A2(G233gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(G127gat), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n235), .B1(new_n602), .B2(new_n601), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n606), .A2(new_n607), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n580), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n606), .A2(new_n607), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n612), .A2(new_n608), .A3(new_n579), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n524), .B1(new_n575), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n611), .A2(new_n613), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n574), .A2(new_n616), .A3(KEYINPUT92), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G120gat), .B(G148gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(G176gat), .B(G204gat), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n619), .B(new_n620), .Z(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(G230gat), .A2(G233gat), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n596), .A2(new_n600), .A3(new_n542), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT93), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n538), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n535), .A2(KEYINPUT93), .A3(new_n537), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT94), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n541), .B(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n627), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(KEYINPUT95), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT95), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n627), .A2(new_n630), .A3(new_n633), .A4(new_n628), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n625), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n601), .A2(new_n543), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n624), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(KEYINPUT97), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT97), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n640), .B(new_n624), .C1(new_n635), .C2(new_n637), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n623), .B(KEYINPUT98), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT10), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n632), .A2(new_n634), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n644), .B(new_n636), .C1(new_n645), .C2(new_n625), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n543), .A2(new_n644), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n647), .A2(KEYINPUT96), .A3(new_n596), .A4(new_n600), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT96), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n540), .A2(KEYINPUT10), .A3(new_n542), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n649), .B1(new_n601), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n643), .B1(new_n646), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n622), .B1(new_n642), .B2(new_n653), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n635), .A2(new_n637), .A3(KEYINPUT10), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n648), .A2(new_n651), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n623), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n657), .A2(new_n641), .A3(new_n639), .A4(new_n621), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT99), .ZN(new_n659));
  AND3_X1   g458(.A1(new_n654), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n659), .B1(new_n654), .B2(new_n658), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n618), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n523), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n493), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g467(.A(new_n234), .B1(new_n666), .B2(new_n480), .ZN(new_n669));
  INV_X1    g468(.A(new_n480), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT16), .B(G8gat), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n665), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(KEYINPUT42), .B1(new_n669), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n673), .B1(KEYINPUT42), .B2(new_n672), .ZN(G1325gat));
  NAND2_X1  g473(.A1(new_n518), .A2(new_n520), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT100), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n518), .A2(KEYINPUT100), .A3(new_n520), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(G15gat), .B1(new_n665), .B2(new_n680), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n517), .A2(G15gat), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n681), .B1(new_n665), .B2(new_n682), .ZN(G1326gat));
  NOR2_X1   g482(.A1(new_n665), .A2(new_n332), .ZN(new_n684));
  XOR2_X1   g483(.A(KEYINPUT43), .B(G22gat), .Z(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1327gat));
  NAND2_X1  g485(.A1(new_n497), .A2(new_n522), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n575), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(KEYINPUT44), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n574), .A2(KEYINPUT103), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT103), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n568), .A2(new_n573), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n696), .B1(new_n522), .B2(new_n497), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n689), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n614), .A2(new_n662), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(new_n259), .ZN(new_n701));
  XOR2_X1   g500(.A(new_n701), .B(KEYINPUT102), .Z(new_n702));
  AND2_X1   g501(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n493), .ZN(new_n705));
  OAI21_X1  g504(.A(G29gat), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n700), .A2(new_n574), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n707), .B(KEYINPUT101), .Z(new_n708));
  AND2_X1   g507(.A1(new_n708), .A2(new_n523), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n709), .A2(new_n216), .A3(new_n493), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT45), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n706), .A2(new_n711), .ZN(G1328gat));
  NAND3_X1  g511(.A1(new_n709), .A2(new_n217), .A3(new_n480), .ZN(new_n713));
  XOR2_X1   g512(.A(new_n713), .B(KEYINPUT46), .Z(new_n714));
  OAI21_X1  g513(.A(G36gat), .B1(new_n704), .B2(new_n670), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(G1329gat));
  INV_X1    g515(.A(new_n675), .ZN(new_n717));
  OAI21_X1  g516(.A(G43gat), .B1(new_n704), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n517), .A2(G43gat), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n709), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n718), .A2(KEYINPUT47), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n202), .B1(new_n703), .B2(new_n679), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n722), .B1(new_n709), .B2(new_n719), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n721), .B1(new_n723), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g523(.A1(new_n487), .A2(new_n488), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n709), .A2(new_n203), .A3(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT106), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n726), .A2(new_n727), .ZN(new_n729));
  OAI21_X1  g528(.A(KEYINPUT48), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n703), .A2(new_n725), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT48), .ZN(new_n732));
  AOI22_X1  g531(.A1(new_n731), .A2(G50gat), .B1(KEYINPUT104), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n731), .A2(KEYINPUT104), .A3(G50gat), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT105), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n726), .B(new_n736), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n734), .B1(new_n738), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g538(.A1(new_n618), .A2(new_n258), .A3(new_n662), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n687), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n741), .A2(new_n705), .ZN(new_n742));
  XOR2_X1   g541(.A(KEYINPUT107), .B(G57gat), .Z(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(G1332gat));
  NOR2_X1   g543(.A1(new_n741), .A2(new_n670), .ZN(new_n745));
  NOR2_X1   g544(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n746));
  AND2_X1   g545(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(new_n745), .B2(new_n746), .ZN(G1333gat));
  INV_X1    g548(.A(new_n741), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n750), .A2(G71gat), .A3(new_n679), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n741), .A2(new_n517), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n752), .A2(KEYINPUT108), .ZN(new_n753));
  INV_X1    g552(.A(G71gat), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n752), .B2(KEYINPUT108), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n751), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g556(.A1(new_n750), .A2(new_n725), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g558(.A1(new_n616), .A2(new_n258), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n761), .A2(new_n662), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n763), .B1(new_n689), .B2(new_n698), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(G85gat), .B1(new_n765), .B2(new_n705), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n687), .A2(new_n575), .A3(new_n760), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT51), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n574), .B1(new_n497), .B2(new_n522), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n770), .A2(KEYINPUT51), .A3(new_n760), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n663), .A2(new_n530), .A3(new_n493), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n766), .B1(new_n773), .B2(new_n774), .ZN(G1336gat));
  AOI21_X1  g574(.A(new_n531), .B1(new_n764), .B2(new_n480), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n776), .A2(KEYINPUT52), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n663), .A2(new_n531), .A3(new_n480), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n773), .A2(new_n778), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n779), .A2(KEYINPUT110), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n779), .A2(KEYINPUT110), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n777), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  XOR2_X1   g581(.A(new_n778), .B(KEYINPUT109), .Z(new_n783));
  NOR2_X1   g582(.A1(new_n773), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT52), .B1(new_n784), .B2(new_n776), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n782), .A2(new_n785), .ZN(G1337gat));
  OAI21_X1  g585(.A(G99gat), .B1(new_n765), .B2(new_n680), .ZN(new_n787));
  OR3_X1    g586(.A1(new_n517), .A2(G99gat), .A3(new_n662), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n787), .B1(new_n773), .B2(new_n788), .ZN(G1338gat));
  AOI21_X1  g588(.A(new_n695), .B1(new_n687), .B2(new_n575), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n725), .B(new_n762), .C1(new_n790), .C2(new_n697), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(G106gat), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n332), .A2(G106gat), .A3(new_n662), .ZN(new_n793));
  XOR2_X1   g592(.A(new_n793), .B(KEYINPUT111), .Z(new_n794));
  OAI21_X1  g593(.A(new_n792), .B1(new_n773), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT53), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT112), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n798));
  INV_X1    g597(.A(new_n771), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT51), .B1(new_n770), .B2(new_n760), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n793), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AND4_X1   g600(.A1(new_n797), .A2(new_n792), .A3(new_n798), .A4(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT53), .B1(new_n772), .B2(new_n793), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n797), .B1(new_n803), .B2(new_n792), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n796), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(KEYINPUT113), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT113), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n796), .B(new_n807), .C1(new_n802), .C2(new_n804), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(G1339gat));
  NAND4_X1  g608(.A1(new_n615), .A2(new_n259), .A3(new_n617), .A4(new_n662), .ZN(new_n810));
  AND3_X1   g609(.A1(new_n568), .A2(new_n573), .A3(new_n691), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n691), .B1(new_n568), .B2(new_n573), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n646), .A2(new_n643), .A3(new_n652), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n657), .A2(KEYINPUT54), .A3(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n653), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n814), .A2(new_n622), .A3(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n240), .A2(new_n241), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n243), .A2(new_n244), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n253), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n257), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n814), .A2(KEYINPUT55), .A3(new_n622), .A4(new_n816), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n819), .A2(new_n658), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n811), .A2(new_n812), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n823), .B1(new_n660), .B2(new_n661), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT114), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n819), .A2(new_n258), .A3(new_n658), .A4(new_n824), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT114), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n830), .B(new_n823), .C1(new_n660), .C2(new_n661), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n828), .A2(new_n829), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n826), .B1(new_n693), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n810), .B1(new_n833), .B2(new_n616), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n517), .A2(new_n725), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NOR4_X1   g636(.A1(new_n835), .A2(new_n705), .A3(new_n480), .A4(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(G113gat), .B1(new_n838), .B2(new_n258), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n705), .A2(new_n480), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n332), .A2(new_n431), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n835), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n259), .A2(new_n377), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n839), .B1(new_n842), .B2(new_n843), .ZN(G1340gat));
  AOI21_X1  g643(.A(G120gat), .B1(new_n838), .B2(new_n663), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n662), .A2(new_n375), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n845), .B1(new_n842), .B2(new_n846), .ZN(G1341gat));
  NAND3_X1  g646(.A1(new_n838), .A2(new_n383), .A3(new_n616), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n835), .A2(new_n614), .A3(new_n841), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n848), .B1(new_n383), .B2(new_n849), .ZN(G1342gat));
  NOR3_X1   g649(.A1(new_n835), .A2(new_n574), .A3(new_n841), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n851), .A2(new_n381), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n838), .A2(new_n381), .A3(new_n575), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(new_n853), .B2(KEYINPUT56), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n854), .B1(KEYINPUT56), .B2(new_n853), .ZN(G1343gat));
  NOR2_X1   g654(.A1(new_n835), .A2(new_n705), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n679), .A2(new_n332), .A3(new_n480), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n858), .A2(G141gat), .A3(new_n259), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n859), .A2(KEYINPUT58), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n717), .A2(new_n840), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(KEYINPUT57), .B1(new_n834), .B2(new_n725), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n725), .A2(KEYINPUT57), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n575), .B1(new_n829), .B2(new_n827), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n614), .B1(new_n826), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n864), .B1(new_n866), .B2(new_n810), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n862), .B1(new_n863), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(G141gat), .B1(new_n868), .B2(new_n259), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n860), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT115), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n832), .A2(new_n693), .ZN(new_n872));
  OR3_X1    g671(.A1(new_n811), .A2(new_n812), .A3(new_n825), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n616), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n810), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n725), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n867), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n871), .B1(new_n878), .B2(new_n861), .ZN(new_n879));
  OAI211_X1 g678(.A(KEYINPUT115), .B(new_n862), .C1(new_n863), .C2(new_n867), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n879), .A2(new_n880), .A3(new_n258), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n859), .B1(new_n881), .B2(G141gat), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT58), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n870), .B1(new_n882), .B2(new_n883), .ZN(G1344gat));
  AND3_X1   g683(.A1(new_n834), .A2(KEYINPUT57), .A3(new_n725), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n574), .A2(new_n825), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n614), .B1(new_n865), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(new_n810), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT57), .B1(new_n888), .B2(new_n725), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n890), .A2(new_n662), .A3(new_n861), .ZN(new_n891));
  INV_X1    g690(.A(G148gat), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT59), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n879), .A2(new_n880), .A3(new_n663), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n894), .A2(new_n895), .A3(G148gat), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n663), .A2(new_n892), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n897), .B1(new_n858), .B2(new_n898), .ZN(G1345gat));
  NAND3_X1  g698(.A1(new_n879), .A2(new_n880), .A3(new_n616), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(G155gat), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n857), .A2(new_n493), .A3(new_n834), .A4(new_n616), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT116), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n902), .A2(new_n903), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n290), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n901), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(KEYINPUT117), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT117), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n901), .A2(new_n909), .A3(new_n906), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(G1346gat));
  AND2_X1   g710(.A1(new_n879), .A2(new_n880), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n693), .A2(new_n298), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n856), .A2(new_n575), .A3(new_n857), .ZN(new_n914));
  AOI22_X1  g713(.A1(new_n912), .A2(new_n913), .B1(new_n298), .B2(new_n914), .ZN(G1347gat));
  NAND2_X1  g714(.A1(new_n836), .A2(new_n480), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT118), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n917), .A2(new_n493), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n918), .A2(new_n834), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n333), .A3(new_n258), .ZN(new_n920));
  XOR2_X1   g719(.A(new_n920), .B(KEYINPUT119), .Z(new_n921));
  NOR2_X1   g720(.A1(new_n670), .A2(new_n493), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n837), .A2(new_n923), .ZN(new_n924));
  AND3_X1   g723(.A1(new_n834), .A2(new_n258), .A3(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n921), .B1(new_n333), .B2(new_n925), .ZN(G1348gat));
  NAND4_X1  g725(.A1(new_n834), .A2(G176gat), .A3(new_n663), .A4(new_n924), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n918), .A2(new_n663), .A3(new_n834), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n928), .A2(KEYINPUT120), .A3(new_n334), .ZN(new_n929));
  AOI21_X1  g728(.A(KEYINPUT120), .B1(new_n928), .B2(new_n334), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n927), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT121), .ZN(G1349gat));
  INV_X1    g731(.A(new_n367), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n919), .A2(new_n933), .A3(new_n616), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n834), .A2(new_n616), .A3(new_n924), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n934), .B1(new_n340), .B2(new_n935), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n936), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g736(.A1(new_n919), .A2(new_n341), .A3(new_n694), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n834), .A2(new_n575), .A3(new_n924), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT61), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n939), .A2(new_n940), .A3(G190gat), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n940), .B1(new_n939), .B2(G190gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n938), .B1(new_n941), .B2(new_n942), .ZN(G1351gat));
  OR2_X1    g742(.A1(new_n885), .A2(new_n889), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n923), .B1(new_n677), .B2(new_n678), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(G197gat), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n946), .A2(new_n947), .A3(new_n259), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n945), .B(new_n725), .C1(new_n874), .C2(new_n875), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT122), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n834), .A2(KEYINPUT122), .A3(new_n725), .A4(new_n945), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n951), .A2(new_n952), .A3(new_n258), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n948), .B1(new_n947), .B2(new_n953), .ZN(G1352gat));
  OR3_X1    g753(.A1(new_n949), .A2(G204gat), .A3(new_n662), .ZN(new_n955));
  OR2_X1    g754(.A1(new_n955), .A2(KEYINPUT123), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(KEYINPUT123), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT62), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g759(.A(G204gat), .B1(new_n946), .B2(new_n662), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n956), .A2(KEYINPUT62), .A3(new_n957), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(G1353gat));
  NAND4_X1  g762(.A1(new_n951), .A2(new_n952), .A3(new_n264), .A4(new_n616), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n944), .A2(new_n616), .A3(new_n945), .ZN(new_n965));
  AND4_X1   g764(.A1(KEYINPUT124), .A2(new_n965), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n966));
  OAI21_X1  g765(.A(G211gat), .B1(KEYINPUT124), .B2(KEYINPUT63), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  AOI22_X1  g767(.A1(new_n965), .A2(new_n968), .B1(KEYINPUT124), .B2(KEYINPUT63), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n964), .B1(new_n966), .B2(new_n969), .ZN(G1354gat));
  NAND4_X1  g769(.A1(new_n944), .A2(G218gat), .A3(new_n575), .A4(new_n945), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n951), .A2(new_n952), .A3(new_n694), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT125), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n972), .A2(new_n973), .A3(new_n265), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n973), .B1(new_n972), .B2(new_n265), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n971), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT126), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI211_X1 g777(.A(new_n971), .B(KEYINPUT126), .C1(new_n974), .C2(new_n975), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(G1355gat));
endmodule


