//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 1 0 0 0 0 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n641, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n819, new_n820, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968;
  XOR2_X1   g000(.A(G15gat), .B(G22gat), .Z(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G15gat), .B(G22gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n205), .B1(new_n206), .B2(G1gat), .ZN(new_n207));
  INV_X1    g006(.A(G8gat), .ZN(new_n208));
  AND3_X1   g007(.A1(new_n204), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n208), .B1(new_n204), .B2(new_n207), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT86), .ZN(new_n212));
  INV_X1    g011(.A(G50gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n212), .B1(new_n213), .B2(G43gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(G43gat), .ZN(new_n215));
  INV_X1    g014(.A(G43gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n216), .A2(KEYINPUT86), .A3(G50gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n214), .A2(new_n215), .A3(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT15), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT15), .B1(new_n213), .B2(G43gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n216), .A2(G50gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G29gat), .ZN(new_n225));
  INV_X1    g024(.A(G36gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(new_n226), .A3(KEYINPUT14), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT14), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n228), .B1(G29gat), .B2(G36gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(G29gat), .A2(G36gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n227), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n220), .A2(new_n224), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT85), .ZN(new_n234));
  AND3_X1   g033(.A1(new_n231), .A2(new_n223), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n234), .B1(new_n231), .B2(new_n223), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n233), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n211), .A2(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n209), .A2(new_n210), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n231), .A2(new_n223), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT85), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n231), .A2(new_n223), .A3(new_n234), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n231), .A2(new_n223), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n241), .A2(new_n242), .B1(new_n220), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n239), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n238), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(G229gat), .A2(G233gat), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n247), .B(KEYINPUT13), .Z(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G113gat), .B(G141gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(G169gat), .B(G197gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(KEYINPUT12), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n233), .B(KEYINPUT17), .C1(new_n236), .C2(new_n235), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT87), .B(KEYINPUT17), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n257), .B(new_n239), .C1(new_n244), .C2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT88), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n258), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n237), .A2(new_n262), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n263), .A2(KEYINPUT88), .A3(new_n239), .A4(new_n257), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n238), .A2(new_n247), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT18), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n249), .B(new_n256), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n268), .A2(KEYINPUT89), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n266), .B1(new_n261), .B2(new_n264), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT89), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n271), .A2(new_n269), .A3(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT90), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n270), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT91), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n271), .A2(KEYINPUT90), .A3(new_n269), .A4(new_n274), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n269), .B1(new_n272), .B2(new_n273), .ZN(new_n281));
  AOI211_X1 g080(.A(KEYINPUT89), .B(new_n266), .C1(new_n261), .C2(new_n264), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n276), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n249), .ZN(new_n284));
  AOI211_X1 g083(.A(new_n255), .B(new_n284), .C1(new_n272), .C2(KEYINPUT18), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n283), .A2(new_n279), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT91), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n275), .B(new_n249), .C1(new_n269), .C2(new_n268), .ZN(new_n288));
  AOI22_X1  g087(.A1(new_n280), .A2(new_n287), .B1(new_n288), .B2(new_n255), .ZN(new_n289));
  NAND2_X1  g088(.A1(G226gat), .A2(G233gat), .ZN(new_n290));
  INV_X1    g089(.A(G169gat), .ZN(new_n291));
  INV_X1    g090(.A(G176gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n293), .B(KEYINPUT65), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT26), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297));
  INV_X1    g096(.A(new_n293), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n296), .B(new_n297), .C1(new_n295), .C2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT27), .B(G183gat), .ZN(new_n300));
  INV_X1    g099(.A(G190gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT28), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT67), .ZN(new_n304));
  AOI22_X1  g103(.A1(new_n302), .A2(new_n304), .B1(G183gat), .B2(G190gat), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n299), .B(new_n305), .C1(new_n302), .C2(new_n304), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n294), .A2(KEYINPUT23), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT24), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n308), .A2(G183gat), .A3(G190gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(G183gat), .B(G190gat), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n309), .B1(new_n310), .B2(new_n308), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT66), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT23), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n293), .A2(new_n313), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n314), .A2(KEYINPUT25), .ZN(new_n315));
  XOR2_X1   g114(.A(new_n297), .B(KEYINPUT64), .Z(new_n316));
  NAND4_X1  g115(.A1(new_n307), .A2(new_n312), .A3(new_n315), .A4(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n311), .A2(KEYINPUT66), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n298), .A2(KEYINPUT23), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n319), .A2(new_n314), .A3(new_n297), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n320), .A2(new_n311), .ZN(new_n321));
  OAI22_X1  g120(.A1(new_n317), .A2(new_n318), .B1(KEYINPUT25), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n290), .B1(new_n324), .B2(KEYINPUT29), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n323), .A2(G226gat), .A3(G233gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT22), .ZN(new_n328));
  INV_X1    g127(.A(G211gat), .ZN(new_n329));
  INV_X1    g128(.A(G218gat), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT72), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT72), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n333), .B(new_n328), .C1(new_n329), .C2(new_n330), .ZN(new_n334));
  XNOR2_X1  g133(.A(G197gat), .B(G204gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n332), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G211gat), .B(G218gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n336), .B(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n327), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n338), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n325), .A2(new_n340), .A3(new_n326), .ZN(new_n341));
  XNOR2_X1  g140(.A(G8gat), .B(G36gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(G64gat), .B(G92gat), .ZN(new_n343));
  XOR2_X1   g142(.A(new_n342), .B(new_n343), .Z(new_n344));
  NAND3_X1  g143(.A1(new_n339), .A2(new_n341), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT73), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n339), .A2(new_n341), .ZN(new_n348));
  INV_X1    g147(.A(new_n344), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n347), .A2(KEYINPUT30), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT30), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n345), .A2(new_n346), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  XOR2_X1   g153(.A(G113gat), .B(G120gat), .Z(new_n355));
  INV_X1    g154(.A(KEYINPUT1), .ZN(new_n356));
  XNOR2_X1  g155(.A(G127gat), .B(G134gat), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n358), .B(KEYINPUT69), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n355), .A2(new_n356), .ZN(new_n360));
  XOR2_X1   g159(.A(KEYINPUT68), .B(G134gat), .Z(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(G127gat), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n360), .B(new_n362), .C1(G127gat), .C2(G134gat), .ZN(new_n363));
  AND2_X1   g162(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(G155gat), .B(G162gat), .ZN(new_n365));
  XOR2_X1   g164(.A(G141gat), .B(G148gat), .Z(new_n366));
  AOI21_X1  g165(.A(new_n365), .B1(new_n366), .B2(KEYINPUT74), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT2), .ZN(new_n368));
  AND2_X1   g167(.A1(G155gat), .A2(G162gat), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n366), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OR2_X1    g169(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n367), .A2(new_n370), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n364), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT4), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n364), .A2(KEYINPUT4), .A3(new_n374), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n373), .A2(KEYINPUT3), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n359), .A2(new_n363), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT3), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n380), .B1(new_n374), .B2(new_n381), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n377), .B(new_n378), .C1(new_n379), .C2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(G225gat), .A2(G233gat), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT5), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n380), .A2(new_n373), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n375), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(KEYINPUT5), .B1(new_n390), .B2(new_n384), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n391), .B1(new_n385), .B2(new_n383), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n387), .A2(new_n392), .ZN(new_n393));
  XOR2_X1   g192(.A(G1gat), .B(G29gat), .Z(new_n394));
  XNOR2_X1  g193(.A(G57gat), .B(G85gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(KEYINPUT75), .B(KEYINPUT0), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n396), .B(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT6), .B1(new_n393), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n398), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n387), .A2(new_n400), .A3(new_n392), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n387), .A2(KEYINPUT6), .A3(new_n392), .A4(new_n400), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n354), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n338), .B1(new_n379), .B2(KEYINPUT29), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n381), .B1(new_n338), .B2(KEYINPUT29), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n373), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(G22gat), .ZN(new_n410));
  INV_X1    g209(.A(G22gat), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n406), .A2(new_n411), .A3(new_n408), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(G228gat), .ZN(new_n414));
  INV_X1    g213(.A(G233gat), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n410), .A2(G228gat), .A3(G233gat), .A4(new_n412), .ZN(new_n417));
  XNOR2_X1  g216(.A(G78gat), .B(G106gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n418), .B(G50gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(KEYINPUT76), .B(KEYINPUT31), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n419), .B(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n416), .A2(new_n417), .A3(new_n421), .ZN(new_n422));
  AND2_X1   g221(.A1(new_n422), .A2(KEYINPUT79), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(KEYINPUT79), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n416), .A2(new_n417), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n421), .B(KEYINPUT77), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT78), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT78), .ZN(new_n428));
  INV_X1    g227(.A(new_n426), .ZN(new_n429));
  AOI211_X1 g228(.A(new_n428), .B(new_n429), .C1(new_n416), .C2(new_n417), .ZN(new_n430));
  OAI22_X1  g229(.A1(new_n423), .A2(new_n424), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n323), .B(new_n380), .ZN(new_n433));
  INV_X1    g232(.A(G227gat), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n434), .A2(new_n415), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT32), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT33), .B1(new_n433), .B2(new_n435), .ZN(new_n439));
  XNOR2_X1  g238(.A(G15gat), .B(G43gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n440), .B(KEYINPUT70), .ZN(new_n441));
  INV_X1    g240(.A(G71gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n441), .B(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n443), .B(G99gat), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n439), .A2(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n323), .B(new_n364), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT34), .ZN(new_n447));
  INV_X1    g246(.A(new_n435), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n447), .B1(new_n446), .B2(new_n448), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n445), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT34), .B1(new_n433), .B2(new_n435), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n453), .B(new_n449), .C1(new_n439), .C2(new_n444), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n438), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n452), .A2(new_n438), .A3(new_n454), .ZN(new_n457));
  NOR2_X1   g256(.A1(KEYINPUT71), .A2(KEYINPUT36), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT71), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT36), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n456), .B(new_n457), .C1(new_n458), .C2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n457), .ZN(new_n463));
  OAI22_X1  g262(.A1(new_n463), .A2(new_n455), .B1(new_n459), .B2(new_n460), .ZN(new_n464));
  AOI22_X1  g263(.A1(new_n405), .A2(new_n432), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n383), .A2(new_n385), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT80), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT80), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n383), .A2(new_n468), .A3(new_n385), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT39), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n470), .B1(new_n390), .B2(new_n384), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n467), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n467), .A2(new_n469), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n398), .B(new_n472), .C1(new_n473), .C2(KEYINPUT39), .ZN(new_n474));
  XOR2_X1   g273(.A(new_n474), .B(KEYINPUT40), .Z(new_n475));
  NAND2_X1  g274(.A1(new_n401), .A2(KEYINPUT81), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT81), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n387), .A2(new_n477), .A3(new_n392), .A4(new_n400), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n353), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n431), .B1(new_n475), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n348), .A2(KEYINPUT37), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT37), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n339), .A2(new_n482), .A3(new_n341), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n481), .A2(new_n483), .A3(new_n349), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT82), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT82), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n481), .A2(new_n486), .A3(new_n483), .A4(new_n349), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n485), .A2(KEYINPUT38), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT38), .B1(new_n485), .B2(new_n487), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n399), .A2(new_n476), .A3(new_n478), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n490), .A2(new_n403), .A3(new_n345), .ZN(new_n491));
  NOR3_X1   g290(.A1(new_n488), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n465), .B1(new_n480), .B2(new_n492), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n431), .A2(new_n457), .A3(new_n456), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT35), .B1(new_n490), .B2(new_n403), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n494), .A2(KEYINPUT83), .A3(new_n354), .A4(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT83), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(new_n354), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n431), .A2(new_n457), .A3(new_n456), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT35), .B1(new_n405), .B2(new_n499), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n496), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n289), .B1(new_n493), .B2(new_n502), .ZN(new_n503));
  XOR2_X1   g302(.A(G183gat), .B(G211gat), .Z(new_n504));
  AOI21_X1  g303(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n505));
  XOR2_X1   g304(.A(new_n505), .B(KEYINPUT92), .Z(new_n506));
  XOR2_X1   g305(.A(G57gat), .B(G64gat), .Z(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XOR2_X1   g307(.A(G71gat), .B(G78gat), .Z(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT93), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n511), .A2(G57gat), .A3(G64gat), .ZN(new_n512));
  AOI21_X1  g311(.A(G64gat), .B1(new_n511), .B2(G57gat), .ZN(new_n513));
  NOR3_X1   g312(.A1(new_n509), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(new_n506), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  XOR2_X1   g315(.A(KEYINPUT94), .B(KEYINPUT21), .Z(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n518), .A2(G231gat), .A3(G233gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(G127gat), .B(G155gat), .ZN(new_n520));
  XOR2_X1   g319(.A(new_n520), .B(KEYINPUT20), .Z(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(G231gat), .A2(G233gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n516), .A2(new_n523), .A3(new_n517), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n519), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n522), .B1(new_n519), .B2(new_n524), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n504), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n527), .ZN(new_n529));
  INV_X1    g328(.A(new_n504), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n529), .A2(new_n530), .A3(new_n525), .ZN(new_n531));
  AOI22_X1  g330(.A1(new_n508), .A2(new_n509), .B1(new_n514), .B2(new_n506), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n211), .B1(KEYINPUT21), .B2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n528), .A2(new_n531), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n535), .B1(new_n528), .B2(new_n531), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G134gat), .B(G162gat), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT98), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT7), .ZN(new_n545));
  INV_X1    g344(.A(G85gat), .ZN(new_n546));
  INV_X1    g345(.A(G92gat), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(G99gat), .A2(G106gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT8), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT96), .ZN(new_n553));
  OR2_X1    g352(.A1(G85gat), .A2(G92gat), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n553), .B1(new_n552), .B2(new_n554), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n550), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT97), .ZN(new_n558));
  XOR2_X1   g357(.A(G99gat), .B(G106gat), .Z(new_n559));
  INV_X1    g358(.A(KEYINPUT97), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n550), .B(new_n560), .C1(new_n555), .C2(new_n556), .ZN(new_n561));
  AND3_X1   g360(.A1(new_n558), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n559), .B1(new_n558), .B2(new_n561), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n544), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n559), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n552), .A2(new_n554), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT96), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n552), .A2(new_n554), .A3(new_n553), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n560), .B1(new_n569), .B2(new_n550), .ZN(new_n570));
  INV_X1    g369(.A(new_n561), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n565), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n558), .A2(new_n559), .A3(new_n561), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n572), .A2(KEYINPUT98), .A3(new_n573), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n564), .A2(new_n574), .A3(new_n257), .A4(new_n263), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n572), .A2(new_n237), .A3(new_n573), .ZN(new_n576));
  NAND3_X1  g375(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G190gat), .B(G218gat), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n579), .B(KEYINPUT99), .Z(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n575), .A2(new_n578), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n581), .B1(new_n575), .B2(new_n578), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n543), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n584), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n586), .A2(new_n542), .A3(new_n582), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n539), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G230gat), .A2(G233gat), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n516), .B1(new_n562), .B2(new_n563), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n572), .A2(new_n532), .A3(new_n573), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT10), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n572), .A2(KEYINPUT10), .A3(new_n532), .A4(new_n573), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n591), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n590), .B1(new_n592), .B2(new_n593), .ZN(new_n598));
  XNOR2_X1  g397(.A(G120gat), .B(G148gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(G176gat), .B(G204gat), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n599), .B(new_n600), .Z(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  OR3_X1    g401(.A1(new_n597), .A2(new_n598), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT100), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n602), .B1(new_n597), .B2(new_n598), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  OAI211_X1 g405(.A(KEYINPUT100), .B(new_n602), .C1(new_n597), .C2(new_n598), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n589), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(KEYINPUT101), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n606), .A2(new_n607), .ZN(new_n611));
  NOR3_X1   g410(.A1(new_n539), .A2(new_n611), .A3(new_n588), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT101), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n503), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n404), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g418(.A1(new_n616), .A2(new_n353), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(G8gat), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT42), .ZN(new_n622));
  XOR2_X1   g421(.A(KEYINPUT16), .B(G8gat), .Z(new_n623));
  NAND3_X1  g422(.A1(new_n616), .A2(new_n353), .A3(new_n623), .ZN(new_n624));
  AND3_X1   g423(.A1(new_n624), .A2(KEYINPUT102), .A3(new_n622), .ZN(new_n625));
  AOI21_X1  g424(.A(KEYINPUT102), .B1(new_n624), .B2(new_n622), .ZN(new_n626));
  OAI221_X1 g425(.A(new_n621), .B1(new_n622), .B2(new_n624), .C1(new_n625), .C2(new_n626), .ZN(G1325gat));
  NAND2_X1  g426(.A1(new_n462), .A2(new_n464), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n616), .A2(G15gat), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n456), .A2(new_n457), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n503), .A2(new_n632), .A3(new_n615), .ZN(new_n633));
  INV_X1    g432(.A(G15gat), .ZN(new_n634));
  AND3_X1   g433(.A1(new_n633), .A2(KEYINPUT103), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT103), .B1(new_n633), .B2(new_n634), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n630), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT104), .ZN(G1326gat));
  AND2_X1   g437(.A1(new_n503), .A2(new_n432), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n615), .ZN(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT43), .B(G22gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(G1327gat));
  AND2_X1   g441(.A1(new_n611), .A2(KEYINPUT105), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n611), .A2(KEYINPUT105), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n288), .A2(new_n255), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n278), .B1(new_n277), .B2(new_n279), .ZN(new_n648));
  AND4_X1   g447(.A1(new_n278), .A2(new_n283), .A3(new_n279), .A4(new_n285), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n646), .A2(new_n650), .A3(new_n539), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n493), .A2(new_n502), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT106), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n493), .A2(new_n502), .A3(KEYINPUT106), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT107), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n588), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n585), .A2(new_n587), .A3(KEYINPUT107), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n660), .A2(KEYINPUT44), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n654), .A2(new_n655), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n663), .B1(new_n652), .B2(new_n588), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n651), .B1(new_n662), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n225), .B1(new_n666), .B2(new_n617), .ZN(new_n667));
  INV_X1    g466(.A(new_n588), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n611), .A2(new_n538), .A3(new_n668), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n503), .A2(new_n225), .A3(new_n617), .A4(new_n669), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n670), .B(KEYINPUT45), .Z(new_n671));
  OAI21_X1  g470(.A(KEYINPUT108), .B1(new_n667), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT108), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n670), .B(KEYINPUT45), .ZN(new_n674));
  AOI211_X1 g473(.A(new_n404), .B(new_n651), .C1(new_n662), .C2(new_n665), .ZN(new_n675));
  OAI211_X1 g474(.A(new_n673), .B(new_n674), .C1(new_n675), .C2(new_n225), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n672), .A2(new_n676), .ZN(G1328gat));
  INV_X1    g476(.A(KEYINPUT109), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n226), .B1(new_n666), .B2(new_n353), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n503), .A2(new_n226), .A3(new_n353), .A4(new_n669), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT46), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n678), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT46), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n680), .B(new_n683), .ZN(new_n684));
  AOI211_X1 g483(.A(new_n354), .B(new_n651), .C1(new_n662), .C2(new_n665), .ZN(new_n685));
  OAI211_X1 g484(.A(KEYINPUT109), .B(new_n684), .C1(new_n685), .C2(new_n226), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n682), .A2(new_n686), .ZN(G1329gat));
  NOR2_X1   g486(.A1(new_n628), .A2(new_n216), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n666), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n503), .A2(new_n632), .A3(new_n669), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(new_n216), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(KEYINPUT47), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT47), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n689), .A2(new_n694), .A3(new_n691), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n695), .ZN(G1330gat));
  INV_X1    g495(.A(KEYINPUT48), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n213), .B1(new_n666), .B2(new_n432), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n639), .A2(new_n213), .A3(new_n669), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n697), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  AOI211_X1 g500(.A(new_n431), .B(new_n651), .C1(new_n662), .C2(new_n665), .ZN(new_n702));
  OAI211_X1 g501(.A(KEYINPUT48), .B(new_n699), .C1(new_n702), .C2(new_n213), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n701), .A2(new_n703), .ZN(G1331gat));
  AND3_X1   g503(.A1(new_n493), .A2(new_n502), .A3(KEYINPUT106), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT106), .B1(new_n493), .B2(new_n502), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n645), .A2(new_n289), .A3(new_n589), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n617), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n353), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n713), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n714));
  XOR2_X1   g513(.A(KEYINPUT49), .B(G64gat), .Z(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(new_n713), .B2(new_n715), .ZN(G1333gat));
  OAI21_X1  g515(.A(G71gat), .B1(new_n709), .B2(new_n628), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n707), .A2(new_n442), .A3(new_n632), .A4(new_n708), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(G1334gat));
  NAND2_X1  g523(.A1(new_n710), .A2(new_n432), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g525(.A1(new_n650), .A2(new_n538), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n652), .A2(new_n588), .A3(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT51), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT112), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n652), .A2(KEYINPUT51), .A3(new_n588), .A4(new_n727), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n728), .A2(KEYINPUT112), .A3(new_n729), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n404), .A2(G85gat), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n733), .A2(new_n611), .A3(new_n734), .A4(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n727), .A2(new_n611), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n661), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n705), .A2(new_n706), .A3(new_n739), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n617), .B(new_n738), .C1(new_n740), .C2(new_n664), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT111), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(G85gat), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n741), .A2(new_n742), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n736), .B1(new_n744), .B2(new_n745), .ZN(G1336gat));
  OAI211_X1 g545(.A(new_n353), .B(new_n738), .C1(new_n740), .C2(new_n664), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(G92gat), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT52), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n646), .A2(G92gat), .A3(new_n354), .ZN(new_n751));
  AND3_X1   g550(.A1(new_n733), .A2(new_n734), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n730), .A2(new_n732), .ZN(new_n753));
  AOI22_X1  g552(.A1(new_n747), .A2(G92gat), .B1(new_n753), .B2(new_n751), .ZN(new_n754));
  OAI22_X1  g553(.A1(new_n750), .A2(new_n752), .B1(new_n754), .B2(new_n749), .ZN(G1337gat));
  NOR2_X1   g554(.A1(new_n631), .A2(G99gat), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n733), .A2(new_n611), .A3(new_n734), .A4(new_n756), .ZN(new_n757));
  AOI211_X1 g556(.A(new_n628), .B(new_n737), .C1(new_n662), .C2(new_n665), .ZN(new_n758));
  INV_X1    g557(.A(G99gat), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(G1338gat));
  OAI211_X1 g559(.A(new_n432), .B(new_n738), .C1(new_n740), .C2(new_n664), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G106gat), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT53), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n646), .A2(G106gat), .A3(new_n431), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n733), .A2(new_n734), .A3(new_n765), .ZN(new_n766));
  AOI22_X1  g565(.A1(new_n761), .A2(G106gat), .B1(new_n753), .B2(new_n765), .ZN(new_n767));
  OAI22_X1  g566(.A1(new_n764), .A2(new_n766), .B1(new_n767), .B2(new_n763), .ZN(G1339gat));
  NOR2_X1   g567(.A1(new_n609), .A2(new_n650), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n265), .A2(new_n238), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n771), .A2(G229gat), .A3(G233gat), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n246), .A2(new_n248), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n775), .A2(new_n254), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n611), .B(new_n777), .C1(new_n648), .C2(new_n649), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n595), .A2(new_n596), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n590), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n595), .A2(new_n596), .A3(new_n591), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n781), .A2(KEYINPUT54), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n601), .B1(new_n597), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n783), .A2(KEYINPUT55), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n603), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT55), .B1(new_n783), .B2(new_n785), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n779), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n790));
  INV_X1    g589(.A(new_n782), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n791), .A2(new_n597), .A3(new_n784), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n780), .A2(new_n784), .A3(new_n590), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n602), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n790), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n795), .A2(KEYINPUT113), .A3(new_n603), .A4(new_n786), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n789), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n778), .B1(new_n797), .B2(new_n289), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n777), .B1(new_n648), .B2(new_n649), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n789), .A2(new_n659), .A3(new_n796), .ZN(new_n801));
  AOI22_X1  g600(.A1(new_n798), .A2(new_n660), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n770), .B1(new_n802), .B2(new_n538), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n804), .A2(new_n432), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n404), .A2(new_n353), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n805), .A2(new_n632), .A3(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(G113gat), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n807), .A2(new_n808), .A3(new_n289), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n804), .A2(new_n404), .A3(new_n499), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n354), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n650), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n809), .B1(new_n813), .B2(new_n808), .ZN(G1340gat));
  INV_X1    g613(.A(G120gat), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n807), .A2(new_n815), .A3(new_n646), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n812), .A2(new_n611), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n816), .B1(new_n817), .B2(new_n815), .ZN(G1341gat));
  OAI21_X1  g617(.A(G127gat), .B1(new_n807), .B2(new_n539), .ZN(new_n819));
  OR2_X1    g618(.A1(new_n539), .A2(G127gat), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n819), .B1(new_n811), .B2(new_n820), .ZN(G1342gat));
  NOR2_X1   g620(.A1(new_n353), .A2(new_n668), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n822), .B(KEYINPUT114), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n823), .A2(new_n361), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n810), .A2(new_n824), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n825), .A2(KEYINPUT56), .ZN(new_n826));
  OAI21_X1  g625(.A(G134gat), .B1(new_n807), .B2(new_n668), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(KEYINPUT56), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(G1343gat));
  AND2_X1   g628(.A1(new_n628), .A2(new_n806), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n788), .A2(KEYINPUT116), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n832));
  AOI211_X1 g631(.A(new_n832), .B(KEYINPUT55), .C1(new_n783), .C2(new_n785), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n603), .B(new_n786), .C1(new_n831), .C2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n289), .A2(new_n834), .ZN(new_n835));
  AOI211_X1 g634(.A(new_n776), .B(new_n608), .C1(new_n287), .C2(new_n280), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n668), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n801), .A2(new_n800), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n538), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI211_X1 g638(.A(KEYINPUT57), .B(new_n432), .C1(new_n839), .C2(new_n769), .ZN(new_n840));
  AOI21_X1  g639(.A(KEYINPUT57), .B1(new_n803), .B2(new_n432), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n840), .B1(new_n841), .B2(KEYINPUT115), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n798), .A2(new_n660), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n538), .B1(new_n843), .B2(new_n838), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n432), .B1(new_n844), .B2(new_n769), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n845), .A2(KEYINPUT115), .A3(new_n846), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n650), .B(new_n830), .C1(new_n842), .C2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(G141gat), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n629), .A2(new_n431), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n803), .A2(new_n850), .A3(new_n617), .A4(new_n354), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n289), .A2(G141gat), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT117), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT118), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n854), .B(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n849), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(KEYINPUT58), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n854), .A2(KEYINPUT119), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n851), .A2(new_n860), .A3(new_n853), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n859), .A2(KEYINPUT58), .A3(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT120), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n849), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n863), .B1(new_n849), .B2(new_n862), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n858), .B1(new_n864), .B2(new_n865), .ZN(G1344gat));
  INV_X1    g665(.A(G148gat), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n867), .A2(KEYINPUT59), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n830), .B1(new_n842), .B2(new_n847), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n868), .B1(new_n869), .B2(new_n608), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT123), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n431), .A2(KEYINPUT57), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n795), .A2(new_n588), .A3(new_n603), .A4(new_n786), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n799), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n538), .B1(new_n837), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n610), .A2(new_n289), .A3(new_n614), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n872), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n461), .B1(new_n456), .B2(new_n457), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n461), .A2(new_n458), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n463), .A2(new_n455), .A3(new_n881), .ZN(new_n882));
  OAI211_X1 g681(.A(KEYINPUT121), .B(new_n806), .C1(new_n880), .C2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n611), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT121), .B1(new_n628), .B2(new_n806), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n650), .A2(new_n789), .A3(new_n796), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n659), .B1(new_n887), .B2(new_n778), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n797), .A2(new_n799), .A3(new_n660), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n539), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n431), .B1(new_n890), .B2(new_n770), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n879), .B(new_n886), .C1(new_n891), .C2(new_n846), .ZN(new_n892));
  OAI21_X1  g691(.A(G148gat), .B1(new_n892), .B2(KEYINPUT122), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT122), .ZN(new_n894));
  INV_X1    g693(.A(new_n872), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n795), .A2(new_n832), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n788), .A2(KEYINPUT116), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n787), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n650), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n588), .B1(new_n899), .B2(new_n778), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n539), .B1(new_n900), .B2(new_n874), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n895), .B1(new_n901), .B2(new_n877), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n902), .B1(new_n845), .B2(KEYINPUT57), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n894), .B1(new_n903), .B2(new_n886), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n871), .B(KEYINPUT59), .C1(new_n893), .C2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n892), .A2(KEYINPUT122), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n845), .A2(KEYINPUT57), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n908), .A2(new_n894), .A3(new_n879), .A4(new_n886), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n907), .A2(G148gat), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n871), .B1(new_n910), .B2(KEYINPUT59), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n870), .B1(new_n906), .B2(new_n911), .ZN(new_n912));
  OR3_X1    g711(.A1(new_n851), .A2(G148gat), .A3(new_n608), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(G1345gat));
  OAI21_X1  g713(.A(G155gat), .B1(new_n869), .B2(new_n539), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n539), .A2(G155gat), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n915), .B1(new_n851), .B2(new_n916), .ZN(G1346gat));
  OAI21_X1  g716(.A(G162gat), .B1(new_n869), .B2(new_n660), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n823), .A2(G162gat), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n919), .A2(new_n803), .A3(new_n617), .A4(new_n850), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(G1347gat));
  NAND2_X1  g720(.A1(new_n404), .A2(new_n353), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT124), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n923), .A2(new_n631), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n805), .A2(new_n924), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n925), .A2(new_n291), .A3(new_n289), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n804), .A2(new_n617), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n499), .A2(new_n354), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n650), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n926), .B1(new_n931), .B2(new_n291), .ZN(G1348gat));
  OAI21_X1  g731(.A(new_n292), .B1(new_n929), .B2(new_n608), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT125), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n925), .A2(new_n292), .A3(new_n646), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n934), .A2(new_n935), .ZN(G1349gat));
  NAND3_X1  g735(.A1(new_n930), .A2(new_n300), .A3(new_n538), .ZN(new_n937));
  OAI21_X1  g736(.A(G183gat), .B1(new_n925), .B2(new_n539), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n937), .A2(KEYINPUT126), .A3(new_n938), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g739(.A(G190gat), .B1(new_n925), .B2(new_n668), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT61), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n659), .A2(new_n301), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n942), .B1(new_n929), .B2(new_n943), .ZN(G1351gat));
  NOR3_X1   g743(.A1(new_n629), .A2(new_n431), .A3(new_n354), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n927), .A2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(G197gat), .B1(new_n947), .B2(new_n650), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n908), .A2(new_n879), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n923), .A2(new_n629), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n650), .A2(G197gat), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n948), .B1(new_n951), .B2(new_n952), .ZN(G1352gat));
  INV_X1    g752(.A(G204gat), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n951), .A2(new_n645), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT127), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n957), .B1(new_n956), .B2(new_n955), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n946), .A2(G204gat), .A3(new_n608), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT62), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n960), .ZN(G1353gat));
  NAND3_X1  g760(.A1(new_n947), .A2(new_n329), .A3(new_n538), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n951), .A2(new_n538), .ZN(new_n963));
  AND3_X1   g762(.A1(new_n963), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n964));
  AOI21_X1  g763(.A(KEYINPUT63), .B1(new_n963), .B2(G211gat), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(G1354gat));
  NAND3_X1  g765(.A1(new_n947), .A2(new_n330), .A3(new_n659), .ZN(new_n967));
  NOR3_X1   g766(.A1(new_n949), .A2(new_n668), .A3(new_n950), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n967), .B1(new_n968), .B2(new_n330), .ZN(G1355gat));
endmodule


